VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO meta_srlatch_array_row
  CLASS BLOCK ;
  FOREIGN meta_srlatch_array_row ;
  ORIGIN 310.220 182.150 ;
  SIZE 474.570 BY 547.550 ;
  SITE unithd ;
  PIN o_ranQ[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 18.315 89.065 18.820 89.145 ;
        RECT 19.620 89.065 20.525 89.155 ;
        RECT 18.315 88.885 20.525 89.065 ;
      LAYER mcon ;
        RECT 18.505 88.975 18.675 89.145 ;
        RECT 19.870 88.975 20.040 89.145 ;
      LAYER met1 ;
        RECT 18.440 88.880 20.130 89.180 ;
        RECT 18.620 88.180 19.620 88.880 ;
    END
  END o_ranQ[1]
  PIN o_ranQ[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 13.355 94.875 15.565 95.055 ;
        RECT 13.355 94.795 13.860 94.875 ;
        RECT 14.660 94.785 15.565 94.875 ;
      LAYER mcon ;
        RECT 13.545 94.795 13.715 94.965 ;
        RECT 14.910 94.795 15.080 94.965 ;
      LAYER met1 ;
        RECT 13.660 95.060 14.660 95.760 ;
        RECT 13.480 94.760 15.170 95.060 ;
    END
  END o_ranQ[2]
  PIN o_ranQ[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 8.395 89.065 8.900 89.145 ;
        RECT 9.700 89.065 10.605 89.155 ;
        RECT 8.395 88.885 10.605 89.065 ;
      LAYER mcon ;
        RECT 8.585 88.975 8.755 89.145 ;
        RECT 9.950 88.975 10.120 89.145 ;
      LAYER met1 ;
        RECT 8.520 88.880 10.210 89.180 ;
        RECT 8.700 88.180 9.700 88.880 ;
    END
  END o_ranQ[3]
  PIN o_ranQ[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 23.275 94.875 25.485 95.055 ;
        RECT 23.275 94.795 23.780 94.875 ;
        RECT 24.580 94.785 25.485 94.875 ;
      LAYER mcon ;
        RECT 23.465 94.795 23.635 94.965 ;
        RECT 24.830 94.795 25.000 94.965 ;
      LAYER met1 ;
        RECT 23.580 95.060 24.580 95.760 ;
        RECT 23.400 94.760 25.090 95.060 ;
    END
  END o_ranQ[0]
  PIN o_ranQ[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 3.435 94.875 5.645 95.055 ;
        RECT 3.435 94.795 3.940 94.875 ;
        RECT 4.740 94.785 5.645 94.875 ;
      LAYER mcon ;
        RECT 3.625 94.795 3.795 94.965 ;
        RECT 4.990 94.795 5.160 94.965 ;
      LAYER met1 ;
        RECT 3.740 95.060 4.740 95.760 ;
        RECT 3.560 94.760 5.250 95.060 ;
    END
  END o_ranQ[4]
  PIN o_ranQ[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -1.525 89.065 -1.020 89.145 ;
        RECT -0.220 89.065 0.685 89.155 ;
        RECT -1.525 88.885 0.685 89.065 ;
      LAYER mcon ;
        RECT -1.335 88.975 -1.165 89.145 ;
        RECT 0.030 88.975 0.200 89.145 ;
      LAYER met1 ;
        RECT -1.400 88.880 0.290 89.180 ;
        RECT -1.220 88.180 -0.220 88.880 ;
    END
  END o_ranQ[5]
  PIN o_ranQ[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -6.485 94.875 -4.275 95.055 ;
        RECT -6.485 94.795 -5.980 94.875 ;
        RECT -5.180 94.785 -4.275 94.875 ;
      LAYER mcon ;
        RECT -6.295 94.795 -6.125 94.965 ;
        RECT -4.930 94.795 -4.760 94.965 ;
      LAYER met1 ;
        RECT -6.180 95.060 -5.180 95.760 ;
        RECT -6.360 94.760 -4.670 95.060 ;
    END
  END o_ranQ[6]
  PIN o_ranQ[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -11.445 89.065 -10.940 89.145 ;
        RECT -10.140 89.065 -9.235 89.155 ;
        RECT -11.445 88.885 -9.235 89.065 ;
      LAYER mcon ;
        RECT -11.255 88.975 -11.085 89.145 ;
        RECT -9.890 88.975 -9.720 89.145 ;
      LAYER met1 ;
        RECT -11.320 88.880 -9.630 89.180 ;
        RECT -11.140 88.180 -10.140 88.880 ;
    END
  END o_ranQ[7]
  PIN o_ranQ[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -16.405 94.875 -14.195 95.055 ;
        RECT -16.405 94.795 -15.900 94.875 ;
        RECT -15.100 94.785 -14.195 94.875 ;
      LAYER mcon ;
        RECT -16.215 94.795 -16.045 94.965 ;
        RECT -14.850 94.795 -14.680 94.965 ;
      LAYER met1 ;
        RECT -16.100 95.060 -15.100 95.760 ;
        RECT -16.280 94.760 -14.590 95.060 ;
    END
  END o_ranQ[8]
  PIN o_ranQ[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -21.365 89.065 -20.860 89.145 ;
        RECT -20.060 89.065 -19.155 89.155 ;
        RECT -21.365 88.885 -19.155 89.065 ;
      LAYER mcon ;
        RECT -21.175 88.975 -21.005 89.145 ;
        RECT -19.810 88.975 -19.640 89.145 ;
      LAYER met1 ;
        RECT -21.240 88.880 -19.550 89.180 ;
        RECT -21.060 88.180 -20.060 88.880 ;
    END
  END o_ranQ[9]
  PIN o_ranQ[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -26.325 94.875 -24.115 95.055 ;
        RECT -26.325 94.795 -25.820 94.875 ;
        RECT -25.020 94.785 -24.115 94.875 ;
      LAYER mcon ;
        RECT -26.135 94.795 -25.965 94.965 ;
        RECT -24.770 94.795 -24.600 94.965 ;
      LAYER met1 ;
        RECT -26.020 95.060 -25.020 95.760 ;
        RECT -26.200 94.760 -24.510 95.060 ;
    END
  END o_ranQ[10]
  PIN o_ranQ[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -31.285 89.065 -30.780 89.145 ;
        RECT -29.980 89.065 -29.075 89.155 ;
        RECT -31.285 88.885 -29.075 89.065 ;
      LAYER mcon ;
        RECT -31.095 88.975 -30.925 89.145 ;
        RECT -29.730 88.975 -29.560 89.145 ;
      LAYER met1 ;
        RECT -31.160 88.880 -29.470 89.180 ;
        RECT -30.980 88.180 -29.980 88.880 ;
    END
  END o_ranQ[11]
  PIN o_ranQ[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -36.245 94.875 -34.035 95.055 ;
        RECT -36.245 94.795 -35.740 94.875 ;
        RECT -34.940 94.785 -34.035 94.875 ;
      LAYER mcon ;
        RECT -36.055 94.795 -35.885 94.965 ;
        RECT -34.690 94.795 -34.520 94.965 ;
      LAYER met1 ;
        RECT -35.940 95.060 -34.940 95.760 ;
        RECT -36.120 94.760 -34.430 95.060 ;
    END
  END o_ranQ[12]
  PIN o_ranQ[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -41.205 89.065 -40.700 89.145 ;
        RECT -39.900 89.065 -38.995 89.155 ;
        RECT -41.205 88.885 -38.995 89.065 ;
      LAYER mcon ;
        RECT -41.015 88.975 -40.845 89.145 ;
        RECT -39.650 88.975 -39.480 89.145 ;
      LAYER met1 ;
        RECT -41.080 88.880 -39.390 89.180 ;
        RECT -40.900 88.180 -39.900 88.880 ;
    END
  END o_ranQ[13]
  PIN o_ranQ[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -46.165 94.875 -43.955 95.055 ;
        RECT -46.165 94.795 -45.660 94.875 ;
        RECT -44.860 94.785 -43.955 94.875 ;
      LAYER mcon ;
        RECT -45.975 94.795 -45.805 94.965 ;
        RECT -44.610 94.795 -44.440 94.965 ;
      LAYER met1 ;
        RECT -45.860 95.060 -44.860 95.760 ;
        RECT -46.040 94.760 -44.350 95.060 ;
    END
  END o_ranQ[14]
  PIN o_ranQ[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -51.125 89.065 -50.620 89.145 ;
        RECT -49.820 89.065 -48.915 89.155 ;
        RECT -51.125 88.885 -48.915 89.065 ;
      LAYER mcon ;
        RECT -50.935 88.975 -50.765 89.145 ;
        RECT -49.570 88.975 -49.400 89.145 ;
      LAYER met1 ;
        RECT -51.000 88.880 -49.310 89.180 ;
        RECT -50.820 88.180 -49.820 88.880 ;
    END
  END o_ranQ[15]
  PIN o_ranQ[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -61.045 89.065 -60.540 89.145 ;
        RECT -59.740 89.065 -58.835 89.155 ;
        RECT -61.045 88.885 -58.835 89.065 ;
      LAYER mcon ;
        RECT -60.855 88.975 -60.685 89.145 ;
        RECT -59.490 88.975 -59.320 89.145 ;
      LAYER met1 ;
        RECT -60.920 88.880 -59.230 89.180 ;
        RECT -60.740 88.180 -59.740 88.880 ;
    END
  END o_ranQ[17]
  PIN o_ranQ[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -66.005 94.875 -63.795 95.055 ;
        RECT -66.005 94.795 -65.500 94.875 ;
        RECT -64.700 94.785 -63.795 94.875 ;
      LAYER mcon ;
        RECT -65.815 94.795 -65.645 94.965 ;
        RECT -64.450 94.795 -64.280 94.965 ;
      LAYER met1 ;
        RECT -65.700 95.060 -64.700 95.760 ;
        RECT -65.880 94.760 -64.190 95.060 ;
    END
  END o_ranQ[18]
  PIN o_ranQ[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -70.965 89.065 -70.460 89.145 ;
        RECT -69.660 89.065 -68.755 89.155 ;
        RECT -70.965 88.885 -68.755 89.065 ;
      LAYER mcon ;
        RECT -70.775 88.975 -70.605 89.145 ;
        RECT -69.410 88.975 -69.240 89.145 ;
      LAYER met1 ;
        RECT -70.840 88.880 -69.150 89.180 ;
        RECT -70.660 88.180 -69.660 88.880 ;
    END
  END o_ranQ[19]
  PIN o_ranQ[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -56.085 94.875 -53.875 95.055 ;
        RECT -56.085 94.795 -55.580 94.875 ;
        RECT -54.780 94.785 -53.875 94.875 ;
      LAYER mcon ;
        RECT -55.895 94.795 -55.725 94.965 ;
        RECT -54.530 94.795 -54.360 94.965 ;
      LAYER met1 ;
        RECT -55.780 95.060 -54.780 95.760 ;
        RECT -55.960 94.760 -54.270 95.060 ;
    END
  END o_ranQ[16]
  PIN o_ranQ[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -75.925 94.875 -73.715 95.055 ;
        RECT -75.925 94.795 -75.420 94.875 ;
        RECT -74.620 94.785 -73.715 94.875 ;
      LAYER mcon ;
        RECT -75.735 94.795 -75.565 94.965 ;
        RECT -74.370 94.795 -74.200 94.965 ;
      LAYER met1 ;
        RECT -75.620 95.060 -74.620 95.760 ;
        RECT -75.800 94.760 -74.110 95.060 ;
    END
  END o_ranQ[20]
  PIN o_ranQ[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -80.885 89.065 -80.380 89.145 ;
        RECT -79.580 89.065 -78.675 89.155 ;
        RECT -80.885 88.885 -78.675 89.065 ;
      LAYER mcon ;
        RECT -80.695 88.975 -80.525 89.145 ;
        RECT -79.330 88.975 -79.160 89.145 ;
      LAYER met1 ;
        RECT -80.760 88.880 -79.070 89.180 ;
        RECT -80.580 88.180 -79.580 88.880 ;
    END
  END o_ranQ[21]
  PIN o_ranQ[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -85.845 94.875 -83.635 95.055 ;
        RECT -85.845 94.795 -85.340 94.875 ;
        RECT -84.540 94.785 -83.635 94.875 ;
      LAYER mcon ;
        RECT -85.655 94.795 -85.485 94.965 ;
        RECT -84.290 94.795 -84.120 94.965 ;
      LAYER met1 ;
        RECT -85.540 95.060 -84.540 95.760 ;
        RECT -85.720 94.760 -84.030 95.060 ;
    END
  END o_ranQ[22]
  PIN o_ranQ[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -90.805 89.065 -90.300 89.145 ;
        RECT -89.500 89.065 -88.595 89.155 ;
        RECT -90.805 88.885 -88.595 89.065 ;
      LAYER mcon ;
        RECT -90.615 88.975 -90.445 89.145 ;
        RECT -89.250 88.975 -89.080 89.145 ;
      LAYER met1 ;
        RECT -90.680 88.880 -88.990 89.180 ;
        RECT -90.500 88.180 -89.500 88.880 ;
    END
  END o_ranQ[23]
  PIN o_ranQ[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -95.765 94.875 -93.555 95.055 ;
        RECT -95.765 94.795 -95.260 94.875 ;
        RECT -94.460 94.785 -93.555 94.875 ;
      LAYER mcon ;
        RECT -95.575 94.795 -95.405 94.965 ;
        RECT -94.210 94.795 -94.040 94.965 ;
      LAYER met1 ;
        RECT -95.460 95.060 -94.460 95.760 ;
        RECT -95.640 94.760 -93.950 95.060 ;
    END
  END o_ranQ[24]
  PIN o_ranQ[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -100.725 89.065 -100.220 89.145 ;
        RECT -99.420 89.065 -98.515 89.155 ;
        RECT -100.725 88.885 -98.515 89.065 ;
      LAYER mcon ;
        RECT -100.535 88.975 -100.365 89.145 ;
        RECT -99.170 88.975 -99.000 89.145 ;
      LAYER met1 ;
        RECT -100.600 88.880 -98.910 89.180 ;
        RECT -100.420 88.180 -99.420 88.880 ;
    END
  END o_ranQ[25]
  PIN o_ranQ[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -105.685 94.875 -103.475 95.055 ;
        RECT -105.685 94.795 -105.180 94.875 ;
        RECT -104.380 94.785 -103.475 94.875 ;
      LAYER mcon ;
        RECT -105.495 94.795 -105.325 94.965 ;
        RECT -104.130 94.795 -103.960 94.965 ;
      LAYER met1 ;
        RECT -105.380 95.060 -104.380 95.760 ;
        RECT -105.560 94.760 -103.870 95.060 ;
    END
  END o_ranQ[26]
  PIN o_ranQ[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -110.645 89.065 -110.140 89.145 ;
        RECT -109.340 89.065 -108.435 89.155 ;
        RECT -110.645 88.885 -108.435 89.065 ;
      LAYER mcon ;
        RECT -110.455 88.975 -110.285 89.145 ;
        RECT -109.090 88.975 -108.920 89.145 ;
      LAYER met1 ;
        RECT -110.520 88.880 -108.830 89.180 ;
        RECT -110.340 88.180 -109.340 88.880 ;
    END
  END o_ranQ[27]
  PIN o_ranQ[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -115.605 94.875 -113.395 95.055 ;
        RECT -115.605 94.795 -115.100 94.875 ;
        RECT -114.300 94.785 -113.395 94.875 ;
      LAYER mcon ;
        RECT -115.415 94.795 -115.245 94.965 ;
        RECT -114.050 94.795 -113.880 94.965 ;
      LAYER met1 ;
        RECT -115.300 95.060 -114.300 95.760 ;
        RECT -115.480 94.760 -113.790 95.060 ;
    END
  END o_ranQ[28]
  PIN o_ranQ[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -120.565 89.065 -120.060 89.145 ;
        RECT -119.260 89.065 -118.355 89.155 ;
        RECT -120.565 88.885 -118.355 89.065 ;
      LAYER mcon ;
        RECT -120.375 88.975 -120.205 89.145 ;
        RECT -119.010 88.975 -118.840 89.145 ;
      LAYER met1 ;
        RECT -120.440 88.880 -118.750 89.180 ;
        RECT -120.260 88.180 -119.260 88.880 ;
    END
  END o_ranQ[29]
  PIN o_ranQ[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -125.525 94.875 -123.315 95.055 ;
        RECT -125.525 94.795 -125.020 94.875 ;
        RECT -124.220 94.785 -123.315 94.875 ;
      LAYER mcon ;
        RECT -125.335 94.795 -125.165 94.965 ;
        RECT -123.970 94.795 -123.800 94.965 ;
      LAYER met1 ;
        RECT -125.220 95.060 -124.220 95.760 ;
        RECT -125.400 94.760 -123.710 95.060 ;
    END
  END o_ranQ[30]
  PIN o_ranQ[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -130.485 89.065 -129.980 89.145 ;
        RECT -129.180 89.065 -128.275 89.155 ;
        RECT -130.485 88.885 -128.275 89.065 ;
      LAYER mcon ;
        RECT -130.295 88.975 -130.125 89.145 ;
        RECT -128.930 88.975 -128.760 89.145 ;
      LAYER met1 ;
        RECT -130.360 88.880 -128.670 89.180 ;
        RECT -130.180 88.180 -129.180 88.880 ;
    END
  END o_ranQ[31]
  PIN o_ranQ[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -140.405 89.065 -139.900 89.145 ;
        RECT -139.100 89.065 -138.195 89.155 ;
        RECT -140.405 88.885 -138.195 89.065 ;
      LAYER mcon ;
        RECT -140.215 88.975 -140.045 89.145 ;
        RECT -138.850 88.975 -138.680 89.145 ;
      LAYER met1 ;
        RECT -140.280 88.880 -138.590 89.180 ;
        RECT -140.100 88.180 -139.100 88.880 ;
    END
  END o_ranQ[33]
  PIN o_ranQ[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -145.365 94.875 -143.155 95.055 ;
        RECT -145.365 94.795 -144.860 94.875 ;
        RECT -144.060 94.785 -143.155 94.875 ;
      LAYER mcon ;
        RECT -145.175 94.795 -145.005 94.965 ;
        RECT -143.810 94.795 -143.640 94.965 ;
      LAYER met1 ;
        RECT -145.060 95.060 -144.060 95.760 ;
        RECT -145.240 94.760 -143.550 95.060 ;
    END
  END o_ranQ[34]
  PIN o_ranQ[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -150.325 89.065 -149.820 89.145 ;
        RECT -149.020 89.065 -148.115 89.155 ;
        RECT -150.325 88.885 -148.115 89.065 ;
      LAYER mcon ;
        RECT -150.135 88.975 -149.965 89.145 ;
        RECT -148.770 88.975 -148.600 89.145 ;
      LAYER met1 ;
        RECT -150.200 88.880 -148.510 89.180 ;
        RECT -150.020 88.180 -149.020 88.880 ;
    END
  END o_ranQ[35]
  PIN o_ranQ[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -135.445 94.875 -133.235 95.055 ;
        RECT -135.445 94.795 -134.940 94.875 ;
        RECT -134.140 94.785 -133.235 94.875 ;
      LAYER mcon ;
        RECT -135.255 94.795 -135.085 94.965 ;
        RECT -133.890 94.795 -133.720 94.965 ;
      LAYER met1 ;
        RECT -135.140 95.060 -134.140 95.760 ;
        RECT -135.320 94.760 -133.630 95.060 ;
    END
  END o_ranQ[32]
  PIN o_ranQ[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -155.285 94.875 -153.075 95.055 ;
        RECT -155.285 94.795 -154.780 94.875 ;
        RECT -153.980 94.785 -153.075 94.875 ;
      LAYER mcon ;
        RECT -155.095 94.795 -154.925 94.965 ;
        RECT -153.730 94.795 -153.560 94.965 ;
      LAYER met1 ;
        RECT -154.980 95.060 -153.980 95.760 ;
        RECT -155.160 94.760 -153.470 95.060 ;
    END
  END o_ranQ[36]
  PIN o_ranQ[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -160.245 89.065 -159.740 89.145 ;
        RECT -158.940 89.065 -158.035 89.155 ;
        RECT -160.245 88.885 -158.035 89.065 ;
      LAYER mcon ;
        RECT -160.055 88.975 -159.885 89.145 ;
        RECT -158.690 88.975 -158.520 89.145 ;
      LAYER met1 ;
        RECT -160.120 88.880 -158.430 89.180 ;
        RECT -159.940 88.180 -158.940 88.880 ;
    END
  END o_ranQ[37]
  PIN o_ranQ[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -165.205 94.875 -162.995 95.055 ;
        RECT -165.205 94.795 -164.700 94.875 ;
        RECT -163.900 94.785 -162.995 94.875 ;
      LAYER mcon ;
        RECT -165.015 94.795 -164.845 94.965 ;
        RECT -163.650 94.795 -163.480 94.965 ;
      LAYER met1 ;
        RECT -164.900 95.060 -163.900 95.760 ;
        RECT -165.080 94.760 -163.390 95.060 ;
    END
  END o_ranQ[38]
  PIN o_ranQ[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -170.165 89.065 -169.660 89.145 ;
        RECT -168.860 89.065 -167.955 89.155 ;
        RECT -170.165 88.885 -167.955 89.065 ;
      LAYER mcon ;
        RECT -169.975 88.975 -169.805 89.145 ;
        RECT -168.610 88.975 -168.440 89.145 ;
      LAYER met1 ;
        RECT -170.040 88.880 -168.350 89.180 ;
        RECT -169.860 88.180 -168.860 88.880 ;
    END
  END o_ranQ[39]
  PIN o_ranQ[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -175.125 94.875 -172.915 95.055 ;
        RECT -175.125 94.795 -174.620 94.875 ;
        RECT -173.820 94.785 -172.915 94.875 ;
      LAYER mcon ;
        RECT -174.935 94.795 -174.765 94.965 ;
        RECT -173.570 94.795 -173.400 94.965 ;
      LAYER met1 ;
        RECT -174.820 95.060 -173.820 95.760 ;
        RECT -175.000 94.760 -173.310 95.060 ;
    END
  END o_ranQ[40]
  PIN o_ranQ[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -180.085 89.065 -179.580 89.145 ;
        RECT -178.780 89.065 -177.875 89.155 ;
        RECT -180.085 88.885 -177.875 89.065 ;
      LAYER mcon ;
        RECT -179.895 88.975 -179.725 89.145 ;
        RECT -178.530 88.975 -178.360 89.145 ;
      LAYER met1 ;
        RECT -179.960 88.880 -178.270 89.180 ;
        RECT -179.780 88.180 -178.780 88.880 ;
    END
  END o_ranQ[41]
  PIN o_ranQ[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -185.045 94.875 -182.835 95.055 ;
        RECT -185.045 94.795 -184.540 94.875 ;
        RECT -183.740 94.785 -182.835 94.875 ;
      LAYER mcon ;
        RECT -184.855 94.795 -184.685 94.965 ;
        RECT -183.490 94.795 -183.320 94.965 ;
      LAYER met1 ;
        RECT -184.740 95.060 -183.740 95.760 ;
        RECT -184.920 94.760 -183.230 95.060 ;
    END
  END o_ranQ[42]
  PIN o_ranQ[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -190.005 89.065 -189.500 89.145 ;
        RECT -188.700 89.065 -187.795 89.155 ;
        RECT -190.005 88.885 -187.795 89.065 ;
      LAYER mcon ;
        RECT -189.815 88.975 -189.645 89.145 ;
        RECT -188.450 88.975 -188.280 89.145 ;
      LAYER met1 ;
        RECT -189.880 88.880 -188.190 89.180 ;
        RECT -189.700 88.180 -188.700 88.880 ;
    END
  END o_ranQ[43]
  PIN o_ranQ[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -194.965 94.875 -192.755 95.055 ;
        RECT -194.965 94.795 -194.460 94.875 ;
        RECT -193.660 94.785 -192.755 94.875 ;
      LAYER mcon ;
        RECT -194.775 94.795 -194.605 94.965 ;
        RECT -193.410 94.795 -193.240 94.965 ;
      LAYER met1 ;
        RECT -194.660 95.060 -193.660 95.760 ;
        RECT -194.840 94.760 -193.150 95.060 ;
    END
  END o_ranQ[44]
  PIN o_ranQ[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -199.925 89.065 -199.420 89.145 ;
        RECT -198.620 89.065 -197.715 89.155 ;
        RECT -199.925 88.885 -197.715 89.065 ;
      LAYER mcon ;
        RECT -199.735 88.975 -199.565 89.145 ;
        RECT -198.370 88.975 -198.200 89.145 ;
      LAYER met1 ;
        RECT -199.800 88.880 -198.110 89.180 ;
        RECT -199.620 88.180 -198.620 88.880 ;
    END
  END o_ranQ[45]
  PIN o_ranQ[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -204.885 94.875 -202.675 95.055 ;
        RECT -204.885 94.795 -204.380 94.875 ;
        RECT -203.580 94.785 -202.675 94.875 ;
      LAYER mcon ;
        RECT -204.695 94.795 -204.525 94.965 ;
        RECT -203.330 94.795 -203.160 94.965 ;
      LAYER met1 ;
        RECT -204.580 95.060 -203.580 95.760 ;
        RECT -204.760 94.760 -203.070 95.060 ;
    END
  END o_ranQ[46]
  PIN o_ranQ[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -209.845 89.065 -209.340 89.145 ;
        RECT -208.540 89.065 -207.635 89.155 ;
        RECT -209.845 88.885 -207.635 89.065 ;
      LAYER mcon ;
        RECT -209.655 88.975 -209.485 89.145 ;
        RECT -208.290 88.975 -208.120 89.145 ;
      LAYER met1 ;
        RECT -209.720 88.880 -208.030 89.180 ;
        RECT -209.540 88.180 -208.540 88.880 ;
    END
  END o_ranQ[47]
  PIN o_ranQ[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -219.765 89.065 -219.260 89.145 ;
        RECT -218.460 89.065 -217.555 89.155 ;
        RECT -219.765 88.885 -217.555 89.065 ;
      LAYER mcon ;
        RECT -219.575 88.975 -219.405 89.145 ;
        RECT -218.210 88.975 -218.040 89.145 ;
      LAYER met1 ;
        RECT -219.640 88.880 -217.950 89.180 ;
        RECT -219.460 88.180 -218.460 88.880 ;
    END
  END o_ranQ[49]
  PIN o_ranQ[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -224.725 94.875 -222.515 95.055 ;
        RECT -224.725 94.795 -224.220 94.875 ;
        RECT -223.420 94.785 -222.515 94.875 ;
      LAYER mcon ;
        RECT -224.535 94.795 -224.365 94.965 ;
        RECT -223.170 94.795 -223.000 94.965 ;
      LAYER met1 ;
        RECT -224.420 95.060 -223.420 95.760 ;
        RECT -224.600 94.760 -222.910 95.060 ;
    END
  END o_ranQ[50]
  PIN o_ranQ[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -229.685 89.065 -229.180 89.145 ;
        RECT -228.380 89.065 -227.475 89.155 ;
        RECT -229.685 88.885 -227.475 89.065 ;
      LAYER mcon ;
        RECT -229.495 88.975 -229.325 89.145 ;
        RECT -228.130 88.975 -227.960 89.145 ;
      LAYER met1 ;
        RECT -229.560 88.880 -227.870 89.180 ;
        RECT -229.380 88.180 -228.380 88.880 ;
    END
  END o_ranQ[51]
  PIN o_ranQ[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -214.805 94.875 -212.595 95.055 ;
        RECT -214.805 94.795 -214.300 94.875 ;
        RECT -213.500 94.785 -212.595 94.875 ;
      LAYER mcon ;
        RECT -214.615 94.795 -214.445 94.965 ;
        RECT -213.250 94.795 -213.080 94.965 ;
      LAYER met1 ;
        RECT -214.500 95.060 -213.500 95.760 ;
        RECT -214.680 94.760 -212.990 95.060 ;
    END
  END o_ranQ[48]
  PIN o_ranQ[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -234.645 94.875 -232.435 95.055 ;
        RECT -234.645 94.795 -234.140 94.875 ;
        RECT -233.340 94.785 -232.435 94.875 ;
      LAYER mcon ;
        RECT -234.455 94.795 -234.285 94.965 ;
        RECT -233.090 94.795 -232.920 94.965 ;
      LAYER met1 ;
        RECT -234.340 95.060 -233.340 95.760 ;
        RECT -234.520 94.760 -232.830 95.060 ;
    END
  END o_ranQ[52]
  PIN o_ranQ[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -239.605 89.065 -239.100 89.145 ;
        RECT -238.300 89.065 -237.395 89.155 ;
        RECT -239.605 88.885 -237.395 89.065 ;
      LAYER mcon ;
        RECT -239.415 88.975 -239.245 89.145 ;
        RECT -238.050 88.975 -237.880 89.145 ;
      LAYER met1 ;
        RECT -239.480 88.880 -237.790 89.180 ;
        RECT -239.300 88.180 -238.300 88.880 ;
    END
  END o_ranQ[53]
  PIN o_ranQ[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -244.565 94.875 -242.355 95.055 ;
        RECT -244.565 94.795 -244.060 94.875 ;
        RECT -243.260 94.785 -242.355 94.875 ;
      LAYER mcon ;
        RECT -244.375 94.795 -244.205 94.965 ;
        RECT -243.010 94.795 -242.840 94.965 ;
      LAYER met1 ;
        RECT -244.260 95.060 -243.260 95.760 ;
        RECT -244.440 94.760 -242.750 95.060 ;
    END
  END o_ranQ[54]
  PIN o_ranQ[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -249.525 89.065 -249.020 89.145 ;
        RECT -248.220 89.065 -247.315 89.155 ;
        RECT -249.525 88.885 -247.315 89.065 ;
      LAYER mcon ;
        RECT -249.335 88.975 -249.165 89.145 ;
        RECT -247.970 88.975 -247.800 89.145 ;
      LAYER met1 ;
        RECT -249.400 88.880 -247.710 89.180 ;
        RECT -249.220 88.180 -248.220 88.880 ;
    END
  END o_ranQ[55]
  PIN o_ranQ[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -254.485 94.875 -252.275 95.055 ;
        RECT -254.485 94.795 -253.980 94.875 ;
        RECT -253.180 94.785 -252.275 94.875 ;
      LAYER mcon ;
        RECT -254.295 94.795 -254.125 94.965 ;
        RECT -252.930 94.795 -252.760 94.965 ;
      LAYER met1 ;
        RECT -254.180 95.060 -253.180 95.760 ;
        RECT -254.360 94.760 -252.670 95.060 ;
    END
  END o_ranQ[56]
  PIN o_ranQ[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -259.445 89.065 -258.940 89.145 ;
        RECT -258.140 89.065 -257.235 89.155 ;
        RECT -259.445 88.885 -257.235 89.065 ;
      LAYER mcon ;
        RECT -259.255 88.975 -259.085 89.145 ;
        RECT -257.890 88.975 -257.720 89.145 ;
      LAYER met1 ;
        RECT -259.320 88.880 -257.630 89.180 ;
        RECT -259.140 88.180 -258.140 88.880 ;
    END
  END o_ranQ[57]
  PIN o_ranQ[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -264.405 94.875 -262.195 95.055 ;
        RECT -264.405 94.795 -263.900 94.875 ;
        RECT -263.100 94.785 -262.195 94.875 ;
      LAYER mcon ;
        RECT -264.215 94.795 -264.045 94.965 ;
        RECT -262.850 94.795 -262.680 94.965 ;
      LAYER met1 ;
        RECT -264.100 95.060 -263.100 95.760 ;
        RECT -264.280 94.760 -262.590 95.060 ;
    END
  END o_ranQ[58]
  PIN o_ranQ[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -269.365 89.065 -268.860 89.145 ;
        RECT -268.060 89.065 -267.155 89.155 ;
        RECT -269.365 88.885 -267.155 89.065 ;
      LAYER mcon ;
        RECT -269.175 88.975 -269.005 89.145 ;
        RECT -267.810 88.975 -267.640 89.145 ;
      LAYER met1 ;
        RECT -269.240 88.880 -267.550 89.180 ;
        RECT -269.060 88.180 -268.060 88.880 ;
    END
  END o_ranQ[59]
  PIN o_ranQ[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -274.325 94.875 -272.115 95.055 ;
        RECT -274.325 94.795 -273.820 94.875 ;
        RECT -273.020 94.785 -272.115 94.875 ;
      LAYER mcon ;
        RECT -274.135 94.795 -273.965 94.965 ;
        RECT -272.770 94.795 -272.600 94.965 ;
      LAYER met1 ;
        RECT -274.020 95.060 -273.020 95.760 ;
        RECT -274.200 94.760 -272.510 95.060 ;
    END
  END o_ranQ[60]
  PIN o_ranQ[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -279.285 89.065 -278.780 89.145 ;
        RECT -277.980 89.065 -277.075 89.155 ;
        RECT -279.285 88.885 -277.075 89.065 ;
      LAYER mcon ;
        RECT -279.095 88.975 -278.925 89.145 ;
        RECT -277.730 88.975 -277.560 89.145 ;
      LAYER met1 ;
        RECT -279.160 88.880 -277.470 89.180 ;
        RECT -278.980 88.180 -277.980 88.880 ;
    END
  END o_ranQ[61]
  PIN o_ranQ[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -284.245 94.875 -282.035 95.055 ;
        RECT -284.245 94.795 -283.740 94.875 ;
        RECT -282.940 94.785 -282.035 94.875 ;
      LAYER mcon ;
        RECT -284.055 94.795 -283.885 94.965 ;
        RECT -282.690 94.795 -282.520 94.965 ;
      LAYER met1 ;
        RECT -283.940 95.060 -282.940 95.760 ;
        RECT -284.120 94.760 -282.430 95.060 ;
    END
  END o_ranQ[62]
  PIN o_ranQ[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -289.205 89.065 -288.700 89.145 ;
        RECT -287.900 89.065 -286.995 89.155 ;
        RECT -289.205 88.885 -286.995 89.065 ;
      LAYER mcon ;
        RECT -289.015 88.975 -288.845 89.145 ;
        RECT -287.650 88.975 -287.480 89.145 ;
      LAYER met1 ;
        RECT -289.080 88.880 -287.390 89.180 ;
        RECT -288.900 88.180 -287.900 88.880 ;
    END
  END o_ranQ[63]
  PIN i_srclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 31.679998 ;
    PORT
      LAYER li1 ;
        RECT -290.905 92.005 -290.570 92.275 ;
        RECT -281.970 92.005 -281.635 92.275 ;
        RECT -280.985 92.005 -280.650 92.275 ;
        RECT -272.050 92.005 -271.715 92.275 ;
        RECT -271.065 92.005 -270.730 92.275 ;
        RECT -262.130 92.005 -261.795 92.275 ;
        RECT -261.145 92.005 -260.810 92.275 ;
        RECT -252.210 92.005 -251.875 92.275 ;
        RECT -251.225 92.005 -250.890 92.275 ;
        RECT -242.290 92.005 -241.955 92.275 ;
        RECT -241.305 92.005 -240.970 92.275 ;
        RECT -232.370 92.005 -232.035 92.275 ;
        RECT -231.385 92.005 -231.050 92.275 ;
        RECT -222.450 92.005 -222.115 92.275 ;
        RECT -221.465 92.005 -221.130 92.275 ;
        RECT -212.530 92.005 -212.195 92.275 ;
        RECT -211.545 92.005 -211.210 92.275 ;
        RECT -202.610 92.005 -202.275 92.275 ;
        RECT -201.625 92.005 -201.290 92.275 ;
        RECT -192.690 92.005 -192.355 92.275 ;
        RECT -191.705 92.005 -191.370 92.275 ;
        RECT -182.770 92.005 -182.435 92.275 ;
        RECT -181.785 92.005 -181.450 92.275 ;
        RECT -172.850 92.005 -172.515 92.275 ;
        RECT -171.865 92.005 -171.530 92.275 ;
        RECT -162.930 92.005 -162.595 92.275 ;
        RECT -161.945 92.005 -161.610 92.275 ;
        RECT -153.010 92.005 -152.675 92.275 ;
        RECT -152.025 92.005 -151.690 92.275 ;
        RECT -143.090 92.005 -142.755 92.275 ;
        RECT -142.105 92.005 -141.770 92.275 ;
        RECT -133.170 92.005 -132.835 92.275 ;
        RECT -132.185 92.005 -131.850 92.275 ;
        RECT -123.250 92.005 -122.915 92.275 ;
        RECT -122.265 92.005 -121.930 92.275 ;
        RECT -113.330 92.005 -112.995 92.275 ;
        RECT -112.345 92.005 -112.010 92.275 ;
        RECT -103.410 92.005 -103.075 92.275 ;
        RECT -102.425 92.005 -102.090 92.275 ;
        RECT -93.490 92.005 -93.155 92.275 ;
        RECT -92.505 92.005 -92.170 92.275 ;
        RECT -83.570 92.005 -83.235 92.275 ;
        RECT -82.585 92.005 -82.250 92.275 ;
        RECT -73.650 92.005 -73.315 92.275 ;
        RECT -72.665 92.005 -72.330 92.275 ;
        RECT -63.730 92.005 -63.395 92.275 ;
        RECT -62.745 92.005 -62.410 92.275 ;
        RECT -53.810 92.005 -53.475 92.275 ;
        RECT -52.825 92.005 -52.490 92.275 ;
        RECT -43.890 92.005 -43.555 92.275 ;
        RECT -42.905 92.005 -42.570 92.275 ;
        RECT -33.970 92.005 -33.635 92.275 ;
        RECT -32.985 92.005 -32.650 92.275 ;
        RECT -24.050 92.005 -23.715 92.275 ;
        RECT -23.065 92.005 -22.730 92.275 ;
        RECT -14.130 92.005 -13.795 92.275 ;
        RECT -13.145 92.005 -12.810 92.275 ;
        RECT -4.210 92.005 -3.875 92.275 ;
        RECT -3.225 92.005 -2.890 92.275 ;
        RECT 5.710 92.005 6.045 92.275 ;
        RECT 6.695 92.005 7.030 92.275 ;
        RECT 15.630 92.005 15.965 92.275 ;
        RECT 16.615 92.005 16.950 92.275 ;
        RECT 25.550 92.005 25.885 92.275 ;
        RECT -286.930 91.665 -286.595 91.935 ;
        RECT -285.945 91.665 -285.610 91.935 ;
        RECT -277.010 91.665 -276.675 91.935 ;
        RECT -276.025 91.665 -275.690 91.935 ;
        RECT -267.090 91.665 -266.755 91.935 ;
        RECT -266.105 91.665 -265.770 91.935 ;
        RECT -257.170 91.665 -256.835 91.935 ;
        RECT -256.185 91.665 -255.850 91.935 ;
        RECT -247.250 91.665 -246.915 91.935 ;
        RECT -246.265 91.665 -245.930 91.935 ;
        RECT -237.330 91.665 -236.995 91.935 ;
        RECT -236.345 91.665 -236.010 91.935 ;
        RECT -227.410 91.665 -227.075 91.935 ;
        RECT -226.425 91.665 -226.090 91.935 ;
        RECT -217.490 91.665 -217.155 91.935 ;
        RECT -216.505 91.665 -216.170 91.935 ;
        RECT -207.570 91.665 -207.235 91.935 ;
        RECT -206.585 91.665 -206.250 91.935 ;
        RECT -197.650 91.665 -197.315 91.935 ;
        RECT -196.665 91.665 -196.330 91.935 ;
        RECT -187.730 91.665 -187.395 91.935 ;
        RECT -186.745 91.665 -186.410 91.935 ;
        RECT -177.810 91.665 -177.475 91.935 ;
        RECT -176.825 91.665 -176.490 91.935 ;
        RECT -167.890 91.665 -167.555 91.935 ;
        RECT -166.905 91.665 -166.570 91.935 ;
        RECT -157.970 91.665 -157.635 91.935 ;
        RECT -156.985 91.665 -156.650 91.935 ;
        RECT -148.050 91.665 -147.715 91.935 ;
        RECT -147.065 91.665 -146.730 91.935 ;
        RECT -138.130 91.665 -137.795 91.935 ;
        RECT -137.145 91.665 -136.810 91.935 ;
        RECT -128.210 91.665 -127.875 91.935 ;
        RECT -127.225 91.665 -126.890 91.935 ;
        RECT -118.290 91.665 -117.955 91.935 ;
        RECT -117.305 91.665 -116.970 91.935 ;
        RECT -108.370 91.665 -108.035 91.935 ;
        RECT -107.385 91.665 -107.050 91.935 ;
        RECT -98.450 91.665 -98.115 91.935 ;
        RECT -97.465 91.665 -97.130 91.935 ;
        RECT -88.530 91.665 -88.195 91.935 ;
        RECT -87.545 91.665 -87.210 91.935 ;
        RECT -78.610 91.665 -78.275 91.935 ;
        RECT -77.625 91.665 -77.290 91.935 ;
        RECT -68.690 91.665 -68.355 91.935 ;
        RECT -67.705 91.665 -67.370 91.935 ;
        RECT -58.770 91.665 -58.435 91.935 ;
        RECT -57.785 91.665 -57.450 91.935 ;
        RECT -48.850 91.665 -48.515 91.935 ;
        RECT -47.865 91.665 -47.530 91.935 ;
        RECT -38.930 91.665 -38.595 91.935 ;
        RECT -37.945 91.665 -37.610 91.935 ;
        RECT -29.010 91.665 -28.675 91.935 ;
        RECT -28.025 91.665 -27.690 91.935 ;
        RECT -19.090 91.665 -18.755 91.935 ;
        RECT -18.105 91.665 -17.770 91.935 ;
        RECT -9.170 91.665 -8.835 91.935 ;
        RECT -8.185 91.665 -7.850 91.935 ;
        RECT 0.750 91.665 1.085 91.935 ;
        RECT 1.735 91.665 2.070 91.935 ;
        RECT 10.670 91.665 11.005 91.935 ;
        RECT 11.655 91.665 11.990 91.935 ;
        RECT 20.590 91.665 20.925 91.935 ;
        RECT 21.575 91.665 21.910 91.935 ;
      LAYER mcon ;
        RECT -290.820 92.085 -290.650 92.255 ;
        RECT -281.890 92.085 -281.720 92.255 ;
        RECT -280.900 92.085 -280.730 92.255 ;
        RECT -271.970 92.085 -271.800 92.255 ;
        RECT -270.980 92.085 -270.810 92.255 ;
        RECT -262.050 92.085 -261.880 92.255 ;
        RECT -261.060 92.085 -260.890 92.255 ;
        RECT -252.130 92.085 -251.960 92.255 ;
        RECT -251.140 92.085 -250.970 92.255 ;
        RECT -242.210 92.085 -242.040 92.255 ;
        RECT -241.220 92.085 -241.050 92.255 ;
        RECT -232.290 92.085 -232.120 92.255 ;
        RECT -231.300 92.085 -231.130 92.255 ;
        RECT -222.370 92.085 -222.200 92.255 ;
        RECT -221.380 92.085 -221.210 92.255 ;
        RECT -212.450 92.085 -212.280 92.255 ;
        RECT -211.460 92.085 -211.290 92.255 ;
        RECT -202.530 92.085 -202.360 92.255 ;
        RECT -201.540 92.085 -201.370 92.255 ;
        RECT -192.610 92.085 -192.440 92.255 ;
        RECT -191.620 92.085 -191.450 92.255 ;
        RECT -182.690 92.085 -182.520 92.255 ;
        RECT -181.700 92.085 -181.530 92.255 ;
        RECT -172.770 92.085 -172.600 92.255 ;
        RECT -171.780 92.085 -171.610 92.255 ;
        RECT -162.850 92.085 -162.680 92.255 ;
        RECT -161.860 92.085 -161.690 92.255 ;
        RECT -152.930 92.085 -152.760 92.255 ;
        RECT -151.940 92.085 -151.770 92.255 ;
        RECT -143.010 92.085 -142.840 92.255 ;
        RECT -142.020 92.085 -141.850 92.255 ;
        RECT -133.090 92.085 -132.920 92.255 ;
        RECT -132.100 92.085 -131.930 92.255 ;
        RECT -123.170 92.085 -123.000 92.255 ;
        RECT -122.180 92.085 -122.010 92.255 ;
        RECT -113.250 92.085 -113.080 92.255 ;
        RECT -112.260 92.085 -112.090 92.255 ;
        RECT -103.330 92.085 -103.160 92.255 ;
        RECT -102.340 92.085 -102.170 92.255 ;
        RECT -93.410 92.085 -93.240 92.255 ;
        RECT -92.420 92.085 -92.250 92.255 ;
        RECT -83.490 92.085 -83.320 92.255 ;
        RECT -82.500 92.085 -82.330 92.255 ;
        RECT -73.570 92.085 -73.400 92.255 ;
        RECT -72.580 92.085 -72.410 92.255 ;
        RECT -63.650 92.085 -63.480 92.255 ;
        RECT -62.660 92.085 -62.490 92.255 ;
        RECT -53.730 92.085 -53.560 92.255 ;
        RECT -52.740 92.085 -52.570 92.255 ;
        RECT -43.810 92.085 -43.640 92.255 ;
        RECT -42.820 92.085 -42.650 92.255 ;
        RECT -33.890 92.085 -33.720 92.255 ;
        RECT -32.900 92.085 -32.730 92.255 ;
        RECT -23.970 92.085 -23.800 92.255 ;
        RECT -22.980 92.085 -22.810 92.255 ;
        RECT -14.050 92.085 -13.880 92.255 ;
        RECT -13.060 92.085 -12.890 92.255 ;
        RECT -4.130 92.085 -3.960 92.255 ;
        RECT -3.140 92.085 -2.970 92.255 ;
        RECT 5.790 92.085 5.960 92.255 ;
        RECT 6.780 92.085 6.950 92.255 ;
        RECT 15.710 92.085 15.880 92.255 ;
        RECT 16.700 92.085 16.870 92.255 ;
        RECT 25.630 92.085 25.800 92.255 ;
        RECT -286.850 91.685 -286.680 91.855 ;
        RECT -285.860 91.685 -285.690 91.855 ;
        RECT -276.930 91.685 -276.760 91.855 ;
        RECT -275.940 91.685 -275.770 91.855 ;
        RECT -267.010 91.685 -266.840 91.855 ;
        RECT -266.020 91.685 -265.850 91.855 ;
        RECT -257.090 91.685 -256.920 91.855 ;
        RECT -256.100 91.685 -255.930 91.855 ;
        RECT -247.170 91.685 -247.000 91.855 ;
        RECT -246.180 91.685 -246.010 91.855 ;
        RECT -237.250 91.685 -237.080 91.855 ;
        RECT -236.260 91.685 -236.090 91.855 ;
        RECT -227.330 91.685 -227.160 91.855 ;
        RECT -226.340 91.685 -226.170 91.855 ;
        RECT -217.410 91.685 -217.240 91.855 ;
        RECT -216.420 91.685 -216.250 91.855 ;
        RECT -207.490 91.685 -207.320 91.855 ;
        RECT -206.500 91.685 -206.330 91.855 ;
        RECT -197.570 91.685 -197.400 91.855 ;
        RECT -196.580 91.685 -196.410 91.855 ;
        RECT -187.650 91.685 -187.480 91.855 ;
        RECT -186.660 91.685 -186.490 91.855 ;
        RECT -177.730 91.685 -177.560 91.855 ;
        RECT -176.740 91.685 -176.570 91.855 ;
        RECT -167.810 91.685 -167.640 91.855 ;
        RECT -166.820 91.685 -166.650 91.855 ;
        RECT -157.890 91.685 -157.720 91.855 ;
        RECT -156.900 91.685 -156.730 91.855 ;
        RECT -147.970 91.685 -147.800 91.855 ;
        RECT -146.980 91.685 -146.810 91.855 ;
        RECT -138.050 91.685 -137.880 91.855 ;
        RECT -137.060 91.685 -136.890 91.855 ;
        RECT -128.130 91.685 -127.960 91.855 ;
        RECT -127.140 91.685 -126.970 91.855 ;
        RECT -118.210 91.685 -118.040 91.855 ;
        RECT -117.220 91.685 -117.050 91.855 ;
        RECT -108.290 91.685 -108.120 91.855 ;
        RECT -107.300 91.685 -107.130 91.855 ;
        RECT -98.370 91.685 -98.200 91.855 ;
        RECT -97.380 91.685 -97.210 91.855 ;
        RECT -88.450 91.685 -88.280 91.855 ;
        RECT -87.460 91.685 -87.290 91.855 ;
        RECT -78.530 91.685 -78.360 91.855 ;
        RECT -77.540 91.685 -77.370 91.855 ;
        RECT -68.610 91.685 -68.440 91.855 ;
        RECT -67.620 91.685 -67.450 91.855 ;
        RECT -58.690 91.685 -58.520 91.855 ;
        RECT -57.700 91.685 -57.530 91.855 ;
        RECT -48.770 91.685 -48.600 91.855 ;
        RECT -47.780 91.685 -47.610 91.855 ;
        RECT -38.850 91.685 -38.680 91.855 ;
        RECT -37.860 91.685 -37.690 91.855 ;
        RECT -28.930 91.685 -28.760 91.855 ;
        RECT -27.940 91.685 -27.770 91.855 ;
        RECT -19.010 91.685 -18.840 91.855 ;
        RECT -18.020 91.685 -17.850 91.855 ;
        RECT -9.090 91.685 -8.920 91.855 ;
        RECT -8.100 91.685 -7.930 91.855 ;
        RECT 0.830 91.685 1.000 91.855 ;
        RECT 1.820 91.685 1.990 91.855 ;
        RECT 10.750 91.685 10.920 91.855 ;
        RECT 11.740 91.685 11.910 91.855 ;
        RECT 20.670 91.685 20.840 91.855 ;
        RECT 21.660 91.685 21.830 91.855 ;
      LAYER met1 ;
        RECT -291.010 91.900 -290.550 92.350 ;
        RECT -286.950 91.590 -286.490 92.040 ;
        RECT -286.050 91.590 -285.590 92.040 ;
        RECT -281.990 91.900 -281.530 92.350 ;
        RECT -281.090 91.900 -280.630 92.350 ;
        RECT -277.030 91.590 -276.570 92.040 ;
        RECT -276.130 91.590 -275.670 92.040 ;
        RECT -272.070 91.900 -271.610 92.350 ;
        RECT -271.170 91.900 -270.710 92.350 ;
        RECT -267.110 91.590 -266.650 92.040 ;
        RECT -266.210 91.590 -265.750 92.040 ;
        RECT -262.150 91.900 -261.690 92.350 ;
        RECT -261.250 91.900 -260.790 92.350 ;
        RECT -257.190 91.590 -256.730 92.040 ;
        RECT -256.290 91.590 -255.830 92.040 ;
        RECT -252.230 91.900 -251.770 92.350 ;
        RECT -251.330 91.900 -250.870 92.350 ;
        RECT -247.270 91.590 -246.810 92.040 ;
        RECT -246.370 91.590 -245.910 92.040 ;
        RECT -242.310 91.900 -241.850 92.350 ;
        RECT -241.410 91.900 -240.950 92.350 ;
        RECT -237.350 91.590 -236.890 92.040 ;
        RECT -236.450 91.590 -235.990 92.040 ;
        RECT -232.390 91.900 -231.930 92.350 ;
        RECT -231.490 91.900 -231.030 92.350 ;
        RECT -227.430 91.590 -226.970 92.040 ;
        RECT -226.530 91.590 -226.070 92.040 ;
        RECT -222.470 91.900 -222.010 92.350 ;
        RECT -221.570 91.900 -221.110 92.350 ;
        RECT -217.510 91.590 -217.050 92.040 ;
        RECT -216.610 91.590 -216.150 92.040 ;
        RECT -212.550 91.900 -212.090 92.350 ;
        RECT -211.650 91.900 -211.190 92.350 ;
        RECT -207.590 91.590 -207.130 92.040 ;
        RECT -206.690 91.590 -206.230 92.040 ;
        RECT -202.630 91.900 -202.170 92.350 ;
        RECT -201.730 91.900 -201.270 92.350 ;
        RECT -197.670 91.590 -197.210 92.040 ;
        RECT -196.770 91.590 -196.310 92.040 ;
        RECT -192.710 91.900 -192.250 92.350 ;
        RECT -191.810 91.900 -191.350 92.350 ;
        RECT -187.750 91.590 -187.290 92.040 ;
        RECT -186.850 91.590 -186.390 92.040 ;
        RECT -182.790 91.900 -182.330 92.350 ;
        RECT -181.890 91.900 -181.430 92.350 ;
        RECT -177.830 91.590 -177.370 92.040 ;
        RECT -176.930 91.590 -176.470 92.040 ;
        RECT -172.870 91.900 -172.410 92.350 ;
        RECT -171.970 91.900 -171.510 92.350 ;
        RECT -167.910 91.590 -167.450 92.040 ;
        RECT -167.010 91.590 -166.550 92.040 ;
        RECT -162.950 91.900 -162.490 92.350 ;
        RECT -162.050 91.900 -161.590 92.350 ;
        RECT -157.990 91.590 -157.530 92.040 ;
        RECT -157.090 91.590 -156.630 92.040 ;
        RECT -153.030 91.900 -152.570 92.350 ;
        RECT -152.130 91.900 -151.670 92.350 ;
        RECT -148.070 91.590 -147.610 92.040 ;
        RECT -147.170 91.590 -146.710 92.040 ;
        RECT -143.110 91.900 -142.650 92.350 ;
        RECT -142.210 91.900 -141.750 92.350 ;
        RECT -138.150 91.590 -137.690 92.040 ;
        RECT -137.250 91.590 -136.790 92.040 ;
        RECT -133.190 91.900 -132.730 92.350 ;
        RECT -132.290 91.900 -131.830 92.350 ;
        RECT -128.230 91.590 -127.770 92.040 ;
        RECT -127.330 91.590 -126.870 92.040 ;
        RECT -123.270 91.900 -122.810 92.350 ;
        RECT -122.370 91.900 -121.910 92.350 ;
        RECT -118.310 91.590 -117.850 92.040 ;
        RECT -117.410 91.590 -116.950 92.040 ;
        RECT -113.350 91.900 -112.890 92.350 ;
        RECT -112.450 91.900 -111.990 92.350 ;
        RECT -108.390 91.590 -107.930 92.040 ;
        RECT -107.490 91.590 -107.030 92.040 ;
        RECT -103.430 91.900 -102.970 92.350 ;
        RECT -102.530 91.900 -102.070 92.350 ;
        RECT -98.470 91.590 -98.010 92.040 ;
        RECT -97.570 91.590 -97.110 92.040 ;
        RECT -93.510 91.900 -93.050 92.350 ;
        RECT -92.610 91.900 -92.150 92.350 ;
        RECT -88.550 91.590 -88.090 92.040 ;
        RECT -87.650 91.590 -87.190 92.040 ;
        RECT -83.590 91.900 -83.130 92.350 ;
        RECT -82.690 91.900 -82.230 92.350 ;
        RECT -78.630 91.590 -78.170 92.040 ;
        RECT -77.730 91.590 -77.270 92.040 ;
        RECT -73.670 91.900 -73.210 92.350 ;
        RECT -72.770 91.900 -72.310 92.350 ;
        RECT -68.710 91.590 -68.250 92.040 ;
        RECT -67.810 91.590 -67.350 92.040 ;
        RECT -63.750 91.900 -63.290 92.350 ;
        RECT -62.850 91.900 -62.390 92.350 ;
        RECT -58.790 91.590 -58.330 92.040 ;
        RECT -57.890 91.590 -57.430 92.040 ;
        RECT -53.830 91.900 -53.370 92.350 ;
        RECT -52.930 91.900 -52.470 92.350 ;
        RECT -48.870 91.590 -48.410 92.040 ;
        RECT -47.970 91.590 -47.510 92.040 ;
        RECT -43.910 91.900 -43.450 92.350 ;
        RECT -43.010 91.900 -42.550 92.350 ;
        RECT -38.950 91.590 -38.490 92.040 ;
        RECT -38.050 91.590 -37.590 92.040 ;
        RECT -33.990 91.900 -33.530 92.350 ;
        RECT -33.090 91.900 -32.630 92.350 ;
        RECT -29.030 91.590 -28.570 92.040 ;
        RECT -28.130 91.590 -27.670 92.040 ;
        RECT -24.070 91.900 -23.610 92.350 ;
        RECT -23.170 91.900 -22.710 92.350 ;
        RECT -19.110 91.590 -18.650 92.040 ;
        RECT -18.210 91.590 -17.750 92.040 ;
        RECT -14.150 91.900 -13.690 92.350 ;
        RECT -13.250 91.900 -12.790 92.350 ;
        RECT -9.190 91.590 -8.730 92.040 ;
        RECT -8.290 91.590 -7.830 92.040 ;
        RECT -4.230 91.900 -3.770 92.350 ;
        RECT -3.330 91.900 -2.870 92.350 ;
        RECT 0.730 91.590 1.190 92.040 ;
        RECT 1.630 91.590 2.090 92.040 ;
        RECT 5.690 91.900 6.150 92.350 ;
        RECT 6.590 91.900 7.050 92.350 ;
        RECT 10.650 91.590 11.110 92.040 ;
        RECT 11.550 91.590 12.010 92.040 ;
        RECT 15.610 91.900 16.070 92.350 ;
        RECT 16.510 91.900 16.970 92.350 ;
        RECT 20.570 91.590 21.030 92.040 ;
        RECT 21.470 91.590 21.930 92.040 ;
        RECT 25.530 91.900 25.990 92.350 ;
      LAYER via ;
        RECT -290.940 92.000 -290.640 92.300 ;
        RECT -286.860 91.640 -286.560 91.940 ;
        RECT -285.980 91.640 -285.680 91.940 ;
        RECT -281.900 92.000 -281.600 92.300 ;
        RECT -281.020 92.000 -280.720 92.300 ;
        RECT -276.940 91.640 -276.640 91.940 ;
        RECT -276.060 91.640 -275.760 91.940 ;
        RECT -271.980 92.000 -271.680 92.300 ;
        RECT -271.100 92.000 -270.800 92.300 ;
        RECT -267.020 91.640 -266.720 91.940 ;
        RECT -266.140 91.640 -265.840 91.940 ;
        RECT -262.060 92.000 -261.760 92.300 ;
        RECT -261.180 92.000 -260.880 92.300 ;
        RECT -257.100 91.640 -256.800 91.940 ;
        RECT -256.220 91.640 -255.920 91.940 ;
        RECT -252.140 92.000 -251.840 92.300 ;
        RECT -251.260 92.000 -250.960 92.300 ;
        RECT -247.180 91.640 -246.880 91.940 ;
        RECT -246.300 91.640 -246.000 91.940 ;
        RECT -242.220 92.000 -241.920 92.300 ;
        RECT -241.340 92.000 -241.040 92.300 ;
        RECT -237.260 91.640 -236.960 91.940 ;
        RECT -236.380 91.640 -236.080 91.940 ;
        RECT -232.300 92.000 -232.000 92.300 ;
        RECT -231.420 92.000 -231.120 92.300 ;
        RECT -227.340 91.640 -227.040 91.940 ;
        RECT -226.460 91.640 -226.160 91.940 ;
        RECT -222.380 92.000 -222.080 92.300 ;
        RECT -221.500 92.000 -221.200 92.300 ;
        RECT -217.420 91.640 -217.120 91.940 ;
        RECT -216.540 91.640 -216.240 91.940 ;
        RECT -212.460 92.000 -212.160 92.300 ;
        RECT -211.580 92.000 -211.280 92.300 ;
        RECT -207.500 91.640 -207.200 91.940 ;
        RECT -206.620 91.640 -206.320 91.940 ;
        RECT -202.540 92.000 -202.240 92.300 ;
        RECT -201.660 92.000 -201.360 92.300 ;
        RECT -197.580 91.640 -197.280 91.940 ;
        RECT -196.700 91.640 -196.400 91.940 ;
        RECT -192.620 92.000 -192.320 92.300 ;
        RECT -191.740 92.000 -191.440 92.300 ;
        RECT -187.660 91.640 -187.360 91.940 ;
        RECT -186.780 91.640 -186.480 91.940 ;
        RECT -182.700 92.000 -182.400 92.300 ;
        RECT -181.820 92.000 -181.520 92.300 ;
        RECT -177.740 91.640 -177.440 91.940 ;
        RECT -176.860 91.640 -176.560 91.940 ;
        RECT -172.780 92.000 -172.480 92.300 ;
        RECT -171.900 92.000 -171.600 92.300 ;
        RECT -167.820 91.640 -167.520 91.940 ;
        RECT -166.940 91.640 -166.640 91.940 ;
        RECT -162.860 92.000 -162.560 92.300 ;
        RECT -161.980 92.000 -161.680 92.300 ;
        RECT -157.900 91.640 -157.600 91.940 ;
        RECT -157.020 91.640 -156.720 91.940 ;
        RECT -152.940 92.000 -152.640 92.300 ;
        RECT -152.060 92.000 -151.760 92.300 ;
        RECT -147.980 91.640 -147.680 91.940 ;
        RECT -147.100 91.640 -146.800 91.940 ;
        RECT -143.020 92.000 -142.720 92.300 ;
        RECT -142.140 92.000 -141.840 92.300 ;
        RECT -138.060 91.640 -137.760 91.940 ;
        RECT -137.180 91.640 -136.880 91.940 ;
        RECT -133.100 92.000 -132.800 92.300 ;
        RECT -132.220 92.000 -131.920 92.300 ;
        RECT -128.140 91.640 -127.840 91.940 ;
        RECT -127.260 91.640 -126.960 91.940 ;
        RECT -123.180 92.000 -122.880 92.300 ;
        RECT -122.300 92.000 -122.000 92.300 ;
        RECT -118.220 91.640 -117.920 91.940 ;
        RECT -117.340 91.640 -117.040 91.940 ;
        RECT -113.260 92.000 -112.960 92.300 ;
        RECT -112.380 92.000 -112.080 92.300 ;
        RECT -108.300 91.640 -108.000 91.940 ;
        RECT -107.420 91.640 -107.120 91.940 ;
        RECT -103.340 92.000 -103.040 92.300 ;
        RECT -102.460 92.000 -102.160 92.300 ;
        RECT -98.380 91.640 -98.080 91.940 ;
        RECT -97.500 91.640 -97.200 91.940 ;
        RECT -93.420 92.000 -93.120 92.300 ;
        RECT -92.540 92.000 -92.240 92.300 ;
        RECT -88.460 91.640 -88.160 91.940 ;
        RECT -87.580 91.640 -87.280 91.940 ;
        RECT -83.500 92.000 -83.200 92.300 ;
        RECT -82.620 92.000 -82.320 92.300 ;
        RECT -78.540 91.640 -78.240 91.940 ;
        RECT -77.660 91.640 -77.360 91.940 ;
        RECT -73.580 92.000 -73.280 92.300 ;
        RECT -72.700 92.000 -72.400 92.300 ;
        RECT -68.620 91.640 -68.320 91.940 ;
        RECT -67.740 91.640 -67.440 91.940 ;
        RECT -63.660 92.000 -63.360 92.300 ;
        RECT -62.780 92.000 -62.480 92.300 ;
        RECT -58.700 91.640 -58.400 91.940 ;
        RECT -57.820 91.640 -57.520 91.940 ;
        RECT -53.740 92.000 -53.440 92.300 ;
        RECT -52.860 92.000 -52.560 92.300 ;
        RECT -48.780 91.640 -48.480 91.940 ;
        RECT -47.900 91.640 -47.600 91.940 ;
        RECT -43.820 92.000 -43.520 92.300 ;
        RECT -42.940 92.000 -42.640 92.300 ;
        RECT -38.860 91.640 -38.560 91.940 ;
        RECT -37.980 91.640 -37.680 91.940 ;
        RECT -33.900 92.000 -33.600 92.300 ;
        RECT -33.020 92.000 -32.720 92.300 ;
        RECT -28.940 91.640 -28.640 91.940 ;
        RECT -28.060 91.640 -27.760 91.940 ;
        RECT -23.980 92.000 -23.680 92.300 ;
        RECT -23.100 92.000 -22.800 92.300 ;
        RECT -19.020 91.640 -18.720 91.940 ;
        RECT -18.140 91.640 -17.840 91.940 ;
        RECT -14.060 92.000 -13.760 92.300 ;
        RECT -13.180 92.000 -12.880 92.300 ;
        RECT -9.100 91.640 -8.800 91.940 ;
        RECT -8.220 91.640 -7.920 91.940 ;
        RECT -4.140 92.000 -3.840 92.300 ;
        RECT -3.260 92.000 -2.960 92.300 ;
        RECT 0.820 91.640 1.120 91.940 ;
        RECT 1.700 91.640 2.000 91.940 ;
        RECT 5.780 92.000 6.080 92.300 ;
        RECT 6.660 92.000 6.960 92.300 ;
        RECT 10.740 91.640 11.040 91.940 ;
        RECT 11.620 91.640 11.920 91.940 ;
        RECT 15.700 92.000 16.000 92.300 ;
        RECT 16.580 92.000 16.880 92.300 ;
        RECT 20.660 91.640 20.960 91.940 ;
        RECT 21.540 91.640 21.840 91.940 ;
        RECT 25.620 92.000 25.920 92.300 ;
      LAYER met2 ;
        RECT -291.010 92.040 -290.550 92.350 ;
        RECT -288.820 92.040 -288.680 92.440 ;
        RECT -283.860 92.040 -283.720 92.440 ;
        RECT -281.990 92.040 -280.630 92.350 ;
        RECT -278.900 92.040 -278.760 92.440 ;
        RECT -273.940 92.040 -273.800 92.440 ;
        RECT -272.070 92.040 -270.710 92.350 ;
        RECT -268.980 92.040 -268.840 92.440 ;
        RECT -264.020 92.040 -263.880 92.440 ;
        RECT -262.150 92.040 -260.790 92.350 ;
        RECT -259.060 92.040 -258.920 92.440 ;
        RECT -254.100 92.040 -253.960 92.440 ;
        RECT -252.230 92.040 -250.870 92.350 ;
        RECT -249.140 92.040 -249.000 92.440 ;
        RECT -244.180 92.040 -244.040 92.440 ;
        RECT -242.310 92.040 -240.950 92.350 ;
        RECT -239.220 92.040 -239.080 92.440 ;
        RECT -234.260 92.040 -234.120 92.440 ;
        RECT -232.390 92.040 -231.030 92.350 ;
        RECT -229.300 92.040 -229.160 92.440 ;
        RECT -224.340 92.040 -224.200 92.440 ;
        RECT -222.470 92.040 -221.110 92.350 ;
        RECT -219.380 92.040 -219.240 92.440 ;
        RECT -214.420 92.040 -214.280 92.440 ;
        RECT -212.550 92.040 -211.190 92.350 ;
        RECT -209.460 92.040 -209.320 92.440 ;
        RECT -204.500 92.040 -204.360 92.440 ;
        RECT -202.630 92.040 -201.270 92.350 ;
        RECT -199.540 92.040 -199.400 92.440 ;
        RECT -194.580 92.040 -194.440 92.440 ;
        RECT -192.710 92.040 -191.350 92.350 ;
        RECT -189.620 92.040 -189.480 92.440 ;
        RECT -184.660 92.040 -184.520 92.440 ;
        RECT -182.790 92.040 -181.430 92.350 ;
        RECT -179.700 92.040 -179.560 92.440 ;
        RECT -174.740 92.040 -174.600 92.440 ;
        RECT -172.870 92.040 -171.510 92.350 ;
        RECT -169.780 92.040 -169.640 92.440 ;
        RECT -164.820 92.040 -164.680 92.440 ;
        RECT -162.950 92.040 -161.590 92.350 ;
        RECT -159.860 92.040 -159.720 92.440 ;
        RECT -154.900 92.040 -154.760 92.440 ;
        RECT -153.030 92.040 -151.670 92.350 ;
        RECT -149.940 92.040 -149.800 92.440 ;
        RECT -144.980 92.040 -144.840 92.440 ;
        RECT -143.110 92.040 -141.750 92.350 ;
        RECT -140.020 92.040 -139.880 92.440 ;
        RECT -135.060 92.040 -134.920 92.440 ;
        RECT -133.190 92.040 -131.830 92.350 ;
        RECT -130.100 92.040 -129.960 92.440 ;
        RECT -125.140 92.040 -125.000 92.440 ;
        RECT -123.270 92.040 -121.910 92.350 ;
        RECT -120.180 92.040 -120.040 92.440 ;
        RECT -115.220 92.040 -115.080 92.440 ;
        RECT -113.350 92.040 -111.990 92.350 ;
        RECT -110.260 92.040 -110.120 92.440 ;
        RECT -105.300 92.040 -105.160 92.440 ;
        RECT -103.430 92.040 -102.070 92.350 ;
        RECT -100.340 92.040 -100.200 92.440 ;
        RECT -95.380 92.040 -95.240 92.440 ;
        RECT -93.510 92.040 -92.150 92.350 ;
        RECT -90.420 92.040 -90.280 92.440 ;
        RECT -85.460 92.040 -85.320 92.440 ;
        RECT -83.590 92.040 -82.230 92.350 ;
        RECT -80.500 92.040 -80.360 92.440 ;
        RECT -75.540 92.040 -75.400 92.440 ;
        RECT -73.670 92.040 -72.310 92.350 ;
        RECT -70.580 92.040 -70.440 92.440 ;
        RECT -65.620 92.040 -65.480 92.440 ;
        RECT -63.750 92.040 -62.390 92.350 ;
        RECT -60.660 92.040 -60.520 92.440 ;
        RECT -55.700 92.040 -55.560 92.440 ;
        RECT -53.830 92.040 -52.470 92.350 ;
        RECT -50.740 92.040 -50.600 92.440 ;
        RECT -45.780 92.040 -45.640 92.440 ;
        RECT -43.910 92.040 -42.550 92.350 ;
        RECT -40.820 92.040 -40.680 92.440 ;
        RECT -35.860 92.040 -35.720 92.440 ;
        RECT -33.990 92.040 -32.630 92.350 ;
        RECT -30.900 92.040 -30.760 92.440 ;
        RECT -25.940 92.040 -25.800 92.440 ;
        RECT -24.070 92.040 -22.710 92.350 ;
        RECT -20.980 92.040 -20.840 92.440 ;
        RECT -16.020 92.040 -15.880 92.440 ;
        RECT -14.150 92.040 -12.790 92.350 ;
        RECT -11.060 92.040 -10.920 92.440 ;
        RECT -6.100 92.040 -5.960 92.440 ;
        RECT -4.230 92.040 -2.870 92.350 ;
        RECT -1.140 92.040 -1.000 92.440 ;
        RECT 3.820 92.040 3.960 92.440 ;
        RECT 5.690 92.040 7.050 92.350 ;
        RECT 8.780 92.040 8.920 92.440 ;
        RECT 13.740 92.040 13.880 92.440 ;
        RECT 15.610 92.040 16.970 92.350 ;
        RECT 18.700 92.040 18.840 92.440 ;
        RECT 23.660 92.040 23.800 92.440 ;
        RECT 37.260 92.370 37.720 96.680 ;
        RECT 32.950 92.360 37.720 92.370 ;
        RECT 25.530 92.040 37.720 92.360 ;
        RECT -291.010 91.910 37.720 92.040 ;
        RECT -291.010 91.900 34.270 91.910 ;
        RECT -288.820 91.500 -288.680 91.900 ;
        RECT -286.950 91.590 -285.590 91.900 ;
        RECT -283.860 91.500 -283.720 91.900 ;
        RECT -278.900 91.500 -278.760 91.900 ;
        RECT -277.030 91.590 -275.670 91.900 ;
        RECT -273.940 91.500 -273.800 91.900 ;
        RECT -268.980 91.500 -268.840 91.900 ;
        RECT -267.110 91.590 -265.750 91.900 ;
        RECT -264.020 91.500 -263.880 91.900 ;
        RECT -259.060 91.500 -258.920 91.900 ;
        RECT -257.190 91.590 -255.830 91.900 ;
        RECT -254.100 91.500 -253.960 91.900 ;
        RECT -249.140 91.500 -249.000 91.900 ;
        RECT -247.270 91.590 -245.910 91.900 ;
        RECT -244.180 91.500 -244.040 91.900 ;
        RECT -239.220 91.500 -239.080 91.900 ;
        RECT -237.350 91.590 -235.990 91.900 ;
        RECT -234.260 91.500 -234.120 91.900 ;
        RECT -229.300 91.500 -229.160 91.900 ;
        RECT -227.430 91.590 -226.070 91.900 ;
        RECT -224.340 91.500 -224.200 91.900 ;
        RECT -219.380 91.500 -219.240 91.900 ;
        RECT -217.510 91.590 -216.150 91.900 ;
        RECT -214.420 91.500 -214.280 91.900 ;
        RECT -209.460 91.500 -209.320 91.900 ;
        RECT -207.590 91.590 -206.230 91.900 ;
        RECT -204.500 91.500 -204.360 91.900 ;
        RECT -199.540 91.500 -199.400 91.900 ;
        RECT -197.670 91.590 -196.310 91.900 ;
        RECT -194.580 91.500 -194.440 91.900 ;
        RECT -189.620 91.500 -189.480 91.900 ;
        RECT -187.750 91.590 -186.390 91.900 ;
        RECT -184.660 91.500 -184.520 91.900 ;
        RECT -179.700 91.500 -179.560 91.900 ;
        RECT -177.830 91.590 -176.470 91.900 ;
        RECT -174.740 91.500 -174.600 91.900 ;
        RECT -169.780 91.500 -169.640 91.900 ;
        RECT -167.910 91.590 -166.550 91.900 ;
        RECT -164.820 91.500 -164.680 91.900 ;
        RECT -159.860 91.500 -159.720 91.900 ;
        RECT -157.990 91.590 -156.630 91.900 ;
        RECT -154.900 91.500 -154.760 91.900 ;
        RECT -149.940 91.500 -149.800 91.900 ;
        RECT -148.070 91.590 -146.710 91.900 ;
        RECT -144.980 91.500 -144.840 91.900 ;
        RECT -140.020 91.500 -139.880 91.900 ;
        RECT -138.150 91.590 -136.790 91.900 ;
        RECT -135.060 91.500 -134.920 91.900 ;
        RECT -130.100 91.500 -129.960 91.900 ;
        RECT -128.230 91.590 -126.870 91.900 ;
        RECT -125.140 91.500 -125.000 91.900 ;
        RECT -120.180 91.500 -120.040 91.900 ;
        RECT -118.310 91.590 -116.950 91.900 ;
        RECT -115.220 91.500 -115.080 91.900 ;
        RECT -110.260 91.500 -110.120 91.900 ;
        RECT -108.390 91.590 -107.030 91.900 ;
        RECT -105.300 91.500 -105.160 91.900 ;
        RECT -100.340 91.500 -100.200 91.900 ;
        RECT -98.470 91.590 -97.110 91.900 ;
        RECT -95.380 91.500 -95.240 91.900 ;
        RECT -90.420 91.500 -90.280 91.900 ;
        RECT -88.550 91.590 -87.190 91.900 ;
        RECT -85.460 91.500 -85.320 91.900 ;
        RECT -80.500 91.500 -80.360 91.900 ;
        RECT -78.630 91.590 -77.270 91.900 ;
        RECT -75.540 91.500 -75.400 91.900 ;
        RECT -70.580 91.500 -70.440 91.900 ;
        RECT -68.710 91.590 -67.350 91.900 ;
        RECT -65.620 91.500 -65.480 91.900 ;
        RECT -60.660 91.500 -60.520 91.900 ;
        RECT -58.790 91.590 -57.430 91.900 ;
        RECT -55.700 91.500 -55.560 91.900 ;
        RECT -50.740 91.500 -50.600 91.900 ;
        RECT -48.870 91.590 -47.510 91.900 ;
        RECT -45.780 91.500 -45.640 91.900 ;
        RECT -40.820 91.500 -40.680 91.900 ;
        RECT -38.950 91.590 -37.590 91.900 ;
        RECT -35.860 91.500 -35.720 91.900 ;
        RECT -30.900 91.500 -30.760 91.900 ;
        RECT -29.030 91.590 -27.670 91.900 ;
        RECT -25.940 91.500 -25.800 91.900 ;
        RECT -20.980 91.500 -20.840 91.900 ;
        RECT -19.110 91.590 -17.750 91.900 ;
        RECT -16.020 91.500 -15.880 91.900 ;
        RECT -11.060 91.500 -10.920 91.900 ;
        RECT -9.190 91.590 -7.830 91.900 ;
        RECT -6.100 91.500 -5.960 91.900 ;
        RECT -1.140 91.500 -1.000 91.900 ;
        RECT 0.730 91.590 2.090 91.900 ;
        RECT 3.820 91.500 3.960 91.900 ;
        RECT 8.780 91.500 8.920 91.900 ;
        RECT 10.650 91.590 12.010 91.900 ;
        RECT 13.740 91.500 13.880 91.900 ;
        RECT 18.700 91.500 18.840 91.900 ;
        RECT 20.570 91.590 21.930 91.900 ;
        RECT 23.660 91.500 23.800 91.900 ;
    END
  END i_srclk
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -288.220 95.135 -284.260 95.140 ;
        RECT -278.300 95.135 -274.340 95.140 ;
        RECT -268.380 95.135 -264.420 95.140 ;
        RECT -258.460 95.135 -254.500 95.140 ;
        RECT -248.540 95.135 -244.580 95.140 ;
        RECT -238.620 95.135 -234.660 95.140 ;
        RECT -228.700 95.135 -224.740 95.140 ;
        RECT -218.780 95.135 -214.820 95.140 ;
        RECT -208.860 95.135 -204.900 95.140 ;
        RECT -198.940 95.135 -194.980 95.140 ;
        RECT -189.020 95.135 -185.060 95.140 ;
        RECT -179.100 95.135 -175.140 95.140 ;
        RECT -169.180 95.135 -165.220 95.140 ;
        RECT -159.260 95.135 -155.300 95.140 ;
        RECT -149.340 95.135 -145.380 95.140 ;
        RECT -139.420 95.135 -135.460 95.140 ;
        RECT -129.500 95.135 -125.540 95.140 ;
        RECT -119.580 95.135 -115.620 95.140 ;
        RECT -109.660 95.135 -105.700 95.140 ;
        RECT -99.740 95.135 -95.780 95.140 ;
        RECT -89.820 95.135 -85.860 95.140 ;
        RECT -79.900 95.135 -75.940 95.140 ;
        RECT -69.980 95.135 -66.020 95.140 ;
        RECT -60.060 95.135 -56.100 95.140 ;
        RECT -50.140 95.135 -46.180 95.140 ;
        RECT -40.220 95.135 -36.260 95.140 ;
        RECT -30.300 95.135 -26.340 95.140 ;
        RECT -20.380 95.135 -16.420 95.140 ;
        RECT -10.460 95.135 -6.500 95.140 ;
        RECT -0.540 95.135 3.420 95.140 ;
        RECT 9.380 95.135 13.340 95.140 ;
        RECT 19.300 95.135 23.260 95.140 ;
        RECT -288.925 93.765 -283.615 95.135 ;
        RECT -279.005 93.765 -273.695 95.135 ;
        RECT -269.085 93.765 -263.775 95.135 ;
        RECT -259.165 93.765 -253.855 95.135 ;
        RECT -249.245 93.765 -243.935 95.135 ;
        RECT -239.325 93.765 -234.015 95.135 ;
        RECT -229.405 93.765 -224.095 95.135 ;
        RECT -219.485 93.765 -214.175 95.135 ;
        RECT -209.565 93.765 -204.255 95.135 ;
        RECT -199.645 93.765 -194.335 95.135 ;
        RECT -189.725 93.765 -184.415 95.135 ;
        RECT -179.805 93.765 -174.495 95.135 ;
        RECT -169.885 93.765 -164.575 95.135 ;
        RECT -159.965 93.765 -154.655 95.135 ;
        RECT -150.045 93.765 -144.735 95.135 ;
        RECT -140.125 93.765 -134.815 95.135 ;
        RECT -130.205 93.765 -124.895 95.135 ;
        RECT -120.285 93.765 -114.975 95.135 ;
        RECT -110.365 93.765 -105.055 95.135 ;
        RECT -100.445 93.765 -95.135 95.135 ;
        RECT -90.525 93.765 -85.215 95.135 ;
        RECT -80.605 93.765 -75.295 95.135 ;
        RECT -70.685 93.765 -65.375 95.135 ;
        RECT -60.765 93.765 -55.455 95.135 ;
        RECT -50.845 93.765 -45.535 95.135 ;
        RECT -40.925 93.765 -35.615 95.135 ;
        RECT -31.005 93.765 -25.695 95.135 ;
        RECT -21.085 93.765 -15.775 95.135 ;
        RECT -11.165 93.765 -5.855 95.135 ;
        RECT -1.245 93.765 4.065 95.135 ;
        RECT 8.675 93.765 13.985 95.135 ;
        RECT 18.595 93.765 23.905 95.135 ;
        RECT -288.220 93.760 -284.260 93.765 ;
        RECT -278.300 93.760 -274.340 93.765 ;
        RECT -268.380 93.760 -264.420 93.765 ;
        RECT -258.460 93.760 -254.500 93.765 ;
        RECT -248.540 93.760 -244.580 93.765 ;
        RECT -238.620 93.760 -234.660 93.765 ;
        RECT -228.700 93.760 -224.740 93.765 ;
        RECT -218.780 93.760 -214.820 93.765 ;
        RECT -208.860 93.760 -204.900 93.765 ;
        RECT -198.940 93.760 -194.980 93.765 ;
        RECT -189.020 93.760 -185.060 93.765 ;
        RECT -179.100 93.760 -175.140 93.765 ;
        RECT -169.180 93.760 -165.220 93.765 ;
        RECT -159.260 93.760 -155.300 93.765 ;
        RECT -149.340 93.760 -145.380 93.765 ;
        RECT -139.420 93.760 -135.460 93.765 ;
        RECT -129.500 93.760 -125.540 93.765 ;
        RECT -119.580 93.760 -115.620 93.765 ;
        RECT -109.660 93.760 -105.700 93.765 ;
        RECT -99.740 93.760 -95.780 93.765 ;
        RECT -89.820 93.760 -85.860 93.765 ;
        RECT -79.900 93.760 -75.940 93.765 ;
        RECT -69.980 93.760 -66.020 93.765 ;
        RECT -60.060 93.760 -56.100 93.765 ;
        RECT -50.140 93.760 -46.180 93.765 ;
        RECT -40.220 93.760 -36.260 93.765 ;
        RECT -30.300 93.760 -26.340 93.765 ;
        RECT -20.380 93.760 -16.420 93.765 ;
        RECT -10.460 93.760 -6.500 93.765 ;
        RECT -0.540 93.760 3.420 93.765 ;
        RECT 9.380 93.760 13.340 93.765 ;
        RECT 19.300 93.760 23.260 93.765 ;
        RECT -281.850 93.225 -281.680 93.415 ;
        RECT -280.940 93.225 -280.770 93.415 ;
        RECT -271.930 93.225 -271.760 93.415 ;
        RECT -271.020 93.225 -270.850 93.415 ;
        RECT -262.010 93.225 -261.840 93.415 ;
        RECT -261.100 93.225 -260.930 93.415 ;
        RECT -252.090 93.225 -251.920 93.415 ;
        RECT -251.180 93.225 -251.010 93.415 ;
        RECT -242.170 93.225 -242.000 93.415 ;
        RECT -241.260 93.225 -241.090 93.415 ;
        RECT -232.250 93.225 -232.080 93.415 ;
        RECT -231.340 93.225 -231.170 93.415 ;
        RECT -222.330 93.225 -222.160 93.415 ;
        RECT -221.420 93.225 -221.250 93.415 ;
        RECT -212.410 93.225 -212.240 93.415 ;
        RECT -211.500 93.225 -211.330 93.415 ;
        RECT -202.490 93.225 -202.320 93.415 ;
        RECT -201.580 93.225 -201.410 93.415 ;
        RECT -192.570 93.225 -192.400 93.415 ;
        RECT -191.660 93.225 -191.490 93.415 ;
        RECT -182.650 93.225 -182.480 93.415 ;
        RECT -181.740 93.225 -181.570 93.415 ;
        RECT -172.730 93.225 -172.560 93.415 ;
        RECT -171.820 93.225 -171.650 93.415 ;
        RECT -162.810 93.225 -162.640 93.415 ;
        RECT -161.900 93.225 -161.730 93.415 ;
        RECT -152.890 93.225 -152.720 93.415 ;
        RECT -151.980 93.225 -151.810 93.415 ;
        RECT -142.970 93.225 -142.800 93.415 ;
        RECT -142.060 93.225 -141.890 93.415 ;
        RECT -133.050 93.225 -132.880 93.415 ;
        RECT -132.140 93.225 -131.970 93.415 ;
        RECT -123.130 93.225 -122.960 93.415 ;
        RECT -122.220 93.225 -122.050 93.415 ;
        RECT -113.210 93.225 -113.040 93.415 ;
        RECT -112.300 93.225 -112.130 93.415 ;
        RECT -103.290 93.225 -103.120 93.415 ;
        RECT -102.380 93.225 -102.210 93.415 ;
        RECT -93.370 93.225 -93.200 93.415 ;
        RECT -92.460 93.225 -92.290 93.415 ;
        RECT -83.450 93.225 -83.280 93.415 ;
        RECT -82.540 93.225 -82.370 93.415 ;
        RECT -73.530 93.225 -73.360 93.415 ;
        RECT -72.620 93.225 -72.450 93.415 ;
        RECT -63.610 93.225 -63.440 93.415 ;
        RECT -62.700 93.225 -62.530 93.415 ;
        RECT -53.690 93.225 -53.520 93.415 ;
        RECT -52.780 93.225 -52.610 93.415 ;
        RECT -43.770 93.225 -43.600 93.415 ;
        RECT -42.860 93.225 -42.690 93.415 ;
        RECT -33.850 93.225 -33.680 93.415 ;
        RECT -32.940 93.225 -32.770 93.415 ;
        RECT -23.930 93.225 -23.760 93.415 ;
        RECT -23.020 93.225 -22.850 93.415 ;
        RECT -14.010 93.225 -13.840 93.415 ;
        RECT -13.100 93.225 -12.930 93.415 ;
        RECT -4.090 93.225 -3.920 93.415 ;
        RECT -3.180 93.225 -3.010 93.415 ;
        RECT 5.830 93.225 6.000 93.415 ;
        RECT 6.740 93.225 6.910 93.415 ;
        RECT 15.750 93.225 15.920 93.415 ;
        RECT 16.660 93.225 16.830 93.415 ;
        RECT -282.915 93.220 -281.565 93.225 ;
        RECT -281.055 93.220 -279.705 93.225 ;
        RECT -282.915 92.320 -279.705 93.220 ;
        RECT -282.915 92.315 -281.565 92.320 ;
        RECT -281.055 92.315 -279.705 92.320 ;
        RECT -272.995 93.220 -271.645 93.225 ;
        RECT -271.135 93.220 -269.785 93.225 ;
        RECT -272.995 92.320 -269.785 93.220 ;
        RECT -272.995 92.315 -271.645 92.320 ;
        RECT -271.135 92.315 -269.785 92.320 ;
        RECT -263.075 93.220 -261.725 93.225 ;
        RECT -261.215 93.220 -259.865 93.225 ;
        RECT -263.075 92.320 -259.865 93.220 ;
        RECT -263.075 92.315 -261.725 92.320 ;
        RECT -261.215 92.315 -259.865 92.320 ;
        RECT -253.155 93.220 -251.805 93.225 ;
        RECT -251.295 93.220 -249.945 93.225 ;
        RECT -253.155 92.320 -249.945 93.220 ;
        RECT -253.155 92.315 -251.805 92.320 ;
        RECT -251.295 92.315 -249.945 92.320 ;
        RECT -243.235 93.220 -241.885 93.225 ;
        RECT -241.375 93.220 -240.025 93.225 ;
        RECT -243.235 92.320 -240.025 93.220 ;
        RECT -243.235 92.315 -241.885 92.320 ;
        RECT -241.375 92.315 -240.025 92.320 ;
        RECT -233.315 93.220 -231.965 93.225 ;
        RECT -231.455 93.220 -230.105 93.225 ;
        RECT -233.315 92.320 -230.105 93.220 ;
        RECT -233.315 92.315 -231.965 92.320 ;
        RECT -231.455 92.315 -230.105 92.320 ;
        RECT -223.395 93.220 -222.045 93.225 ;
        RECT -221.535 93.220 -220.185 93.225 ;
        RECT -223.395 92.320 -220.185 93.220 ;
        RECT -223.395 92.315 -222.045 92.320 ;
        RECT -221.535 92.315 -220.185 92.320 ;
        RECT -213.475 93.220 -212.125 93.225 ;
        RECT -211.615 93.220 -210.265 93.225 ;
        RECT -213.475 92.320 -210.265 93.220 ;
        RECT -213.475 92.315 -212.125 92.320 ;
        RECT -211.615 92.315 -210.265 92.320 ;
        RECT -203.555 93.220 -202.205 93.225 ;
        RECT -201.695 93.220 -200.345 93.225 ;
        RECT -203.555 92.320 -200.345 93.220 ;
        RECT -203.555 92.315 -202.205 92.320 ;
        RECT -201.695 92.315 -200.345 92.320 ;
        RECT -193.635 93.220 -192.285 93.225 ;
        RECT -191.775 93.220 -190.425 93.225 ;
        RECT -193.635 92.320 -190.425 93.220 ;
        RECT -193.635 92.315 -192.285 92.320 ;
        RECT -191.775 92.315 -190.425 92.320 ;
        RECT -183.715 93.220 -182.365 93.225 ;
        RECT -181.855 93.220 -180.505 93.225 ;
        RECT -183.715 92.320 -180.505 93.220 ;
        RECT -183.715 92.315 -182.365 92.320 ;
        RECT -181.855 92.315 -180.505 92.320 ;
        RECT -173.795 93.220 -172.445 93.225 ;
        RECT -171.935 93.220 -170.585 93.225 ;
        RECT -173.795 92.320 -170.585 93.220 ;
        RECT -173.795 92.315 -172.445 92.320 ;
        RECT -171.935 92.315 -170.585 92.320 ;
        RECT -163.875 93.220 -162.525 93.225 ;
        RECT -162.015 93.220 -160.665 93.225 ;
        RECT -163.875 92.320 -160.665 93.220 ;
        RECT -163.875 92.315 -162.525 92.320 ;
        RECT -162.015 92.315 -160.665 92.320 ;
        RECT -153.955 93.220 -152.605 93.225 ;
        RECT -152.095 93.220 -150.745 93.225 ;
        RECT -153.955 92.320 -150.745 93.220 ;
        RECT -153.955 92.315 -152.605 92.320 ;
        RECT -152.095 92.315 -150.745 92.320 ;
        RECT -144.035 93.220 -142.685 93.225 ;
        RECT -142.175 93.220 -140.825 93.225 ;
        RECT -144.035 92.320 -140.825 93.220 ;
        RECT -144.035 92.315 -142.685 92.320 ;
        RECT -142.175 92.315 -140.825 92.320 ;
        RECT -134.115 93.220 -132.765 93.225 ;
        RECT -132.255 93.220 -130.905 93.225 ;
        RECT -134.115 92.320 -130.905 93.220 ;
        RECT -134.115 92.315 -132.765 92.320 ;
        RECT -132.255 92.315 -130.905 92.320 ;
        RECT -124.195 93.220 -122.845 93.225 ;
        RECT -122.335 93.220 -120.985 93.225 ;
        RECT -124.195 92.320 -120.985 93.220 ;
        RECT -124.195 92.315 -122.845 92.320 ;
        RECT -122.335 92.315 -120.985 92.320 ;
        RECT -114.275 93.220 -112.925 93.225 ;
        RECT -112.415 93.220 -111.065 93.225 ;
        RECT -114.275 92.320 -111.065 93.220 ;
        RECT -114.275 92.315 -112.925 92.320 ;
        RECT -112.415 92.315 -111.065 92.320 ;
        RECT -104.355 93.220 -103.005 93.225 ;
        RECT -102.495 93.220 -101.145 93.225 ;
        RECT -104.355 92.320 -101.145 93.220 ;
        RECT -104.355 92.315 -103.005 92.320 ;
        RECT -102.495 92.315 -101.145 92.320 ;
        RECT -94.435 93.220 -93.085 93.225 ;
        RECT -92.575 93.220 -91.225 93.225 ;
        RECT -94.435 92.320 -91.225 93.220 ;
        RECT -94.435 92.315 -93.085 92.320 ;
        RECT -92.575 92.315 -91.225 92.320 ;
        RECT -84.515 93.220 -83.165 93.225 ;
        RECT -82.655 93.220 -81.305 93.225 ;
        RECT -84.515 92.320 -81.305 93.220 ;
        RECT -84.515 92.315 -83.165 92.320 ;
        RECT -82.655 92.315 -81.305 92.320 ;
        RECT -74.595 93.220 -73.245 93.225 ;
        RECT -72.735 93.220 -71.385 93.225 ;
        RECT -74.595 92.320 -71.385 93.220 ;
        RECT -74.595 92.315 -73.245 92.320 ;
        RECT -72.735 92.315 -71.385 92.320 ;
        RECT -64.675 93.220 -63.325 93.225 ;
        RECT -62.815 93.220 -61.465 93.225 ;
        RECT -64.675 92.320 -61.465 93.220 ;
        RECT -64.675 92.315 -63.325 92.320 ;
        RECT -62.815 92.315 -61.465 92.320 ;
        RECT -54.755 93.220 -53.405 93.225 ;
        RECT -52.895 93.220 -51.545 93.225 ;
        RECT -54.755 92.320 -51.545 93.220 ;
        RECT -54.755 92.315 -53.405 92.320 ;
        RECT -52.895 92.315 -51.545 92.320 ;
        RECT -44.835 93.220 -43.485 93.225 ;
        RECT -42.975 93.220 -41.625 93.225 ;
        RECT -44.835 92.320 -41.625 93.220 ;
        RECT -44.835 92.315 -43.485 92.320 ;
        RECT -42.975 92.315 -41.625 92.320 ;
        RECT -34.915 93.220 -33.565 93.225 ;
        RECT -33.055 93.220 -31.705 93.225 ;
        RECT -34.915 92.320 -31.705 93.220 ;
        RECT -34.915 92.315 -33.565 92.320 ;
        RECT -33.055 92.315 -31.705 92.320 ;
        RECT -24.995 93.220 -23.645 93.225 ;
        RECT -23.135 93.220 -21.785 93.225 ;
        RECT -24.995 92.320 -21.785 93.220 ;
        RECT -24.995 92.315 -23.645 92.320 ;
        RECT -23.135 92.315 -21.785 92.320 ;
        RECT -15.075 93.220 -13.725 93.225 ;
        RECT -13.215 93.220 -11.865 93.225 ;
        RECT -15.075 92.320 -11.865 93.220 ;
        RECT -15.075 92.315 -13.725 92.320 ;
        RECT -13.215 92.315 -11.865 92.320 ;
        RECT -5.155 93.220 -3.805 93.225 ;
        RECT -3.295 93.220 -1.945 93.225 ;
        RECT -5.155 92.320 -1.945 93.220 ;
        RECT -5.155 92.315 -3.805 92.320 ;
        RECT -3.295 92.315 -1.945 92.320 ;
        RECT 4.765 93.220 6.115 93.225 ;
        RECT 6.625 93.220 7.975 93.225 ;
        RECT 4.765 92.320 7.975 93.220 ;
        RECT 4.765 92.315 6.115 92.320 ;
        RECT 6.625 92.315 7.975 92.320 ;
        RECT 14.685 93.220 16.035 93.225 ;
        RECT 16.545 93.220 17.895 93.225 ;
        RECT 14.685 92.320 17.895 93.220 ;
        RECT 14.685 92.315 16.035 92.320 ;
        RECT 16.545 92.315 17.895 92.320 ;
        RECT -287.875 91.620 -286.525 91.625 ;
        RECT -286.015 91.620 -284.665 91.625 ;
        RECT -287.875 90.720 -284.665 91.620 ;
        RECT -287.875 90.715 -286.525 90.720 ;
        RECT -286.015 90.715 -284.665 90.720 ;
        RECT -277.955 91.620 -276.605 91.625 ;
        RECT -276.095 91.620 -274.745 91.625 ;
        RECT -277.955 90.720 -274.745 91.620 ;
        RECT -277.955 90.715 -276.605 90.720 ;
        RECT -276.095 90.715 -274.745 90.720 ;
        RECT -268.035 91.620 -266.685 91.625 ;
        RECT -266.175 91.620 -264.825 91.625 ;
        RECT -268.035 90.720 -264.825 91.620 ;
        RECT -268.035 90.715 -266.685 90.720 ;
        RECT -266.175 90.715 -264.825 90.720 ;
        RECT -258.115 91.620 -256.765 91.625 ;
        RECT -256.255 91.620 -254.905 91.625 ;
        RECT -258.115 90.720 -254.905 91.620 ;
        RECT -258.115 90.715 -256.765 90.720 ;
        RECT -256.255 90.715 -254.905 90.720 ;
        RECT -248.195 91.620 -246.845 91.625 ;
        RECT -246.335 91.620 -244.985 91.625 ;
        RECT -248.195 90.720 -244.985 91.620 ;
        RECT -248.195 90.715 -246.845 90.720 ;
        RECT -246.335 90.715 -244.985 90.720 ;
        RECT -238.275 91.620 -236.925 91.625 ;
        RECT -236.415 91.620 -235.065 91.625 ;
        RECT -238.275 90.720 -235.065 91.620 ;
        RECT -238.275 90.715 -236.925 90.720 ;
        RECT -236.415 90.715 -235.065 90.720 ;
        RECT -228.355 91.620 -227.005 91.625 ;
        RECT -226.495 91.620 -225.145 91.625 ;
        RECT -228.355 90.720 -225.145 91.620 ;
        RECT -228.355 90.715 -227.005 90.720 ;
        RECT -226.495 90.715 -225.145 90.720 ;
        RECT -218.435 91.620 -217.085 91.625 ;
        RECT -216.575 91.620 -215.225 91.625 ;
        RECT -218.435 90.720 -215.225 91.620 ;
        RECT -218.435 90.715 -217.085 90.720 ;
        RECT -216.575 90.715 -215.225 90.720 ;
        RECT -208.515 91.620 -207.165 91.625 ;
        RECT -206.655 91.620 -205.305 91.625 ;
        RECT -208.515 90.720 -205.305 91.620 ;
        RECT -208.515 90.715 -207.165 90.720 ;
        RECT -206.655 90.715 -205.305 90.720 ;
        RECT -198.595 91.620 -197.245 91.625 ;
        RECT -196.735 91.620 -195.385 91.625 ;
        RECT -198.595 90.720 -195.385 91.620 ;
        RECT -198.595 90.715 -197.245 90.720 ;
        RECT -196.735 90.715 -195.385 90.720 ;
        RECT -188.675 91.620 -187.325 91.625 ;
        RECT -186.815 91.620 -185.465 91.625 ;
        RECT -188.675 90.720 -185.465 91.620 ;
        RECT -188.675 90.715 -187.325 90.720 ;
        RECT -186.815 90.715 -185.465 90.720 ;
        RECT -178.755 91.620 -177.405 91.625 ;
        RECT -176.895 91.620 -175.545 91.625 ;
        RECT -178.755 90.720 -175.545 91.620 ;
        RECT -178.755 90.715 -177.405 90.720 ;
        RECT -176.895 90.715 -175.545 90.720 ;
        RECT -168.835 91.620 -167.485 91.625 ;
        RECT -166.975 91.620 -165.625 91.625 ;
        RECT -168.835 90.720 -165.625 91.620 ;
        RECT -168.835 90.715 -167.485 90.720 ;
        RECT -166.975 90.715 -165.625 90.720 ;
        RECT -158.915 91.620 -157.565 91.625 ;
        RECT -157.055 91.620 -155.705 91.625 ;
        RECT -158.915 90.720 -155.705 91.620 ;
        RECT -158.915 90.715 -157.565 90.720 ;
        RECT -157.055 90.715 -155.705 90.720 ;
        RECT -148.995 91.620 -147.645 91.625 ;
        RECT -147.135 91.620 -145.785 91.625 ;
        RECT -148.995 90.720 -145.785 91.620 ;
        RECT -148.995 90.715 -147.645 90.720 ;
        RECT -147.135 90.715 -145.785 90.720 ;
        RECT -139.075 91.620 -137.725 91.625 ;
        RECT -137.215 91.620 -135.865 91.625 ;
        RECT -139.075 90.720 -135.865 91.620 ;
        RECT -139.075 90.715 -137.725 90.720 ;
        RECT -137.215 90.715 -135.865 90.720 ;
        RECT -129.155 91.620 -127.805 91.625 ;
        RECT -127.295 91.620 -125.945 91.625 ;
        RECT -129.155 90.720 -125.945 91.620 ;
        RECT -129.155 90.715 -127.805 90.720 ;
        RECT -127.295 90.715 -125.945 90.720 ;
        RECT -119.235 91.620 -117.885 91.625 ;
        RECT -117.375 91.620 -116.025 91.625 ;
        RECT -119.235 90.720 -116.025 91.620 ;
        RECT -119.235 90.715 -117.885 90.720 ;
        RECT -117.375 90.715 -116.025 90.720 ;
        RECT -109.315 91.620 -107.965 91.625 ;
        RECT -107.455 91.620 -106.105 91.625 ;
        RECT -109.315 90.720 -106.105 91.620 ;
        RECT -109.315 90.715 -107.965 90.720 ;
        RECT -107.455 90.715 -106.105 90.720 ;
        RECT -99.395 91.620 -98.045 91.625 ;
        RECT -97.535 91.620 -96.185 91.625 ;
        RECT -99.395 90.720 -96.185 91.620 ;
        RECT -99.395 90.715 -98.045 90.720 ;
        RECT -97.535 90.715 -96.185 90.720 ;
        RECT -89.475 91.620 -88.125 91.625 ;
        RECT -87.615 91.620 -86.265 91.625 ;
        RECT -89.475 90.720 -86.265 91.620 ;
        RECT -89.475 90.715 -88.125 90.720 ;
        RECT -87.615 90.715 -86.265 90.720 ;
        RECT -79.555 91.620 -78.205 91.625 ;
        RECT -77.695 91.620 -76.345 91.625 ;
        RECT -79.555 90.720 -76.345 91.620 ;
        RECT -79.555 90.715 -78.205 90.720 ;
        RECT -77.695 90.715 -76.345 90.720 ;
        RECT -69.635 91.620 -68.285 91.625 ;
        RECT -67.775 91.620 -66.425 91.625 ;
        RECT -69.635 90.720 -66.425 91.620 ;
        RECT -69.635 90.715 -68.285 90.720 ;
        RECT -67.775 90.715 -66.425 90.720 ;
        RECT -59.715 91.620 -58.365 91.625 ;
        RECT -57.855 91.620 -56.505 91.625 ;
        RECT -59.715 90.720 -56.505 91.620 ;
        RECT -59.715 90.715 -58.365 90.720 ;
        RECT -57.855 90.715 -56.505 90.720 ;
        RECT -49.795 91.620 -48.445 91.625 ;
        RECT -47.935 91.620 -46.585 91.625 ;
        RECT -49.795 90.720 -46.585 91.620 ;
        RECT -49.795 90.715 -48.445 90.720 ;
        RECT -47.935 90.715 -46.585 90.720 ;
        RECT -39.875 91.620 -38.525 91.625 ;
        RECT -38.015 91.620 -36.665 91.625 ;
        RECT -39.875 90.720 -36.665 91.620 ;
        RECT -39.875 90.715 -38.525 90.720 ;
        RECT -38.015 90.715 -36.665 90.720 ;
        RECT -29.955 91.620 -28.605 91.625 ;
        RECT -28.095 91.620 -26.745 91.625 ;
        RECT -29.955 90.720 -26.745 91.620 ;
        RECT -29.955 90.715 -28.605 90.720 ;
        RECT -28.095 90.715 -26.745 90.720 ;
        RECT -20.035 91.620 -18.685 91.625 ;
        RECT -18.175 91.620 -16.825 91.625 ;
        RECT -20.035 90.720 -16.825 91.620 ;
        RECT -20.035 90.715 -18.685 90.720 ;
        RECT -18.175 90.715 -16.825 90.720 ;
        RECT -10.115 91.620 -8.765 91.625 ;
        RECT -8.255 91.620 -6.905 91.625 ;
        RECT -10.115 90.720 -6.905 91.620 ;
        RECT -10.115 90.715 -8.765 90.720 ;
        RECT -8.255 90.715 -6.905 90.720 ;
        RECT -0.195 91.620 1.155 91.625 ;
        RECT 1.665 91.620 3.015 91.625 ;
        RECT -0.195 90.720 3.015 91.620 ;
        RECT -0.195 90.715 1.155 90.720 ;
        RECT 1.665 90.715 3.015 90.720 ;
        RECT 9.725 91.620 11.075 91.625 ;
        RECT 11.585 91.620 12.935 91.625 ;
        RECT 9.725 90.720 12.935 91.620 ;
        RECT 9.725 90.715 11.075 90.720 ;
        RECT 11.585 90.715 12.935 90.720 ;
        RECT 19.645 91.620 20.995 91.625 ;
        RECT 21.505 91.620 22.855 91.625 ;
        RECT 19.645 90.720 22.855 91.620 ;
        RECT 19.645 90.715 20.995 90.720 ;
        RECT 21.505 90.715 22.855 90.720 ;
        RECT -286.810 90.525 -286.640 90.715 ;
        RECT -285.900 90.525 -285.730 90.715 ;
        RECT -276.890 90.525 -276.720 90.715 ;
        RECT -275.980 90.525 -275.810 90.715 ;
        RECT -266.970 90.525 -266.800 90.715 ;
        RECT -266.060 90.525 -265.890 90.715 ;
        RECT -257.050 90.525 -256.880 90.715 ;
        RECT -256.140 90.525 -255.970 90.715 ;
        RECT -247.130 90.525 -246.960 90.715 ;
        RECT -246.220 90.525 -246.050 90.715 ;
        RECT -237.210 90.525 -237.040 90.715 ;
        RECT -236.300 90.525 -236.130 90.715 ;
        RECT -227.290 90.525 -227.120 90.715 ;
        RECT -226.380 90.525 -226.210 90.715 ;
        RECT -217.370 90.525 -217.200 90.715 ;
        RECT -216.460 90.525 -216.290 90.715 ;
        RECT -207.450 90.525 -207.280 90.715 ;
        RECT -206.540 90.525 -206.370 90.715 ;
        RECT -197.530 90.525 -197.360 90.715 ;
        RECT -196.620 90.525 -196.450 90.715 ;
        RECT -187.610 90.525 -187.440 90.715 ;
        RECT -186.700 90.525 -186.530 90.715 ;
        RECT -177.690 90.525 -177.520 90.715 ;
        RECT -176.780 90.525 -176.610 90.715 ;
        RECT -167.770 90.525 -167.600 90.715 ;
        RECT -166.860 90.525 -166.690 90.715 ;
        RECT -157.850 90.525 -157.680 90.715 ;
        RECT -156.940 90.525 -156.770 90.715 ;
        RECT -147.930 90.525 -147.760 90.715 ;
        RECT -147.020 90.525 -146.850 90.715 ;
        RECT -138.010 90.525 -137.840 90.715 ;
        RECT -137.100 90.525 -136.930 90.715 ;
        RECT -128.090 90.525 -127.920 90.715 ;
        RECT -127.180 90.525 -127.010 90.715 ;
        RECT -118.170 90.525 -118.000 90.715 ;
        RECT -117.260 90.525 -117.090 90.715 ;
        RECT -108.250 90.525 -108.080 90.715 ;
        RECT -107.340 90.525 -107.170 90.715 ;
        RECT -98.330 90.525 -98.160 90.715 ;
        RECT -97.420 90.525 -97.250 90.715 ;
        RECT -88.410 90.525 -88.240 90.715 ;
        RECT -87.500 90.525 -87.330 90.715 ;
        RECT -78.490 90.525 -78.320 90.715 ;
        RECT -77.580 90.525 -77.410 90.715 ;
        RECT -68.570 90.525 -68.400 90.715 ;
        RECT -67.660 90.525 -67.490 90.715 ;
        RECT -58.650 90.525 -58.480 90.715 ;
        RECT -57.740 90.525 -57.570 90.715 ;
        RECT -48.730 90.525 -48.560 90.715 ;
        RECT -47.820 90.525 -47.650 90.715 ;
        RECT -38.810 90.525 -38.640 90.715 ;
        RECT -37.900 90.525 -37.730 90.715 ;
        RECT -28.890 90.525 -28.720 90.715 ;
        RECT -27.980 90.525 -27.810 90.715 ;
        RECT -18.970 90.525 -18.800 90.715 ;
        RECT -18.060 90.525 -17.890 90.715 ;
        RECT -9.050 90.525 -8.880 90.715 ;
        RECT -8.140 90.525 -7.970 90.715 ;
        RECT 0.870 90.525 1.040 90.715 ;
        RECT 1.780 90.525 1.950 90.715 ;
        RECT 10.790 90.525 10.960 90.715 ;
        RECT 11.700 90.525 11.870 90.715 ;
        RECT 20.710 90.525 20.880 90.715 ;
        RECT 21.620 90.525 21.790 90.715 ;
        RECT -281.525 90.180 -281.095 90.195 ;
        RECT -271.605 90.180 -271.175 90.195 ;
        RECT -261.685 90.180 -261.255 90.195 ;
        RECT -251.765 90.180 -251.335 90.195 ;
        RECT -241.845 90.180 -241.415 90.195 ;
        RECT -231.925 90.180 -231.495 90.195 ;
        RECT -222.005 90.180 -221.575 90.195 ;
        RECT -212.085 90.180 -211.655 90.195 ;
        RECT -202.165 90.180 -201.735 90.195 ;
        RECT -192.245 90.180 -191.815 90.195 ;
        RECT -182.325 90.180 -181.895 90.195 ;
        RECT -172.405 90.180 -171.975 90.195 ;
        RECT -162.485 90.180 -162.055 90.195 ;
        RECT -152.565 90.180 -152.135 90.195 ;
        RECT -142.645 90.180 -142.215 90.195 ;
        RECT -132.725 90.180 -132.295 90.195 ;
        RECT -122.805 90.180 -122.375 90.195 ;
        RECT -112.885 90.180 -112.455 90.195 ;
        RECT -102.965 90.180 -102.535 90.195 ;
        RECT -93.045 90.180 -92.615 90.195 ;
        RECT -83.125 90.180 -82.695 90.195 ;
        RECT -73.205 90.180 -72.775 90.195 ;
        RECT -63.285 90.180 -62.855 90.195 ;
        RECT -53.365 90.180 -52.935 90.195 ;
        RECT -43.445 90.180 -43.015 90.195 ;
        RECT -33.525 90.180 -33.095 90.195 ;
        RECT -23.605 90.180 -23.175 90.195 ;
        RECT -13.685 90.180 -13.255 90.195 ;
        RECT -3.765 90.180 -3.335 90.195 ;
        RECT 6.155 90.180 6.585 90.195 ;
        RECT 16.075 90.180 16.505 90.195 ;
        RECT -283.360 90.175 -279.420 90.180 ;
        RECT -273.400 90.175 -269.380 90.180 ;
        RECT -263.520 90.175 -259.580 90.180 ;
        RECT -283.965 88.820 -278.655 90.175 ;
        RECT -283.965 88.805 -283.185 88.820 ;
        RECT -279.435 88.805 -278.655 88.820 ;
        RECT -274.045 88.805 -268.735 90.175 ;
        RECT -264.125 88.820 -258.815 90.175 ;
        RECT -264.125 88.805 -263.345 88.820 ;
        RECT -259.595 88.805 -258.815 88.820 ;
        RECT -254.205 90.170 -253.425 90.175 ;
        RECT -253.360 90.170 -249.910 90.180 ;
        RECT -243.680 90.175 -239.740 90.180 ;
        RECT -233.720 90.175 -229.700 90.180 ;
        RECT -223.840 90.175 -219.900 90.180 ;
        RECT -213.840 90.175 -209.770 90.180 ;
        RECT -204.000 90.175 -200.060 90.180 ;
        RECT -194.040 90.175 -190.020 90.180 ;
        RECT -184.160 90.175 -180.220 90.180 ;
        RECT -249.675 90.170 -248.895 90.175 ;
        RECT -254.205 88.805 -248.895 90.170 ;
        RECT -244.285 88.820 -238.975 90.175 ;
        RECT -244.285 88.805 -243.505 88.820 ;
        RECT -239.755 88.805 -238.975 88.820 ;
        RECT -234.365 88.805 -229.055 90.175 ;
        RECT -224.445 88.820 -219.135 90.175 ;
        RECT -224.445 88.805 -223.665 88.820 ;
        RECT -219.915 88.805 -219.135 88.820 ;
        RECT -214.525 88.810 -209.215 90.175 ;
        RECT -214.525 88.805 -213.745 88.810 ;
        RECT -209.995 88.805 -209.215 88.810 ;
        RECT -204.605 88.820 -199.295 90.175 ;
        RECT -204.605 88.805 -203.825 88.820 ;
        RECT -200.075 88.805 -199.295 88.820 ;
        RECT -194.685 88.805 -189.375 90.175 ;
        RECT -184.765 88.820 -179.455 90.175 ;
        RECT -184.765 88.805 -183.985 88.820 ;
        RECT -180.235 88.805 -179.455 88.820 ;
        RECT -174.845 90.170 -174.065 90.175 ;
        RECT -174.000 90.170 -170.550 90.180 ;
        RECT -164.320 90.175 -160.380 90.180 ;
        RECT -154.360 90.175 -150.340 90.180 ;
        RECT -144.480 90.175 -140.540 90.180 ;
        RECT -134.440 90.175 -130.500 90.180 ;
        RECT -124.640 90.175 -120.700 90.180 ;
        RECT -114.680 90.175 -110.660 90.180 ;
        RECT -104.800 90.175 -100.860 90.180 ;
        RECT -170.315 90.170 -169.535 90.175 ;
        RECT -174.845 88.805 -169.535 90.170 ;
        RECT -164.925 88.820 -159.615 90.175 ;
        RECT -164.925 88.805 -164.145 88.820 ;
        RECT -160.395 88.805 -159.615 88.820 ;
        RECT -155.005 88.805 -149.695 90.175 ;
        RECT -145.085 88.820 -139.775 90.175 ;
        RECT -145.085 88.805 -144.305 88.820 ;
        RECT -140.555 88.805 -139.775 88.820 ;
        RECT -135.165 88.820 -129.855 90.175 ;
        RECT -135.165 88.805 -134.385 88.820 ;
        RECT -130.635 88.805 -129.855 88.820 ;
        RECT -125.245 88.820 -119.935 90.175 ;
        RECT -125.245 88.805 -124.465 88.820 ;
        RECT -120.715 88.805 -119.935 88.820 ;
        RECT -115.325 88.805 -110.015 90.175 ;
        RECT -105.405 88.820 -100.095 90.175 ;
        RECT -105.405 88.805 -104.625 88.820 ;
        RECT -100.875 88.805 -100.095 88.820 ;
        RECT -95.485 90.170 -94.705 90.175 ;
        RECT -94.640 90.170 -91.190 90.180 ;
        RECT -84.960 90.175 -81.020 90.180 ;
        RECT -75.000 90.175 -70.980 90.180 ;
        RECT -65.120 90.175 -61.180 90.180 ;
        RECT -55.120 90.175 -51.050 90.180 ;
        RECT -45.280 90.175 -41.340 90.180 ;
        RECT -35.320 90.175 -31.300 90.180 ;
        RECT -25.440 90.175 -21.500 90.180 ;
        RECT -90.955 90.170 -90.175 90.175 ;
        RECT -95.485 88.805 -90.175 90.170 ;
        RECT -85.565 88.820 -80.255 90.175 ;
        RECT -85.565 88.805 -84.785 88.820 ;
        RECT -81.035 88.805 -80.255 88.820 ;
        RECT -75.645 88.805 -70.335 90.175 ;
        RECT -65.725 88.820 -60.415 90.175 ;
        RECT -65.725 88.805 -64.945 88.820 ;
        RECT -61.195 88.805 -60.415 88.820 ;
        RECT -55.805 88.810 -50.495 90.175 ;
        RECT -55.805 88.805 -55.025 88.810 ;
        RECT -51.275 88.805 -50.495 88.810 ;
        RECT -45.885 88.820 -40.575 90.175 ;
        RECT -45.885 88.805 -45.105 88.820 ;
        RECT -41.355 88.805 -40.575 88.820 ;
        RECT -35.965 88.805 -30.655 90.175 ;
        RECT -26.045 88.820 -20.735 90.175 ;
        RECT -26.045 88.805 -25.265 88.820 ;
        RECT -21.515 88.805 -20.735 88.820 ;
        RECT -16.125 90.170 -15.345 90.175 ;
        RECT -15.280 90.170 -11.830 90.180 ;
        RECT -5.600 90.175 -1.660 90.180 ;
        RECT 4.360 90.175 8.380 90.180 ;
        RECT 14.240 90.175 18.180 90.180 ;
        RECT -11.595 90.170 -10.815 90.175 ;
        RECT -16.125 88.805 -10.815 90.170 ;
        RECT -6.205 88.820 -0.895 90.175 ;
        RECT -6.205 88.805 -5.425 88.820 ;
        RECT -1.675 88.805 -0.895 88.820 ;
        RECT 3.715 88.805 9.025 90.175 ;
        RECT 13.635 88.820 18.945 90.175 ;
        RECT 13.635 88.805 14.415 88.820 ;
        RECT 18.165 88.805 18.945 88.820 ;
        RECT -273.400 88.800 -269.380 88.805 ;
        RECT -253.480 88.800 -249.640 88.805 ;
        RECT -233.720 88.800 -229.700 88.805 ;
        RECT -194.040 88.800 -190.020 88.805 ;
        RECT -174.120 88.800 -170.280 88.805 ;
        RECT -154.360 88.800 -150.340 88.805 ;
        RECT -114.680 88.800 -110.660 88.805 ;
        RECT -94.760 88.800 -90.920 88.805 ;
        RECT -75.000 88.800 -70.980 88.805 ;
        RECT -35.320 88.800 -31.300 88.805 ;
        RECT -15.400 88.800 -11.560 88.805 ;
        RECT 4.360 88.800 8.380 88.805 ;
      LAYER li1 ;
        RECT -288.125 94.615 -287.955 95.140 ;
        RECT -286.500 94.725 -286.040 94.895 ;
        RECT -288.505 94.285 -287.955 94.615 ;
        RECT -288.125 93.760 -287.955 94.285 ;
        RECT -286.415 94.000 -286.125 94.725 ;
        RECT -284.585 94.615 -284.415 95.140 ;
        RECT -278.205 94.615 -278.035 95.140 ;
        RECT -276.580 94.725 -276.120 94.895 ;
        RECT -284.585 94.285 -284.035 94.615 ;
        RECT -278.585 94.285 -278.035 94.615 ;
        RECT -284.585 93.760 -284.415 94.285 ;
        RECT -278.205 93.760 -278.035 94.285 ;
        RECT -276.495 94.000 -276.205 94.725 ;
        RECT -274.665 94.615 -274.495 95.140 ;
        RECT -268.285 94.615 -268.115 95.140 ;
        RECT -266.660 94.725 -266.200 94.895 ;
        RECT -274.665 94.285 -274.115 94.615 ;
        RECT -268.665 94.285 -268.115 94.615 ;
        RECT -274.665 93.760 -274.495 94.285 ;
        RECT -268.285 93.760 -268.115 94.285 ;
        RECT -266.575 94.000 -266.285 94.725 ;
        RECT -264.745 94.615 -264.575 95.140 ;
        RECT -258.365 94.615 -258.195 95.140 ;
        RECT -256.740 94.725 -256.280 94.895 ;
        RECT -264.745 94.285 -264.195 94.615 ;
        RECT -258.745 94.285 -258.195 94.615 ;
        RECT -264.745 93.760 -264.575 94.285 ;
        RECT -258.365 93.760 -258.195 94.285 ;
        RECT -256.655 94.000 -256.365 94.725 ;
        RECT -254.825 94.615 -254.655 95.140 ;
        RECT -248.445 94.615 -248.275 95.140 ;
        RECT -246.820 94.725 -246.360 94.895 ;
        RECT -254.825 94.285 -254.275 94.615 ;
        RECT -248.825 94.285 -248.275 94.615 ;
        RECT -254.825 93.760 -254.655 94.285 ;
        RECT -248.445 93.760 -248.275 94.285 ;
        RECT -246.735 94.000 -246.445 94.725 ;
        RECT -244.905 94.615 -244.735 95.140 ;
        RECT -238.525 94.615 -238.355 95.140 ;
        RECT -236.900 94.725 -236.440 94.895 ;
        RECT -244.905 94.285 -244.355 94.615 ;
        RECT -238.905 94.285 -238.355 94.615 ;
        RECT -244.905 93.760 -244.735 94.285 ;
        RECT -238.525 93.760 -238.355 94.285 ;
        RECT -236.815 94.000 -236.525 94.725 ;
        RECT -234.985 94.615 -234.815 95.140 ;
        RECT -228.605 94.615 -228.435 95.140 ;
        RECT -226.980 94.725 -226.520 94.895 ;
        RECT -234.985 94.285 -234.435 94.615 ;
        RECT -228.985 94.285 -228.435 94.615 ;
        RECT -234.985 93.760 -234.815 94.285 ;
        RECT -228.605 93.760 -228.435 94.285 ;
        RECT -226.895 94.000 -226.605 94.725 ;
        RECT -225.065 94.615 -224.895 95.140 ;
        RECT -218.685 94.615 -218.515 95.140 ;
        RECT -217.060 94.725 -216.600 94.895 ;
        RECT -225.065 94.285 -224.515 94.615 ;
        RECT -219.065 94.285 -218.515 94.615 ;
        RECT -225.065 93.760 -224.895 94.285 ;
        RECT -218.685 93.760 -218.515 94.285 ;
        RECT -216.975 94.000 -216.685 94.725 ;
        RECT -215.145 94.615 -214.975 95.140 ;
        RECT -208.765 94.615 -208.595 95.140 ;
        RECT -207.140 94.725 -206.680 94.895 ;
        RECT -215.145 94.285 -214.595 94.615 ;
        RECT -209.145 94.285 -208.595 94.615 ;
        RECT -215.145 93.760 -214.975 94.285 ;
        RECT -208.765 93.760 -208.595 94.285 ;
        RECT -207.055 94.000 -206.765 94.725 ;
        RECT -205.225 94.615 -205.055 95.140 ;
        RECT -198.845 94.615 -198.675 95.140 ;
        RECT -197.220 94.725 -196.760 94.895 ;
        RECT -205.225 94.285 -204.675 94.615 ;
        RECT -199.225 94.285 -198.675 94.615 ;
        RECT -205.225 93.760 -205.055 94.285 ;
        RECT -198.845 93.760 -198.675 94.285 ;
        RECT -197.135 94.000 -196.845 94.725 ;
        RECT -195.305 94.615 -195.135 95.140 ;
        RECT -188.925 94.615 -188.755 95.140 ;
        RECT -187.300 94.725 -186.840 94.895 ;
        RECT -195.305 94.285 -194.755 94.615 ;
        RECT -189.305 94.285 -188.755 94.615 ;
        RECT -195.305 93.760 -195.135 94.285 ;
        RECT -188.925 93.760 -188.755 94.285 ;
        RECT -187.215 94.000 -186.925 94.725 ;
        RECT -185.385 94.615 -185.215 95.140 ;
        RECT -179.005 94.615 -178.835 95.140 ;
        RECT -177.380 94.725 -176.920 94.895 ;
        RECT -185.385 94.285 -184.835 94.615 ;
        RECT -179.385 94.285 -178.835 94.615 ;
        RECT -185.385 93.760 -185.215 94.285 ;
        RECT -179.005 93.760 -178.835 94.285 ;
        RECT -177.295 94.000 -177.005 94.725 ;
        RECT -175.465 94.615 -175.295 95.140 ;
        RECT -169.085 94.615 -168.915 95.140 ;
        RECT -167.460 94.725 -167.000 94.895 ;
        RECT -175.465 94.285 -174.915 94.615 ;
        RECT -169.465 94.285 -168.915 94.615 ;
        RECT -175.465 93.760 -175.295 94.285 ;
        RECT -169.085 93.760 -168.915 94.285 ;
        RECT -167.375 94.000 -167.085 94.725 ;
        RECT -165.545 94.615 -165.375 95.140 ;
        RECT -159.165 94.615 -158.995 95.140 ;
        RECT -157.540 94.725 -157.080 94.895 ;
        RECT -165.545 94.285 -164.995 94.615 ;
        RECT -159.545 94.285 -158.995 94.615 ;
        RECT -165.545 93.760 -165.375 94.285 ;
        RECT -159.165 93.760 -158.995 94.285 ;
        RECT -157.455 94.000 -157.165 94.725 ;
        RECT -155.625 94.615 -155.455 95.140 ;
        RECT -149.245 94.615 -149.075 95.140 ;
        RECT -147.620 94.725 -147.160 94.895 ;
        RECT -155.625 94.285 -155.075 94.615 ;
        RECT -149.625 94.285 -149.075 94.615 ;
        RECT -155.625 93.760 -155.455 94.285 ;
        RECT -149.245 93.760 -149.075 94.285 ;
        RECT -147.535 94.000 -147.245 94.725 ;
        RECT -145.705 94.615 -145.535 95.140 ;
        RECT -139.325 94.615 -139.155 95.140 ;
        RECT -137.700 94.725 -137.240 94.895 ;
        RECT -145.705 94.285 -145.155 94.615 ;
        RECT -139.705 94.285 -139.155 94.615 ;
        RECT -145.705 93.760 -145.535 94.285 ;
        RECT -139.325 93.760 -139.155 94.285 ;
        RECT -137.615 94.000 -137.325 94.725 ;
        RECT -135.785 94.615 -135.615 95.140 ;
        RECT -129.405 94.615 -129.235 95.140 ;
        RECT -127.780 94.725 -127.320 94.895 ;
        RECT -135.785 94.285 -135.235 94.615 ;
        RECT -129.785 94.285 -129.235 94.615 ;
        RECT -135.785 93.760 -135.615 94.285 ;
        RECT -129.405 93.760 -129.235 94.285 ;
        RECT -127.695 94.000 -127.405 94.725 ;
        RECT -125.865 94.615 -125.695 95.140 ;
        RECT -119.485 94.615 -119.315 95.140 ;
        RECT -117.860 94.725 -117.400 94.895 ;
        RECT -125.865 94.285 -125.315 94.615 ;
        RECT -119.865 94.285 -119.315 94.615 ;
        RECT -125.865 93.760 -125.695 94.285 ;
        RECT -119.485 93.760 -119.315 94.285 ;
        RECT -117.775 94.000 -117.485 94.725 ;
        RECT -115.945 94.615 -115.775 95.140 ;
        RECT -109.565 94.615 -109.395 95.140 ;
        RECT -107.940 94.725 -107.480 94.895 ;
        RECT -115.945 94.285 -115.395 94.615 ;
        RECT -109.945 94.285 -109.395 94.615 ;
        RECT -115.945 93.760 -115.775 94.285 ;
        RECT -109.565 93.760 -109.395 94.285 ;
        RECT -107.855 94.000 -107.565 94.725 ;
        RECT -106.025 94.615 -105.855 95.140 ;
        RECT -99.645 94.615 -99.475 95.140 ;
        RECT -98.020 94.725 -97.560 94.895 ;
        RECT -106.025 94.285 -105.475 94.615 ;
        RECT -100.025 94.285 -99.475 94.615 ;
        RECT -106.025 93.760 -105.855 94.285 ;
        RECT -99.645 93.760 -99.475 94.285 ;
        RECT -97.935 94.000 -97.645 94.725 ;
        RECT -96.105 94.615 -95.935 95.140 ;
        RECT -89.725 94.615 -89.555 95.140 ;
        RECT -88.100 94.725 -87.640 94.895 ;
        RECT -96.105 94.285 -95.555 94.615 ;
        RECT -90.105 94.285 -89.555 94.615 ;
        RECT -96.105 93.760 -95.935 94.285 ;
        RECT -89.725 93.760 -89.555 94.285 ;
        RECT -88.015 94.000 -87.725 94.725 ;
        RECT -86.185 94.615 -86.015 95.140 ;
        RECT -79.805 94.615 -79.635 95.140 ;
        RECT -78.180 94.725 -77.720 94.895 ;
        RECT -86.185 94.285 -85.635 94.615 ;
        RECT -80.185 94.285 -79.635 94.615 ;
        RECT -86.185 93.760 -86.015 94.285 ;
        RECT -79.805 93.760 -79.635 94.285 ;
        RECT -78.095 94.000 -77.805 94.725 ;
        RECT -76.265 94.615 -76.095 95.140 ;
        RECT -69.885 94.615 -69.715 95.140 ;
        RECT -68.260 94.725 -67.800 94.895 ;
        RECT -76.265 94.285 -75.715 94.615 ;
        RECT -70.265 94.285 -69.715 94.615 ;
        RECT -76.265 93.760 -76.095 94.285 ;
        RECT -69.885 93.760 -69.715 94.285 ;
        RECT -68.175 94.000 -67.885 94.725 ;
        RECT -66.345 94.615 -66.175 95.140 ;
        RECT -59.965 94.615 -59.795 95.140 ;
        RECT -58.340 94.725 -57.880 94.895 ;
        RECT -66.345 94.285 -65.795 94.615 ;
        RECT -60.345 94.285 -59.795 94.615 ;
        RECT -66.345 93.760 -66.175 94.285 ;
        RECT -59.965 93.760 -59.795 94.285 ;
        RECT -58.255 94.000 -57.965 94.725 ;
        RECT -56.425 94.615 -56.255 95.140 ;
        RECT -50.045 94.615 -49.875 95.140 ;
        RECT -48.420 94.725 -47.960 94.895 ;
        RECT -56.425 94.285 -55.875 94.615 ;
        RECT -50.425 94.285 -49.875 94.615 ;
        RECT -56.425 93.760 -56.255 94.285 ;
        RECT -50.045 93.760 -49.875 94.285 ;
        RECT -48.335 94.000 -48.045 94.725 ;
        RECT -46.505 94.615 -46.335 95.140 ;
        RECT -40.125 94.615 -39.955 95.140 ;
        RECT -38.500 94.725 -38.040 94.895 ;
        RECT -46.505 94.285 -45.955 94.615 ;
        RECT -40.505 94.285 -39.955 94.615 ;
        RECT -46.505 93.760 -46.335 94.285 ;
        RECT -40.125 93.760 -39.955 94.285 ;
        RECT -38.415 94.000 -38.125 94.725 ;
        RECT -36.585 94.615 -36.415 95.140 ;
        RECT -30.205 94.615 -30.035 95.140 ;
        RECT -28.580 94.725 -28.120 94.895 ;
        RECT -36.585 94.285 -36.035 94.615 ;
        RECT -30.585 94.285 -30.035 94.615 ;
        RECT -36.585 93.760 -36.415 94.285 ;
        RECT -30.205 93.760 -30.035 94.285 ;
        RECT -28.495 94.000 -28.205 94.725 ;
        RECT -26.665 94.615 -26.495 95.140 ;
        RECT -20.285 94.615 -20.115 95.140 ;
        RECT -18.660 94.725 -18.200 94.895 ;
        RECT -26.665 94.285 -26.115 94.615 ;
        RECT -20.665 94.285 -20.115 94.615 ;
        RECT -26.665 93.760 -26.495 94.285 ;
        RECT -20.285 93.760 -20.115 94.285 ;
        RECT -18.575 94.000 -18.285 94.725 ;
        RECT -16.745 94.615 -16.575 95.140 ;
        RECT -10.365 94.615 -10.195 95.140 ;
        RECT -8.740 94.725 -8.280 94.895 ;
        RECT -16.745 94.285 -16.195 94.615 ;
        RECT -10.745 94.285 -10.195 94.615 ;
        RECT -16.745 93.760 -16.575 94.285 ;
        RECT -10.365 93.760 -10.195 94.285 ;
        RECT -8.655 94.000 -8.365 94.725 ;
        RECT -6.825 94.615 -6.655 95.140 ;
        RECT -0.445 94.615 -0.275 95.140 ;
        RECT 1.180 94.725 1.640 94.895 ;
        RECT -6.825 94.285 -6.275 94.615 ;
        RECT -0.825 94.285 -0.275 94.615 ;
        RECT -6.825 93.760 -6.655 94.285 ;
        RECT -0.445 93.760 -0.275 94.285 ;
        RECT 1.265 94.000 1.555 94.725 ;
        RECT 3.095 94.615 3.265 95.140 ;
        RECT 9.475 94.615 9.645 95.140 ;
        RECT 11.100 94.725 11.560 94.895 ;
        RECT 3.095 94.285 3.645 94.615 ;
        RECT 9.095 94.285 9.645 94.615 ;
        RECT 3.095 93.760 3.265 94.285 ;
        RECT 9.475 93.760 9.645 94.285 ;
        RECT 11.185 94.000 11.475 94.725 ;
        RECT 13.015 94.615 13.185 95.140 ;
        RECT 19.395 94.615 19.565 95.140 ;
        RECT 21.020 94.725 21.480 94.895 ;
        RECT 13.015 94.285 13.565 94.615 ;
        RECT 19.015 94.285 19.565 94.615 ;
        RECT 13.015 93.760 13.185 94.285 ;
        RECT 19.395 93.760 19.565 94.285 ;
        RECT 21.105 94.000 21.395 94.725 ;
        RECT 22.935 94.615 23.105 95.140 ;
        RECT 22.935 94.285 23.485 94.615 ;
        RECT 22.935 93.760 23.105 94.285 ;
        RECT -282.920 93.245 -279.700 93.415 ;
        RECT -273.000 93.245 -269.780 93.415 ;
        RECT -263.080 93.245 -259.860 93.415 ;
        RECT -253.160 93.245 -249.940 93.415 ;
        RECT -243.240 93.245 -240.020 93.415 ;
        RECT -233.320 93.245 -230.100 93.415 ;
        RECT -223.400 93.245 -220.180 93.415 ;
        RECT -213.480 93.245 -210.260 93.415 ;
        RECT -203.560 93.245 -200.340 93.415 ;
        RECT -193.640 93.245 -190.420 93.415 ;
        RECT -183.720 93.245 -180.500 93.415 ;
        RECT -173.800 93.245 -170.580 93.415 ;
        RECT -163.880 93.245 -160.660 93.415 ;
        RECT -153.960 93.245 -150.740 93.415 ;
        RECT -144.040 93.245 -140.820 93.415 ;
        RECT -134.120 93.245 -130.900 93.415 ;
        RECT -124.200 93.245 -120.980 93.415 ;
        RECT -114.280 93.245 -111.060 93.415 ;
        RECT -104.360 93.245 -101.140 93.415 ;
        RECT -94.440 93.245 -91.220 93.415 ;
        RECT -84.520 93.245 -81.300 93.415 ;
        RECT -74.600 93.245 -71.380 93.415 ;
        RECT -64.680 93.245 -61.460 93.415 ;
        RECT -54.760 93.245 -51.540 93.415 ;
        RECT -44.840 93.245 -41.620 93.415 ;
        RECT -34.920 93.245 -31.700 93.415 ;
        RECT -25.000 93.245 -21.780 93.415 ;
        RECT -15.080 93.245 -11.860 93.415 ;
        RECT -5.160 93.245 -1.940 93.415 ;
        RECT 4.760 93.245 7.980 93.415 ;
        RECT 14.680 93.245 17.900 93.415 ;
        RECT -281.935 92.445 -281.625 93.245 ;
        RECT -281.455 92.520 -281.165 93.245 ;
        RECT -280.995 92.445 -280.685 93.245 ;
        RECT -272.015 92.445 -271.705 93.245 ;
        RECT -271.535 92.520 -271.245 93.245 ;
        RECT -271.075 92.445 -270.765 93.245 ;
        RECT -262.095 92.445 -261.785 93.245 ;
        RECT -261.615 92.520 -261.325 93.245 ;
        RECT -261.155 92.445 -260.845 93.245 ;
        RECT -252.175 92.445 -251.865 93.245 ;
        RECT -251.695 92.520 -251.405 93.245 ;
        RECT -251.235 92.445 -250.925 93.245 ;
        RECT -242.255 92.445 -241.945 93.245 ;
        RECT -241.775 92.520 -241.485 93.245 ;
        RECT -241.315 92.445 -241.005 93.245 ;
        RECT -232.335 92.445 -232.025 93.245 ;
        RECT -231.855 92.520 -231.565 93.245 ;
        RECT -231.395 92.445 -231.085 93.245 ;
        RECT -222.415 92.445 -222.105 93.245 ;
        RECT -221.935 92.520 -221.645 93.245 ;
        RECT -221.475 92.445 -221.165 93.245 ;
        RECT -212.495 92.445 -212.185 93.245 ;
        RECT -212.015 92.520 -211.725 93.245 ;
        RECT -211.555 92.445 -211.245 93.245 ;
        RECT -202.575 92.445 -202.265 93.245 ;
        RECT -202.095 92.520 -201.805 93.245 ;
        RECT -201.635 92.445 -201.325 93.245 ;
        RECT -192.655 92.445 -192.345 93.245 ;
        RECT -192.175 92.520 -191.885 93.245 ;
        RECT -191.715 92.445 -191.405 93.245 ;
        RECT -182.735 92.445 -182.425 93.245 ;
        RECT -182.255 92.520 -181.965 93.245 ;
        RECT -181.795 92.445 -181.485 93.245 ;
        RECT -172.815 92.445 -172.505 93.245 ;
        RECT -172.335 92.520 -172.045 93.245 ;
        RECT -171.875 92.445 -171.565 93.245 ;
        RECT -162.895 92.445 -162.585 93.245 ;
        RECT -162.415 92.520 -162.125 93.245 ;
        RECT -161.955 92.445 -161.645 93.245 ;
        RECT -152.975 92.445 -152.665 93.245 ;
        RECT -152.495 92.520 -152.205 93.245 ;
        RECT -152.035 92.445 -151.725 93.245 ;
        RECT -143.055 92.445 -142.745 93.245 ;
        RECT -142.575 92.520 -142.285 93.245 ;
        RECT -142.115 92.445 -141.805 93.245 ;
        RECT -133.135 92.445 -132.825 93.245 ;
        RECT -132.655 92.520 -132.365 93.245 ;
        RECT -132.195 92.445 -131.885 93.245 ;
        RECT -123.215 92.445 -122.905 93.245 ;
        RECT -122.735 92.520 -122.445 93.245 ;
        RECT -122.275 92.445 -121.965 93.245 ;
        RECT -113.295 92.445 -112.985 93.245 ;
        RECT -112.815 92.520 -112.525 93.245 ;
        RECT -112.355 92.445 -112.045 93.245 ;
        RECT -103.375 92.445 -103.065 93.245 ;
        RECT -102.895 92.520 -102.605 93.245 ;
        RECT -102.435 92.445 -102.125 93.245 ;
        RECT -93.455 92.445 -93.145 93.245 ;
        RECT -92.975 92.520 -92.685 93.245 ;
        RECT -92.515 92.445 -92.205 93.245 ;
        RECT -83.535 92.445 -83.225 93.245 ;
        RECT -83.055 92.520 -82.765 93.245 ;
        RECT -82.595 92.445 -82.285 93.245 ;
        RECT -73.615 92.445 -73.305 93.245 ;
        RECT -73.135 92.520 -72.845 93.245 ;
        RECT -72.675 92.445 -72.365 93.245 ;
        RECT -63.695 92.445 -63.385 93.245 ;
        RECT -63.215 92.520 -62.925 93.245 ;
        RECT -62.755 92.445 -62.445 93.245 ;
        RECT -53.775 92.445 -53.465 93.245 ;
        RECT -53.295 92.520 -53.005 93.245 ;
        RECT -52.835 92.445 -52.525 93.245 ;
        RECT -43.855 92.445 -43.545 93.245 ;
        RECT -43.375 92.520 -43.085 93.245 ;
        RECT -42.915 92.445 -42.605 93.245 ;
        RECT -33.935 92.445 -33.625 93.245 ;
        RECT -33.455 92.520 -33.165 93.245 ;
        RECT -32.995 92.445 -32.685 93.245 ;
        RECT -24.015 92.445 -23.705 93.245 ;
        RECT -23.535 92.520 -23.245 93.245 ;
        RECT -23.075 92.445 -22.765 93.245 ;
        RECT -14.095 92.445 -13.785 93.245 ;
        RECT -13.615 92.520 -13.325 93.245 ;
        RECT -13.155 92.445 -12.845 93.245 ;
        RECT -4.175 92.445 -3.865 93.245 ;
        RECT -3.695 92.520 -3.405 93.245 ;
        RECT -3.235 92.445 -2.925 93.245 ;
        RECT 5.745 92.445 6.055 93.245 ;
        RECT 6.225 92.520 6.515 93.245 ;
        RECT 6.685 92.445 6.995 93.245 ;
        RECT 15.665 92.445 15.975 93.245 ;
        RECT 16.145 92.520 16.435 93.245 ;
        RECT 16.605 92.445 16.915 93.245 ;
        RECT -286.895 90.695 -286.585 91.495 ;
        RECT -286.415 90.695 -286.125 91.420 ;
        RECT -285.955 90.695 -285.645 91.495 ;
        RECT -276.975 90.695 -276.665 91.495 ;
        RECT -276.495 90.695 -276.205 91.420 ;
        RECT -276.035 90.695 -275.725 91.495 ;
        RECT -267.055 90.695 -266.745 91.495 ;
        RECT -266.575 90.695 -266.285 91.420 ;
        RECT -266.115 90.695 -265.805 91.495 ;
        RECT -257.135 90.695 -256.825 91.495 ;
        RECT -256.655 90.695 -256.365 91.420 ;
        RECT -256.195 90.695 -255.885 91.495 ;
        RECT -247.215 90.695 -246.905 91.495 ;
        RECT -246.735 90.695 -246.445 91.420 ;
        RECT -246.275 90.695 -245.965 91.495 ;
        RECT -237.295 90.695 -236.985 91.495 ;
        RECT -236.815 90.695 -236.525 91.420 ;
        RECT -236.355 90.695 -236.045 91.495 ;
        RECT -227.375 90.695 -227.065 91.495 ;
        RECT -226.895 90.695 -226.605 91.420 ;
        RECT -226.435 90.695 -226.125 91.495 ;
        RECT -217.455 90.695 -217.145 91.495 ;
        RECT -216.975 90.695 -216.685 91.420 ;
        RECT -216.515 90.695 -216.205 91.495 ;
        RECT -207.535 90.695 -207.225 91.495 ;
        RECT -207.055 90.695 -206.765 91.420 ;
        RECT -206.595 90.695 -206.285 91.495 ;
        RECT -197.615 90.695 -197.305 91.495 ;
        RECT -197.135 90.695 -196.845 91.420 ;
        RECT -196.675 90.695 -196.365 91.495 ;
        RECT -187.695 90.695 -187.385 91.495 ;
        RECT -187.215 90.695 -186.925 91.420 ;
        RECT -186.755 90.695 -186.445 91.495 ;
        RECT -177.775 90.695 -177.465 91.495 ;
        RECT -177.295 90.695 -177.005 91.420 ;
        RECT -176.835 90.695 -176.525 91.495 ;
        RECT -167.855 90.695 -167.545 91.495 ;
        RECT -167.375 90.695 -167.085 91.420 ;
        RECT -166.915 90.695 -166.605 91.495 ;
        RECT -157.935 90.695 -157.625 91.495 ;
        RECT -157.455 90.695 -157.165 91.420 ;
        RECT -156.995 90.695 -156.685 91.495 ;
        RECT -148.015 90.695 -147.705 91.495 ;
        RECT -147.535 90.695 -147.245 91.420 ;
        RECT -147.075 90.695 -146.765 91.495 ;
        RECT -138.095 90.695 -137.785 91.495 ;
        RECT -137.615 90.695 -137.325 91.420 ;
        RECT -137.155 90.695 -136.845 91.495 ;
        RECT -128.175 90.695 -127.865 91.495 ;
        RECT -127.695 90.695 -127.405 91.420 ;
        RECT -127.235 90.695 -126.925 91.495 ;
        RECT -118.255 90.695 -117.945 91.495 ;
        RECT -117.775 90.695 -117.485 91.420 ;
        RECT -117.315 90.695 -117.005 91.495 ;
        RECT -108.335 90.695 -108.025 91.495 ;
        RECT -107.855 90.695 -107.565 91.420 ;
        RECT -107.395 90.695 -107.085 91.495 ;
        RECT -98.415 90.695 -98.105 91.495 ;
        RECT -97.935 90.695 -97.645 91.420 ;
        RECT -97.475 90.695 -97.165 91.495 ;
        RECT -88.495 90.695 -88.185 91.495 ;
        RECT -88.015 90.695 -87.725 91.420 ;
        RECT -87.555 90.695 -87.245 91.495 ;
        RECT -78.575 90.695 -78.265 91.495 ;
        RECT -78.095 90.695 -77.805 91.420 ;
        RECT -77.635 90.695 -77.325 91.495 ;
        RECT -68.655 90.695 -68.345 91.495 ;
        RECT -68.175 90.695 -67.885 91.420 ;
        RECT -67.715 90.695 -67.405 91.495 ;
        RECT -58.735 90.695 -58.425 91.495 ;
        RECT -58.255 90.695 -57.965 91.420 ;
        RECT -57.795 90.695 -57.485 91.495 ;
        RECT -48.815 90.695 -48.505 91.495 ;
        RECT -48.335 90.695 -48.045 91.420 ;
        RECT -47.875 90.695 -47.565 91.495 ;
        RECT -38.895 90.695 -38.585 91.495 ;
        RECT -38.415 90.695 -38.125 91.420 ;
        RECT -37.955 90.695 -37.645 91.495 ;
        RECT -28.975 90.695 -28.665 91.495 ;
        RECT -28.495 90.695 -28.205 91.420 ;
        RECT -28.035 90.695 -27.725 91.495 ;
        RECT -19.055 90.695 -18.745 91.495 ;
        RECT -18.575 90.695 -18.285 91.420 ;
        RECT -18.115 90.695 -17.805 91.495 ;
        RECT -9.135 90.695 -8.825 91.495 ;
        RECT -8.655 90.695 -8.365 91.420 ;
        RECT -8.195 90.695 -7.885 91.495 ;
        RECT 0.785 90.695 1.095 91.495 ;
        RECT 1.265 90.695 1.555 91.420 ;
        RECT 1.725 90.695 2.035 91.495 ;
        RECT 10.705 90.695 11.015 91.495 ;
        RECT 11.185 90.695 11.475 91.420 ;
        RECT 11.645 90.695 11.955 91.495 ;
        RECT 20.625 90.695 20.935 91.495 ;
        RECT 21.105 90.695 21.395 91.420 ;
        RECT 21.565 90.695 21.875 91.495 ;
        RECT -287.880 90.525 -284.660 90.695 ;
        RECT -277.960 90.525 -274.740 90.695 ;
        RECT -268.040 90.525 -264.820 90.695 ;
        RECT -258.120 90.525 -254.900 90.695 ;
        RECT -248.200 90.525 -244.980 90.695 ;
        RECT -238.280 90.525 -235.060 90.695 ;
        RECT -228.360 90.525 -225.140 90.695 ;
        RECT -218.440 90.525 -215.220 90.695 ;
        RECT -208.520 90.525 -205.300 90.695 ;
        RECT -198.600 90.525 -195.380 90.695 ;
        RECT -188.680 90.525 -185.460 90.695 ;
        RECT -178.760 90.525 -175.540 90.695 ;
        RECT -168.840 90.525 -165.620 90.695 ;
        RECT -158.920 90.525 -155.700 90.695 ;
        RECT -149.000 90.525 -145.780 90.695 ;
        RECT -139.080 90.525 -135.860 90.695 ;
        RECT -129.160 90.525 -125.940 90.695 ;
        RECT -119.240 90.525 -116.020 90.695 ;
        RECT -109.320 90.525 -106.100 90.695 ;
        RECT -99.400 90.525 -96.180 90.695 ;
        RECT -89.480 90.525 -86.260 90.695 ;
        RECT -79.560 90.525 -76.340 90.695 ;
        RECT -69.640 90.525 -66.420 90.695 ;
        RECT -59.720 90.525 -56.500 90.695 ;
        RECT -49.800 90.525 -46.580 90.695 ;
        RECT -39.880 90.525 -36.660 90.695 ;
        RECT -29.960 90.525 -26.740 90.695 ;
        RECT -20.040 90.525 -16.820 90.695 ;
        RECT -10.120 90.525 -6.900 90.695 ;
        RECT -0.200 90.525 3.020 90.695 ;
        RECT 9.720 90.525 12.940 90.695 ;
        RECT 19.640 90.525 22.860 90.695 ;
        RECT -283.165 89.655 -282.995 90.180 ;
        RECT -283.545 89.325 -282.995 89.655 ;
        RECT -283.165 88.800 -282.995 89.325 ;
        RECT -281.455 89.305 -281.165 90.030 ;
        RECT -279.625 89.655 -279.455 90.180 ;
        RECT -273.245 89.655 -273.075 90.180 ;
        RECT -279.625 89.325 -279.075 89.655 ;
        RECT -273.625 89.325 -273.075 89.655 ;
        RECT -281.540 89.135 -281.080 89.305 ;
        RECT -279.625 88.800 -279.455 89.325 ;
        RECT -273.245 88.800 -273.075 89.325 ;
        RECT -271.535 89.305 -271.245 90.030 ;
        RECT -269.705 89.655 -269.535 90.180 ;
        RECT -263.325 89.655 -263.155 90.180 ;
        RECT -269.705 89.325 -269.155 89.655 ;
        RECT -263.705 89.325 -263.155 89.655 ;
        RECT -271.620 89.135 -271.160 89.305 ;
        RECT -269.705 88.800 -269.535 89.325 ;
        RECT -263.325 88.800 -263.155 89.325 ;
        RECT -261.615 89.305 -261.325 90.030 ;
        RECT -259.785 89.655 -259.615 90.180 ;
        RECT -253.405 89.655 -253.235 90.180 ;
        RECT -259.785 89.325 -259.235 89.655 ;
        RECT -253.785 89.325 -253.235 89.655 ;
        RECT -261.700 89.135 -261.240 89.305 ;
        RECT -259.785 88.800 -259.615 89.325 ;
        RECT -253.405 88.800 -253.235 89.325 ;
        RECT -251.695 89.305 -251.405 90.030 ;
        RECT -249.865 89.655 -249.695 90.180 ;
        RECT -243.485 89.655 -243.315 90.180 ;
        RECT -249.865 89.325 -249.315 89.655 ;
        RECT -243.865 89.325 -243.315 89.655 ;
        RECT -251.780 89.135 -251.320 89.305 ;
        RECT -249.865 88.800 -249.695 89.325 ;
        RECT -243.485 88.800 -243.315 89.325 ;
        RECT -241.775 89.305 -241.485 90.030 ;
        RECT -239.945 89.655 -239.775 90.180 ;
        RECT -233.565 89.655 -233.395 90.180 ;
        RECT -239.945 89.325 -239.395 89.655 ;
        RECT -233.945 89.325 -233.395 89.655 ;
        RECT -241.860 89.135 -241.400 89.305 ;
        RECT -239.945 88.800 -239.775 89.325 ;
        RECT -233.565 88.800 -233.395 89.325 ;
        RECT -231.855 89.305 -231.565 90.030 ;
        RECT -230.025 89.655 -229.855 90.180 ;
        RECT -223.645 89.655 -223.475 90.180 ;
        RECT -230.025 89.325 -229.475 89.655 ;
        RECT -224.025 89.325 -223.475 89.655 ;
        RECT -231.940 89.135 -231.480 89.305 ;
        RECT -230.025 88.800 -229.855 89.325 ;
        RECT -223.645 88.800 -223.475 89.325 ;
        RECT -221.935 89.305 -221.645 90.030 ;
        RECT -220.105 89.655 -219.935 90.180 ;
        RECT -213.725 89.655 -213.555 90.180 ;
        RECT -220.105 89.325 -219.555 89.655 ;
        RECT -214.105 89.325 -213.555 89.655 ;
        RECT -222.020 89.135 -221.560 89.305 ;
        RECT -220.105 88.800 -219.935 89.325 ;
        RECT -213.725 88.800 -213.555 89.325 ;
        RECT -212.015 89.305 -211.725 90.030 ;
        RECT -210.185 89.655 -210.015 90.180 ;
        RECT -203.805 89.655 -203.635 90.180 ;
        RECT -210.185 89.325 -209.635 89.655 ;
        RECT -204.185 89.325 -203.635 89.655 ;
        RECT -212.100 89.135 -211.640 89.305 ;
        RECT -210.185 88.800 -210.015 89.325 ;
        RECT -203.805 88.800 -203.635 89.325 ;
        RECT -202.095 89.305 -201.805 90.030 ;
        RECT -200.265 89.655 -200.095 90.180 ;
        RECT -193.885 89.655 -193.715 90.180 ;
        RECT -200.265 89.325 -199.715 89.655 ;
        RECT -194.265 89.325 -193.715 89.655 ;
        RECT -202.180 89.135 -201.720 89.305 ;
        RECT -200.265 88.800 -200.095 89.325 ;
        RECT -193.885 88.800 -193.715 89.325 ;
        RECT -192.175 89.305 -191.885 90.030 ;
        RECT -190.345 89.655 -190.175 90.180 ;
        RECT -183.965 89.655 -183.795 90.180 ;
        RECT -190.345 89.325 -189.795 89.655 ;
        RECT -184.345 89.325 -183.795 89.655 ;
        RECT -192.260 89.135 -191.800 89.305 ;
        RECT -190.345 88.800 -190.175 89.325 ;
        RECT -183.965 88.800 -183.795 89.325 ;
        RECT -182.255 89.305 -181.965 90.030 ;
        RECT -180.425 89.655 -180.255 90.180 ;
        RECT -174.045 89.655 -173.875 90.180 ;
        RECT -180.425 89.325 -179.875 89.655 ;
        RECT -174.425 89.325 -173.875 89.655 ;
        RECT -182.340 89.135 -181.880 89.305 ;
        RECT -180.425 88.800 -180.255 89.325 ;
        RECT -174.045 88.800 -173.875 89.325 ;
        RECT -172.335 89.305 -172.045 90.030 ;
        RECT -170.505 89.655 -170.335 90.180 ;
        RECT -164.125 89.655 -163.955 90.180 ;
        RECT -170.505 89.325 -169.955 89.655 ;
        RECT -164.505 89.325 -163.955 89.655 ;
        RECT -172.420 89.135 -171.960 89.305 ;
        RECT -170.505 88.800 -170.335 89.325 ;
        RECT -164.125 88.800 -163.955 89.325 ;
        RECT -162.415 89.305 -162.125 90.030 ;
        RECT -160.585 89.655 -160.415 90.180 ;
        RECT -154.205 89.655 -154.035 90.180 ;
        RECT -160.585 89.325 -160.035 89.655 ;
        RECT -154.585 89.325 -154.035 89.655 ;
        RECT -162.500 89.135 -162.040 89.305 ;
        RECT -160.585 88.800 -160.415 89.325 ;
        RECT -154.205 88.800 -154.035 89.325 ;
        RECT -152.495 89.305 -152.205 90.030 ;
        RECT -150.665 89.655 -150.495 90.180 ;
        RECT -144.285 89.655 -144.115 90.180 ;
        RECT -150.665 89.325 -150.115 89.655 ;
        RECT -144.665 89.325 -144.115 89.655 ;
        RECT -152.580 89.135 -152.120 89.305 ;
        RECT -150.665 88.800 -150.495 89.325 ;
        RECT -144.285 88.800 -144.115 89.325 ;
        RECT -142.575 89.305 -142.285 90.030 ;
        RECT -140.745 89.655 -140.575 90.180 ;
        RECT -134.365 89.655 -134.195 90.180 ;
        RECT -140.745 89.325 -140.195 89.655 ;
        RECT -134.745 89.325 -134.195 89.655 ;
        RECT -142.660 89.135 -142.200 89.305 ;
        RECT -140.745 88.800 -140.575 89.325 ;
        RECT -134.365 88.800 -134.195 89.325 ;
        RECT -132.655 89.305 -132.365 90.030 ;
        RECT -130.825 89.655 -130.655 90.180 ;
        RECT -124.445 89.655 -124.275 90.180 ;
        RECT -130.825 89.325 -130.275 89.655 ;
        RECT -124.825 89.325 -124.275 89.655 ;
        RECT -132.740 89.135 -132.280 89.305 ;
        RECT -130.825 88.800 -130.655 89.325 ;
        RECT -124.445 88.800 -124.275 89.325 ;
        RECT -122.735 89.305 -122.445 90.030 ;
        RECT -120.905 89.655 -120.735 90.180 ;
        RECT -114.525 89.655 -114.355 90.180 ;
        RECT -120.905 89.325 -120.355 89.655 ;
        RECT -114.905 89.325 -114.355 89.655 ;
        RECT -122.820 89.135 -122.360 89.305 ;
        RECT -120.905 88.800 -120.735 89.325 ;
        RECT -114.525 88.800 -114.355 89.325 ;
        RECT -112.815 89.305 -112.525 90.030 ;
        RECT -110.985 89.655 -110.815 90.180 ;
        RECT -104.605 89.655 -104.435 90.180 ;
        RECT -110.985 89.325 -110.435 89.655 ;
        RECT -104.985 89.325 -104.435 89.655 ;
        RECT -112.900 89.135 -112.440 89.305 ;
        RECT -110.985 88.800 -110.815 89.325 ;
        RECT -104.605 88.800 -104.435 89.325 ;
        RECT -102.895 89.305 -102.605 90.030 ;
        RECT -101.065 89.655 -100.895 90.180 ;
        RECT -94.685 89.655 -94.515 90.180 ;
        RECT -101.065 89.325 -100.515 89.655 ;
        RECT -95.065 89.325 -94.515 89.655 ;
        RECT -102.980 89.135 -102.520 89.305 ;
        RECT -101.065 88.800 -100.895 89.325 ;
        RECT -94.685 88.800 -94.515 89.325 ;
        RECT -92.975 89.305 -92.685 90.030 ;
        RECT -91.145 89.655 -90.975 90.180 ;
        RECT -84.765 89.655 -84.595 90.180 ;
        RECT -91.145 89.325 -90.595 89.655 ;
        RECT -85.145 89.325 -84.595 89.655 ;
        RECT -93.060 89.135 -92.600 89.305 ;
        RECT -91.145 88.800 -90.975 89.325 ;
        RECT -84.765 88.800 -84.595 89.325 ;
        RECT -83.055 89.305 -82.765 90.030 ;
        RECT -81.225 89.655 -81.055 90.180 ;
        RECT -74.845 89.655 -74.675 90.180 ;
        RECT -81.225 89.325 -80.675 89.655 ;
        RECT -75.225 89.325 -74.675 89.655 ;
        RECT -83.140 89.135 -82.680 89.305 ;
        RECT -81.225 88.800 -81.055 89.325 ;
        RECT -74.845 88.800 -74.675 89.325 ;
        RECT -73.135 89.305 -72.845 90.030 ;
        RECT -71.305 89.655 -71.135 90.180 ;
        RECT -64.925 89.655 -64.755 90.180 ;
        RECT -71.305 89.325 -70.755 89.655 ;
        RECT -65.305 89.325 -64.755 89.655 ;
        RECT -73.220 89.135 -72.760 89.305 ;
        RECT -71.305 88.800 -71.135 89.325 ;
        RECT -64.925 88.800 -64.755 89.325 ;
        RECT -63.215 89.305 -62.925 90.030 ;
        RECT -61.385 89.655 -61.215 90.180 ;
        RECT -55.005 89.655 -54.835 90.180 ;
        RECT -61.385 89.325 -60.835 89.655 ;
        RECT -55.385 89.325 -54.835 89.655 ;
        RECT -63.300 89.135 -62.840 89.305 ;
        RECT -61.385 88.800 -61.215 89.325 ;
        RECT -55.005 88.800 -54.835 89.325 ;
        RECT -53.295 89.305 -53.005 90.030 ;
        RECT -51.465 89.655 -51.295 90.180 ;
        RECT -45.085 89.655 -44.915 90.180 ;
        RECT -51.465 89.325 -50.915 89.655 ;
        RECT -45.465 89.325 -44.915 89.655 ;
        RECT -53.380 89.135 -52.920 89.305 ;
        RECT -51.465 88.800 -51.295 89.325 ;
        RECT -45.085 88.800 -44.915 89.325 ;
        RECT -43.375 89.305 -43.085 90.030 ;
        RECT -41.545 89.655 -41.375 90.180 ;
        RECT -35.165 89.655 -34.995 90.180 ;
        RECT -41.545 89.325 -40.995 89.655 ;
        RECT -35.545 89.325 -34.995 89.655 ;
        RECT -43.460 89.135 -43.000 89.305 ;
        RECT -41.545 88.800 -41.375 89.325 ;
        RECT -35.165 88.800 -34.995 89.325 ;
        RECT -33.455 89.305 -33.165 90.030 ;
        RECT -31.625 89.655 -31.455 90.180 ;
        RECT -25.245 89.655 -25.075 90.180 ;
        RECT -31.625 89.325 -31.075 89.655 ;
        RECT -25.625 89.325 -25.075 89.655 ;
        RECT -33.540 89.135 -33.080 89.305 ;
        RECT -31.625 88.800 -31.455 89.325 ;
        RECT -25.245 88.800 -25.075 89.325 ;
        RECT -23.535 89.305 -23.245 90.030 ;
        RECT -21.705 89.655 -21.535 90.180 ;
        RECT -15.325 89.655 -15.155 90.180 ;
        RECT -21.705 89.325 -21.155 89.655 ;
        RECT -15.705 89.325 -15.155 89.655 ;
        RECT -23.620 89.135 -23.160 89.305 ;
        RECT -21.705 88.800 -21.535 89.325 ;
        RECT -15.325 88.800 -15.155 89.325 ;
        RECT -13.615 89.305 -13.325 90.030 ;
        RECT -11.785 89.655 -11.615 90.180 ;
        RECT -5.405 89.655 -5.235 90.180 ;
        RECT -11.785 89.325 -11.235 89.655 ;
        RECT -5.785 89.325 -5.235 89.655 ;
        RECT -13.700 89.135 -13.240 89.305 ;
        RECT -11.785 88.800 -11.615 89.325 ;
        RECT -5.405 88.800 -5.235 89.325 ;
        RECT -3.695 89.305 -3.405 90.030 ;
        RECT -1.865 89.655 -1.695 90.180 ;
        RECT 4.515 89.655 4.685 90.180 ;
        RECT -1.865 89.325 -1.315 89.655 ;
        RECT 4.135 89.325 4.685 89.655 ;
        RECT -3.780 89.135 -3.320 89.305 ;
        RECT -1.865 88.800 -1.695 89.325 ;
        RECT 4.515 88.800 4.685 89.325 ;
        RECT 6.225 89.305 6.515 90.030 ;
        RECT 8.055 89.655 8.225 90.180 ;
        RECT 14.435 89.655 14.605 90.180 ;
        RECT 8.055 89.325 8.605 89.655 ;
        RECT 14.055 89.325 14.605 89.655 ;
        RECT 6.140 89.135 6.600 89.305 ;
        RECT 8.055 88.800 8.225 89.325 ;
        RECT 14.435 88.800 14.605 89.325 ;
        RECT 16.145 89.305 16.435 90.030 ;
        RECT 17.975 89.655 18.145 90.180 ;
        RECT 17.975 89.325 18.525 89.655 ;
        RECT 16.060 89.135 16.520 89.305 ;
        RECT 17.975 88.800 18.145 89.325 ;
      LAYER mcon ;
        RECT -288.125 94.825 -287.955 94.995 ;
        RECT -286.355 94.725 -286.185 94.895 ;
        RECT -284.585 94.825 -284.415 94.995 ;
        RECT -288.125 94.365 -287.955 94.535 ;
        RECT -288.125 93.905 -287.955 94.075 ;
        RECT -278.205 94.825 -278.035 94.995 ;
        RECT -276.435 94.725 -276.265 94.895 ;
        RECT -274.665 94.825 -274.495 94.995 ;
        RECT -284.585 94.365 -284.415 94.535 ;
        RECT -278.205 94.365 -278.035 94.535 ;
        RECT -284.585 93.905 -284.415 94.075 ;
        RECT -278.205 93.905 -278.035 94.075 ;
        RECT -268.285 94.825 -268.115 94.995 ;
        RECT -266.515 94.725 -266.345 94.895 ;
        RECT -264.745 94.825 -264.575 94.995 ;
        RECT -274.665 94.365 -274.495 94.535 ;
        RECT -268.285 94.365 -268.115 94.535 ;
        RECT -274.665 93.905 -274.495 94.075 ;
        RECT -268.285 93.905 -268.115 94.075 ;
        RECT -258.365 94.825 -258.195 94.995 ;
        RECT -256.595 94.725 -256.425 94.895 ;
        RECT -254.825 94.825 -254.655 94.995 ;
        RECT -264.745 94.365 -264.575 94.535 ;
        RECT -258.365 94.365 -258.195 94.535 ;
        RECT -264.745 93.905 -264.575 94.075 ;
        RECT -258.365 93.905 -258.195 94.075 ;
        RECT -248.445 94.825 -248.275 94.995 ;
        RECT -246.675 94.725 -246.505 94.895 ;
        RECT -244.905 94.825 -244.735 94.995 ;
        RECT -254.825 94.365 -254.655 94.535 ;
        RECT -248.445 94.365 -248.275 94.535 ;
        RECT -254.825 93.905 -254.655 94.075 ;
        RECT -248.445 93.905 -248.275 94.075 ;
        RECT -238.525 94.825 -238.355 94.995 ;
        RECT -236.755 94.725 -236.585 94.895 ;
        RECT -234.985 94.825 -234.815 94.995 ;
        RECT -244.905 94.365 -244.735 94.535 ;
        RECT -238.525 94.365 -238.355 94.535 ;
        RECT -244.905 93.905 -244.735 94.075 ;
        RECT -238.525 93.905 -238.355 94.075 ;
        RECT -228.605 94.825 -228.435 94.995 ;
        RECT -226.835 94.725 -226.665 94.895 ;
        RECT -225.065 94.825 -224.895 94.995 ;
        RECT -234.985 94.365 -234.815 94.535 ;
        RECT -228.605 94.365 -228.435 94.535 ;
        RECT -234.985 93.905 -234.815 94.075 ;
        RECT -228.605 93.905 -228.435 94.075 ;
        RECT -218.685 94.825 -218.515 94.995 ;
        RECT -216.915 94.725 -216.745 94.895 ;
        RECT -215.145 94.825 -214.975 94.995 ;
        RECT -225.065 94.365 -224.895 94.535 ;
        RECT -218.685 94.365 -218.515 94.535 ;
        RECT -225.065 93.905 -224.895 94.075 ;
        RECT -218.685 93.905 -218.515 94.075 ;
        RECT -208.765 94.825 -208.595 94.995 ;
        RECT -206.995 94.725 -206.825 94.895 ;
        RECT -205.225 94.825 -205.055 94.995 ;
        RECT -215.145 94.365 -214.975 94.535 ;
        RECT -208.765 94.365 -208.595 94.535 ;
        RECT -215.145 93.905 -214.975 94.075 ;
        RECT -208.765 93.905 -208.595 94.075 ;
        RECT -198.845 94.825 -198.675 94.995 ;
        RECT -197.075 94.725 -196.905 94.895 ;
        RECT -195.305 94.825 -195.135 94.995 ;
        RECT -205.225 94.365 -205.055 94.535 ;
        RECT -198.845 94.365 -198.675 94.535 ;
        RECT -205.225 93.905 -205.055 94.075 ;
        RECT -198.845 93.905 -198.675 94.075 ;
        RECT -188.925 94.825 -188.755 94.995 ;
        RECT -187.155 94.725 -186.985 94.895 ;
        RECT -185.385 94.825 -185.215 94.995 ;
        RECT -195.305 94.365 -195.135 94.535 ;
        RECT -188.925 94.365 -188.755 94.535 ;
        RECT -195.305 93.905 -195.135 94.075 ;
        RECT -188.925 93.905 -188.755 94.075 ;
        RECT -179.005 94.825 -178.835 94.995 ;
        RECT -177.235 94.725 -177.065 94.895 ;
        RECT -175.465 94.825 -175.295 94.995 ;
        RECT -185.385 94.365 -185.215 94.535 ;
        RECT -179.005 94.365 -178.835 94.535 ;
        RECT -185.385 93.905 -185.215 94.075 ;
        RECT -179.005 93.905 -178.835 94.075 ;
        RECT -169.085 94.825 -168.915 94.995 ;
        RECT -167.315 94.725 -167.145 94.895 ;
        RECT -165.545 94.825 -165.375 94.995 ;
        RECT -175.465 94.365 -175.295 94.535 ;
        RECT -169.085 94.365 -168.915 94.535 ;
        RECT -175.465 93.905 -175.295 94.075 ;
        RECT -169.085 93.905 -168.915 94.075 ;
        RECT -159.165 94.825 -158.995 94.995 ;
        RECT -157.395 94.725 -157.225 94.895 ;
        RECT -155.625 94.825 -155.455 94.995 ;
        RECT -165.545 94.365 -165.375 94.535 ;
        RECT -159.165 94.365 -158.995 94.535 ;
        RECT -165.545 93.905 -165.375 94.075 ;
        RECT -159.165 93.905 -158.995 94.075 ;
        RECT -149.245 94.825 -149.075 94.995 ;
        RECT -147.475 94.725 -147.305 94.895 ;
        RECT -145.705 94.825 -145.535 94.995 ;
        RECT -155.625 94.365 -155.455 94.535 ;
        RECT -149.245 94.365 -149.075 94.535 ;
        RECT -155.625 93.905 -155.455 94.075 ;
        RECT -149.245 93.905 -149.075 94.075 ;
        RECT -139.325 94.825 -139.155 94.995 ;
        RECT -137.555 94.725 -137.385 94.895 ;
        RECT -135.785 94.825 -135.615 94.995 ;
        RECT -145.705 94.365 -145.535 94.535 ;
        RECT -139.325 94.365 -139.155 94.535 ;
        RECT -145.705 93.905 -145.535 94.075 ;
        RECT -139.325 93.905 -139.155 94.075 ;
        RECT -129.405 94.825 -129.235 94.995 ;
        RECT -127.635 94.725 -127.465 94.895 ;
        RECT -125.865 94.825 -125.695 94.995 ;
        RECT -135.785 94.365 -135.615 94.535 ;
        RECT -129.405 94.365 -129.235 94.535 ;
        RECT -135.785 93.905 -135.615 94.075 ;
        RECT -129.405 93.905 -129.235 94.075 ;
        RECT -119.485 94.825 -119.315 94.995 ;
        RECT -117.715 94.725 -117.545 94.895 ;
        RECT -115.945 94.825 -115.775 94.995 ;
        RECT -125.865 94.365 -125.695 94.535 ;
        RECT -119.485 94.365 -119.315 94.535 ;
        RECT -125.865 93.905 -125.695 94.075 ;
        RECT -119.485 93.905 -119.315 94.075 ;
        RECT -109.565 94.825 -109.395 94.995 ;
        RECT -107.795 94.725 -107.625 94.895 ;
        RECT -106.025 94.825 -105.855 94.995 ;
        RECT -115.945 94.365 -115.775 94.535 ;
        RECT -109.565 94.365 -109.395 94.535 ;
        RECT -115.945 93.905 -115.775 94.075 ;
        RECT -109.565 93.905 -109.395 94.075 ;
        RECT -99.645 94.825 -99.475 94.995 ;
        RECT -97.875 94.725 -97.705 94.895 ;
        RECT -96.105 94.825 -95.935 94.995 ;
        RECT -106.025 94.365 -105.855 94.535 ;
        RECT -99.645 94.365 -99.475 94.535 ;
        RECT -106.025 93.905 -105.855 94.075 ;
        RECT -99.645 93.905 -99.475 94.075 ;
        RECT -89.725 94.825 -89.555 94.995 ;
        RECT -87.955 94.725 -87.785 94.895 ;
        RECT -86.185 94.825 -86.015 94.995 ;
        RECT -96.105 94.365 -95.935 94.535 ;
        RECT -89.725 94.365 -89.555 94.535 ;
        RECT -96.105 93.905 -95.935 94.075 ;
        RECT -89.725 93.905 -89.555 94.075 ;
        RECT -79.805 94.825 -79.635 94.995 ;
        RECT -78.035 94.725 -77.865 94.895 ;
        RECT -76.265 94.825 -76.095 94.995 ;
        RECT -86.185 94.365 -86.015 94.535 ;
        RECT -79.805 94.365 -79.635 94.535 ;
        RECT -86.185 93.905 -86.015 94.075 ;
        RECT -79.805 93.905 -79.635 94.075 ;
        RECT -69.885 94.825 -69.715 94.995 ;
        RECT -68.115 94.725 -67.945 94.895 ;
        RECT -66.345 94.825 -66.175 94.995 ;
        RECT -76.265 94.365 -76.095 94.535 ;
        RECT -69.885 94.365 -69.715 94.535 ;
        RECT -76.265 93.905 -76.095 94.075 ;
        RECT -69.885 93.905 -69.715 94.075 ;
        RECT -59.965 94.825 -59.795 94.995 ;
        RECT -58.195 94.725 -58.025 94.895 ;
        RECT -56.425 94.825 -56.255 94.995 ;
        RECT -66.345 94.365 -66.175 94.535 ;
        RECT -59.965 94.365 -59.795 94.535 ;
        RECT -66.345 93.905 -66.175 94.075 ;
        RECT -59.965 93.905 -59.795 94.075 ;
        RECT -50.045 94.825 -49.875 94.995 ;
        RECT -48.275 94.725 -48.105 94.895 ;
        RECT -46.505 94.825 -46.335 94.995 ;
        RECT -56.425 94.365 -56.255 94.535 ;
        RECT -50.045 94.365 -49.875 94.535 ;
        RECT -56.425 93.905 -56.255 94.075 ;
        RECT -50.045 93.905 -49.875 94.075 ;
        RECT -40.125 94.825 -39.955 94.995 ;
        RECT -38.355 94.725 -38.185 94.895 ;
        RECT -36.585 94.825 -36.415 94.995 ;
        RECT -46.505 94.365 -46.335 94.535 ;
        RECT -40.125 94.365 -39.955 94.535 ;
        RECT -46.505 93.905 -46.335 94.075 ;
        RECT -40.125 93.905 -39.955 94.075 ;
        RECT -30.205 94.825 -30.035 94.995 ;
        RECT -28.435 94.725 -28.265 94.895 ;
        RECT -26.665 94.825 -26.495 94.995 ;
        RECT -36.585 94.365 -36.415 94.535 ;
        RECT -30.205 94.365 -30.035 94.535 ;
        RECT -36.585 93.905 -36.415 94.075 ;
        RECT -30.205 93.905 -30.035 94.075 ;
        RECT -20.285 94.825 -20.115 94.995 ;
        RECT -18.515 94.725 -18.345 94.895 ;
        RECT -16.745 94.825 -16.575 94.995 ;
        RECT -26.665 94.365 -26.495 94.535 ;
        RECT -20.285 94.365 -20.115 94.535 ;
        RECT -26.665 93.905 -26.495 94.075 ;
        RECT -20.285 93.905 -20.115 94.075 ;
        RECT -10.365 94.825 -10.195 94.995 ;
        RECT -8.595 94.725 -8.425 94.895 ;
        RECT -6.825 94.825 -6.655 94.995 ;
        RECT -16.745 94.365 -16.575 94.535 ;
        RECT -10.365 94.365 -10.195 94.535 ;
        RECT -16.745 93.905 -16.575 94.075 ;
        RECT -10.365 93.905 -10.195 94.075 ;
        RECT -0.445 94.825 -0.275 94.995 ;
        RECT 1.325 94.725 1.495 94.895 ;
        RECT 3.095 94.825 3.265 94.995 ;
        RECT -6.825 94.365 -6.655 94.535 ;
        RECT -0.445 94.365 -0.275 94.535 ;
        RECT -6.825 93.905 -6.655 94.075 ;
        RECT -0.445 93.905 -0.275 94.075 ;
        RECT 9.475 94.825 9.645 94.995 ;
        RECT 11.245 94.725 11.415 94.895 ;
        RECT 13.015 94.825 13.185 94.995 ;
        RECT 3.095 94.365 3.265 94.535 ;
        RECT 9.475 94.365 9.645 94.535 ;
        RECT 3.095 93.905 3.265 94.075 ;
        RECT 9.475 93.905 9.645 94.075 ;
        RECT 19.395 94.825 19.565 94.995 ;
        RECT 21.165 94.725 21.335 94.895 ;
        RECT 22.935 94.825 23.105 94.995 ;
        RECT 13.015 94.365 13.185 94.535 ;
        RECT 19.395 94.365 19.565 94.535 ;
        RECT 13.015 93.905 13.185 94.075 ;
        RECT 19.395 93.905 19.565 94.075 ;
        RECT 22.935 94.365 23.105 94.535 ;
        RECT 22.935 93.905 23.105 94.075 ;
        RECT -282.775 93.245 -282.605 93.415 ;
        RECT -282.315 93.245 -282.145 93.415 ;
        RECT -281.855 93.245 -281.685 93.415 ;
        RECT -281.395 93.245 -281.225 93.415 ;
        RECT -280.935 93.245 -280.765 93.415 ;
        RECT -280.475 93.245 -280.305 93.415 ;
        RECT -280.015 93.245 -279.845 93.415 ;
        RECT -272.855 93.245 -272.685 93.415 ;
        RECT -272.395 93.245 -272.225 93.415 ;
        RECT -271.935 93.245 -271.765 93.415 ;
        RECT -271.475 93.245 -271.305 93.415 ;
        RECT -271.015 93.245 -270.845 93.415 ;
        RECT -270.555 93.245 -270.385 93.415 ;
        RECT -270.095 93.245 -269.925 93.415 ;
        RECT -262.935 93.245 -262.765 93.415 ;
        RECT -262.475 93.245 -262.305 93.415 ;
        RECT -262.015 93.245 -261.845 93.415 ;
        RECT -261.555 93.245 -261.385 93.415 ;
        RECT -261.095 93.245 -260.925 93.415 ;
        RECT -260.635 93.245 -260.465 93.415 ;
        RECT -260.175 93.245 -260.005 93.415 ;
        RECT -253.015 93.245 -252.845 93.415 ;
        RECT -252.555 93.245 -252.385 93.415 ;
        RECT -252.095 93.245 -251.925 93.415 ;
        RECT -251.635 93.245 -251.465 93.415 ;
        RECT -251.175 93.245 -251.005 93.415 ;
        RECT -250.715 93.245 -250.545 93.415 ;
        RECT -250.255 93.245 -250.085 93.415 ;
        RECT -243.095 93.245 -242.925 93.415 ;
        RECT -242.635 93.245 -242.465 93.415 ;
        RECT -242.175 93.245 -242.005 93.415 ;
        RECT -241.715 93.245 -241.545 93.415 ;
        RECT -241.255 93.245 -241.085 93.415 ;
        RECT -240.795 93.245 -240.625 93.415 ;
        RECT -240.335 93.245 -240.165 93.415 ;
        RECT -233.175 93.245 -233.005 93.415 ;
        RECT -232.715 93.245 -232.545 93.415 ;
        RECT -232.255 93.245 -232.085 93.415 ;
        RECT -231.795 93.245 -231.625 93.415 ;
        RECT -231.335 93.245 -231.165 93.415 ;
        RECT -230.875 93.245 -230.705 93.415 ;
        RECT -230.415 93.245 -230.245 93.415 ;
        RECT -223.255 93.245 -223.085 93.415 ;
        RECT -222.795 93.245 -222.625 93.415 ;
        RECT -222.335 93.245 -222.165 93.415 ;
        RECT -221.875 93.245 -221.705 93.415 ;
        RECT -221.415 93.245 -221.245 93.415 ;
        RECT -220.955 93.245 -220.785 93.415 ;
        RECT -220.495 93.245 -220.325 93.415 ;
        RECT -213.335 93.245 -213.165 93.415 ;
        RECT -212.875 93.245 -212.705 93.415 ;
        RECT -212.415 93.245 -212.245 93.415 ;
        RECT -211.955 93.245 -211.785 93.415 ;
        RECT -211.495 93.245 -211.325 93.415 ;
        RECT -211.035 93.245 -210.865 93.415 ;
        RECT -210.575 93.245 -210.405 93.415 ;
        RECT -203.415 93.245 -203.245 93.415 ;
        RECT -202.955 93.245 -202.785 93.415 ;
        RECT -202.495 93.245 -202.325 93.415 ;
        RECT -202.035 93.245 -201.865 93.415 ;
        RECT -201.575 93.245 -201.405 93.415 ;
        RECT -201.115 93.245 -200.945 93.415 ;
        RECT -200.655 93.245 -200.485 93.415 ;
        RECT -193.495 93.245 -193.325 93.415 ;
        RECT -193.035 93.245 -192.865 93.415 ;
        RECT -192.575 93.245 -192.405 93.415 ;
        RECT -192.115 93.245 -191.945 93.415 ;
        RECT -191.655 93.245 -191.485 93.415 ;
        RECT -191.195 93.245 -191.025 93.415 ;
        RECT -190.735 93.245 -190.565 93.415 ;
        RECT -183.575 93.245 -183.405 93.415 ;
        RECT -183.115 93.245 -182.945 93.415 ;
        RECT -182.655 93.245 -182.485 93.415 ;
        RECT -182.195 93.245 -182.025 93.415 ;
        RECT -181.735 93.245 -181.565 93.415 ;
        RECT -181.275 93.245 -181.105 93.415 ;
        RECT -180.815 93.245 -180.645 93.415 ;
        RECT -173.655 93.245 -173.485 93.415 ;
        RECT -173.195 93.245 -173.025 93.415 ;
        RECT -172.735 93.245 -172.565 93.415 ;
        RECT -172.275 93.245 -172.105 93.415 ;
        RECT -171.815 93.245 -171.645 93.415 ;
        RECT -171.355 93.245 -171.185 93.415 ;
        RECT -170.895 93.245 -170.725 93.415 ;
        RECT -163.735 93.245 -163.565 93.415 ;
        RECT -163.275 93.245 -163.105 93.415 ;
        RECT -162.815 93.245 -162.645 93.415 ;
        RECT -162.355 93.245 -162.185 93.415 ;
        RECT -161.895 93.245 -161.725 93.415 ;
        RECT -161.435 93.245 -161.265 93.415 ;
        RECT -160.975 93.245 -160.805 93.415 ;
        RECT -153.815 93.245 -153.645 93.415 ;
        RECT -153.355 93.245 -153.185 93.415 ;
        RECT -152.895 93.245 -152.725 93.415 ;
        RECT -152.435 93.245 -152.265 93.415 ;
        RECT -151.975 93.245 -151.805 93.415 ;
        RECT -151.515 93.245 -151.345 93.415 ;
        RECT -151.055 93.245 -150.885 93.415 ;
        RECT -143.895 93.245 -143.725 93.415 ;
        RECT -143.435 93.245 -143.265 93.415 ;
        RECT -142.975 93.245 -142.805 93.415 ;
        RECT -142.515 93.245 -142.345 93.415 ;
        RECT -142.055 93.245 -141.885 93.415 ;
        RECT -141.595 93.245 -141.425 93.415 ;
        RECT -141.135 93.245 -140.965 93.415 ;
        RECT -133.975 93.245 -133.805 93.415 ;
        RECT -133.515 93.245 -133.345 93.415 ;
        RECT -133.055 93.245 -132.885 93.415 ;
        RECT -132.595 93.245 -132.425 93.415 ;
        RECT -132.135 93.245 -131.965 93.415 ;
        RECT -131.675 93.245 -131.505 93.415 ;
        RECT -131.215 93.245 -131.045 93.415 ;
        RECT -124.055 93.245 -123.885 93.415 ;
        RECT -123.595 93.245 -123.425 93.415 ;
        RECT -123.135 93.245 -122.965 93.415 ;
        RECT -122.675 93.245 -122.505 93.415 ;
        RECT -122.215 93.245 -122.045 93.415 ;
        RECT -121.755 93.245 -121.585 93.415 ;
        RECT -121.295 93.245 -121.125 93.415 ;
        RECT -114.135 93.245 -113.965 93.415 ;
        RECT -113.675 93.245 -113.505 93.415 ;
        RECT -113.215 93.245 -113.045 93.415 ;
        RECT -112.755 93.245 -112.585 93.415 ;
        RECT -112.295 93.245 -112.125 93.415 ;
        RECT -111.835 93.245 -111.665 93.415 ;
        RECT -111.375 93.245 -111.205 93.415 ;
        RECT -104.215 93.245 -104.045 93.415 ;
        RECT -103.755 93.245 -103.585 93.415 ;
        RECT -103.295 93.245 -103.125 93.415 ;
        RECT -102.835 93.245 -102.665 93.415 ;
        RECT -102.375 93.245 -102.205 93.415 ;
        RECT -101.915 93.245 -101.745 93.415 ;
        RECT -101.455 93.245 -101.285 93.415 ;
        RECT -94.295 93.245 -94.125 93.415 ;
        RECT -93.835 93.245 -93.665 93.415 ;
        RECT -93.375 93.245 -93.205 93.415 ;
        RECT -92.915 93.245 -92.745 93.415 ;
        RECT -92.455 93.245 -92.285 93.415 ;
        RECT -91.995 93.245 -91.825 93.415 ;
        RECT -91.535 93.245 -91.365 93.415 ;
        RECT -84.375 93.245 -84.205 93.415 ;
        RECT -83.915 93.245 -83.745 93.415 ;
        RECT -83.455 93.245 -83.285 93.415 ;
        RECT -82.995 93.245 -82.825 93.415 ;
        RECT -82.535 93.245 -82.365 93.415 ;
        RECT -82.075 93.245 -81.905 93.415 ;
        RECT -81.615 93.245 -81.445 93.415 ;
        RECT -74.455 93.245 -74.285 93.415 ;
        RECT -73.995 93.245 -73.825 93.415 ;
        RECT -73.535 93.245 -73.365 93.415 ;
        RECT -73.075 93.245 -72.905 93.415 ;
        RECT -72.615 93.245 -72.445 93.415 ;
        RECT -72.155 93.245 -71.985 93.415 ;
        RECT -71.695 93.245 -71.525 93.415 ;
        RECT -64.535 93.245 -64.365 93.415 ;
        RECT -64.075 93.245 -63.905 93.415 ;
        RECT -63.615 93.245 -63.445 93.415 ;
        RECT -63.155 93.245 -62.985 93.415 ;
        RECT -62.695 93.245 -62.525 93.415 ;
        RECT -62.235 93.245 -62.065 93.415 ;
        RECT -61.775 93.245 -61.605 93.415 ;
        RECT -54.615 93.245 -54.445 93.415 ;
        RECT -54.155 93.245 -53.985 93.415 ;
        RECT -53.695 93.245 -53.525 93.415 ;
        RECT -53.235 93.245 -53.065 93.415 ;
        RECT -52.775 93.245 -52.605 93.415 ;
        RECT -52.315 93.245 -52.145 93.415 ;
        RECT -51.855 93.245 -51.685 93.415 ;
        RECT -44.695 93.245 -44.525 93.415 ;
        RECT -44.235 93.245 -44.065 93.415 ;
        RECT -43.775 93.245 -43.605 93.415 ;
        RECT -43.315 93.245 -43.145 93.415 ;
        RECT -42.855 93.245 -42.685 93.415 ;
        RECT -42.395 93.245 -42.225 93.415 ;
        RECT -41.935 93.245 -41.765 93.415 ;
        RECT -34.775 93.245 -34.605 93.415 ;
        RECT -34.315 93.245 -34.145 93.415 ;
        RECT -33.855 93.245 -33.685 93.415 ;
        RECT -33.395 93.245 -33.225 93.415 ;
        RECT -32.935 93.245 -32.765 93.415 ;
        RECT -32.475 93.245 -32.305 93.415 ;
        RECT -32.015 93.245 -31.845 93.415 ;
        RECT -24.855 93.245 -24.685 93.415 ;
        RECT -24.395 93.245 -24.225 93.415 ;
        RECT -23.935 93.245 -23.765 93.415 ;
        RECT -23.475 93.245 -23.305 93.415 ;
        RECT -23.015 93.245 -22.845 93.415 ;
        RECT -22.555 93.245 -22.385 93.415 ;
        RECT -22.095 93.245 -21.925 93.415 ;
        RECT -14.935 93.245 -14.765 93.415 ;
        RECT -14.475 93.245 -14.305 93.415 ;
        RECT -14.015 93.245 -13.845 93.415 ;
        RECT -13.555 93.245 -13.385 93.415 ;
        RECT -13.095 93.245 -12.925 93.415 ;
        RECT -12.635 93.245 -12.465 93.415 ;
        RECT -12.175 93.245 -12.005 93.415 ;
        RECT -5.015 93.245 -4.845 93.415 ;
        RECT -4.555 93.245 -4.385 93.415 ;
        RECT -4.095 93.245 -3.925 93.415 ;
        RECT -3.635 93.245 -3.465 93.415 ;
        RECT -3.175 93.245 -3.005 93.415 ;
        RECT -2.715 93.245 -2.545 93.415 ;
        RECT -2.255 93.245 -2.085 93.415 ;
        RECT 4.905 93.245 5.075 93.415 ;
        RECT 5.365 93.245 5.535 93.415 ;
        RECT 5.825 93.245 5.995 93.415 ;
        RECT 6.285 93.245 6.455 93.415 ;
        RECT 6.745 93.245 6.915 93.415 ;
        RECT 7.205 93.245 7.375 93.415 ;
        RECT 7.665 93.245 7.835 93.415 ;
        RECT 14.825 93.245 14.995 93.415 ;
        RECT 15.285 93.245 15.455 93.415 ;
        RECT 15.745 93.245 15.915 93.415 ;
        RECT 16.205 93.245 16.375 93.415 ;
        RECT 16.665 93.245 16.835 93.415 ;
        RECT 17.125 93.245 17.295 93.415 ;
        RECT 17.585 93.245 17.755 93.415 ;
        RECT -287.735 90.525 -287.565 90.695 ;
        RECT -287.275 90.525 -287.105 90.695 ;
        RECT -286.815 90.525 -286.645 90.695 ;
        RECT -286.355 90.525 -286.185 90.695 ;
        RECT -285.895 90.525 -285.725 90.695 ;
        RECT -285.435 90.525 -285.265 90.695 ;
        RECT -284.975 90.525 -284.805 90.695 ;
        RECT -277.815 90.525 -277.645 90.695 ;
        RECT -277.355 90.525 -277.185 90.695 ;
        RECT -276.895 90.525 -276.725 90.695 ;
        RECT -276.435 90.525 -276.265 90.695 ;
        RECT -275.975 90.525 -275.805 90.695 ;
        RECT -275.515 90.525 -275.345 90.695 ;
        RECT -275.055 90.525 -274.885 90.695 ;
        RECT -267.895 90.525 -267.725 90.695 ;
        RECT -267.435 90.525 -267.265 90.695 ;
        RECT -266.975 90.525 -266.805 90.695 ;
        RECT -266.515 90.525 -266.345 90.695 ;
        RECT -266.055 90.525 -265.885 90.695 ;
        RECT -265.595 90.525 -265.425 90.695 ;
        RECT -265.135 90.525 -264.965 90.695 ;
        RECT -257.975 90.525 -257.805 90.695 ;
        RECT -257.515 90.525 -257.345 90.695 ;
        RECT -257.055 90.525 -256.885 90.695 ;
        RECT -256.595 90.525 -256.425 90.695 ;
        RECT -256.135 90.525 -255.965 90.695 ;
        RECT -255.675 90.525 -255.505 90.695 ;
        RECT -255.215 90.525 -255.045 90.695 ;
        RECT -248.055 90.525 -247.885 90.695 ;
        RECT -247.595 90.525 -247.425 90.695 ;
        RECT -247.135 90.525 -246.965 90.695 ;
        RECT -246.675 90.525 -246.505 90.695 ;
        RECT -246.215 90.525 -246.045 90.695 ;
        RECT -245.755 90.525 -245.585 90.695 ;
        RECT -245.295 90.525 -245.125 90.695 ;
        RECT -238.135 90.525 -237.965 90.695 ;
        RECT -237.675 90.525 -237.505 90.695 ;
        RECT -237.215 90.525 -237.045 90.695 ;
        RECT -236.755 90.525 -236.585 90.695 ;
        RECT -236.295 90.525 -236.125 90.695 ;
        RECT -235.835 90.525 -235.665 90.695 ;
        RECT -235.375 90.525 -235.205 90.695 ;
        RECT -228.215 90.525 -228.045 90.695 ;
        RECT -227.755 90.525 -227.585 90.695 ;
        RECT -227.295 90.525 -227.125 90.695 ;
        RECT -226.835 90.525 -226.665 90.695 ;
        RECT -226.375 90.525 -226.205 90.695 ;
        RECT -225.915 90.525 -225.745 90.695 ;
        RECT -225.455 90.525 -225.285 90.695 ;
        RECT -218.295 90.525 -218.125 90.695 ;
        RECT -217.835 90.525 -217.665 90.695 ;
        RECT -217.375 90.525 -217.205 90.695 ;
        RECT -216.915 90.525 -216.745 90.695 ;
        RECT -216.455 90.525 -216.285 90.695 ;
        RECT -215.995 90.525 -215.825 90.695 ;
        RECT -215.535 90.525 -215.365 90.695 ;
        RECT -208.375 90.525 -208.205 90.695 ;
        RECT -207.915 90.525 -207.745 90.695 ;
        RECT -207.455 90.525 -207.285 90.695 ;
        RECT -206.995 90.525 -206.825 90.695 ;
        RECT -206.535 90.525 -206.365 90.695 ;
        RECT -206.075 90.525 -205.905 90.695 ;
        RECT -205.615 90.525 -205.445 90.695 ;
        RECT -198.455 90.525 -198.285 90.695 ;
        RECT -197.995 90.525 -197.825 90.695 ;
        RECT -197.535 90.525 -197.365 90.695 ;
        RECT -197.075 90.525 -196.905 90.695 ;
        RECT -196.615 90.525 -196.445 90.695 ;
        RECT -196.155 90.525 -195.985 90.695 ;
        RECT -195.695 90.525 -195.525 90.695 ;
        RECT -188.535 90.525 -188.365 90.695 ;
        RECT -188.075 90.525 -187.905 90.695 ;
        RECT -187.615 90.525 -187.445 90.695 ;
        RECT -187.155 90.525 -186.985 90.695 ;
        RECT -186.695 90.525 -186.525 90.695 ;
        RECT -186.235 90.525 -186.065 90.695 ;
        RECT -185.775 90.525 -185.605 90.695 ;
        RECT -178.615 90.525 -178.445 90.695 ;
        RECT -178.155 90.525 -177.985 90.695 ;
        RECT -177.695 90.525 -177.525 90.695 ;
        RECT -177.235 90.525 -177.065 90.695 ;
        RECT -176.775 90.525 -176.605 90.695 ;
        RECT -176.315 90.525 -176.145 90.695 ;
        RECT -175.855 90.525 -175.685 90.695 ;
        RECT -168.695 90.525 -168.525 90.695 ;
        RECT -168.235 90.525 -168.065 90.695 ;
        RECT -167.775 90.525 -167.605 90.695 ;
        RECT -167.315 90.525 -167.145 90.695 ;
        RECT -166.855 90.525 -166.685 90.695 ;
        RECT -166.395 90.525 -166.225 90.695 ;
        RECT -165.935 90.525 -165.765 90.695 ;
        RECT -158.775 90.525 -158.605 90.695 ;
        RECT -158.315 90.525 -158.145 90.695 ;
        RECT -157.855 90.525 -157.685 90.695 ;
        RECT -157.395 90.525 -157.225 90.695 ;
        RECT -156.935 90.525 -156.765 90.695 ;
        RECT -156.475 90.525 -156.305 90.695 ;
        RECT -156.015 90.525 -155.845 90.695 ;
        RECT -148.855 90.525 -148.685 90.695 ;
        RECT -148.395 90.525 -148.225 90.695 ;
        RECT -147.935 90.525 -147.765 90.695 ;
        RECT -147.475 90.525 -147.305 90.695 ;
        RECT -147.015 90.525 -146.845 90.695 ;
        RECT -146.555 90.525 -146.385 90.695 ;
        RECT -146.095 90.525 -145.925 90.695 ;
        RECT -138.935 90.525 -138.765 90.695 ;
        RECT -138.475 90.525 -138.305 90.695 ;
        RECT -138.015 90.525 -137.845 90.695 ;
        RECT -137.555 90.525 -137.385 90.695 ;
        RECT -137.095 90.525 -136.925 90.695 ;
        RECT -136.635 90.525 -136.465 90.695 ;
        RECT -136.175 90.525 -136.005 90.695 ;
        RECT -129.015 90.525 -128.845 90.695 ;
        RECT -128.555 90.525 -128.385 90.695 ;
        RECT -128.095 90.525 -127.925 90.695 ;
        RECT -127.635 90.525 -127.465 90.695 ;
        RECT -127.175 90.525 -127.005 90.695 ;
        RECT -126.715 90.525 -126.545 90.695 ;
        RECT -126.255 90.525 -126.085 90.695 ;
        RECT -119.095 90.525 -118.925 90.695 ;
        RECT -118.635 90.525 -118.465 90.695 ;
        RECT -118.175 90.525 -118.005 90.695 ;
        RECT -117.715 90.525 -117.545 90.695 ;
        RECT -117.255 90.525 -117.085 90.695 ;
        RECT -116.795 90.525 -116.625 90.695 ;
        RECT -116.335 90.525 -116.165 90.695 ;
        RECT -109.175 90.525 -109.005 90.695 ;
        RECT -108.715 90.525 -108.545 90.695 ;
        RECT -108.255 90.525 -108.085 90.695 ;
        RECT -107.795 90.525 -107.625 90.695 ;
        RECT -107.335 90.525 -107.165 90.695 ;
        RECT -106.875 90.525 -106.705 90.695 ;
        RECT -106.415 90.525 -106.245 90.695 ;
        RECT -99.255 90.525 -99.085 90.695 ;
        RECT -98.795 90.525 -98.625 90.695 ;
        RECT -98.335 90.525 -98.165 90.695 ;
        RECT -97.875 90.525 -97.705 90.695 ;
        RECT -97.415 90.525 -97.245 90.695 ;
        RECT -96.955 90.525 -96.785 90.695 ;
        RECT -96.495 90.525 -96.325 90.695 ;
        RECT -89.335 90.525 -89.165 90.695 ;
        RECT -88.875 90.525 -88.705 90.695 ;
        RECT -88.415 90.525 -88.245 90.695 ;
        RECT -87.955 90.525 -87.785 90.695 ;
        RECT -87.495 90.525 -87.325 90.695 ;
        RECT -87.035 90.525 -86.865 90.695 ;
        RECT -86.575 90.525 -86.405 90.695 ;
        RECT -79.415 90.525 -79.245 90.695 ;
        RECT -78.955 90.525 -78.785 90.695 ;
        RECT -78.495 90.525 -78.325 90.695 ;
        RECT -78.035 90.525 -77.865 90.695 ;
        RECT -77.575 90.525 -77.405 90.695 ;
        RECT -77.115 90.525 -76.945 90.695 ;
        RECT -76.655 90.525 -76.485 90.695 ;
        RECT -69.495 90.525 -69.325 90.695 ;
        RECT -69.035 90.525 -68.865 90.695 ;
        RECT -68.575 90.525 -68.405 90.695 ;
        RECT -68.115 90.525 -67.945 90.695 ;
        RECT -67.655 90.525 -67.485 90.695 ;
        RECT -67.195 90.525 -67.025 90.695 ;
        RECT -66.735 90.525 -66.565 90.695 ;
        RECT -59.575 90.525 -59.405 90.695 ;
        RECT -59.115 90.525 -58.945 90.695 ;
        RECT -58.655 90.525 -58.485 90.695 ;
        RECT -58.195 90.525 -58.025 90.695 ;
        RECT -57.735 90.525 -57.565 90.695 ;
        RECT -57.275 90.525 -57.105 90.695 ;
        RECT -56.815 90.525 -56.645 90.695 ;
        RECT -49.655 90.525 -49.485 90.695 ;
        RECT -49.195 90.525 -49.025 90.695 ;
        RECT -48.735 90.525 -48.565 90.695 ;
        RECT -48.275 90.525 -48.105 90.695 ;
        RECT -47.815 90.525 -47.645 90.695 ;
        RECT -47.355 90.525 -47.185 90.695 ;
        RECT -46.895 90.525 -46.725 90.695 ;
        RECT -39.735 90.525 -39.565 90.695 ;
        RECT -39.275 90.525 -39.105 90.695 ;
        RECT -38.815 90.525 -38.645 90.695 ;
        RECT -38.355 90.525 -38.185 90.695 ;
        RECT -37.895 90.525 -37.725 90.695 ;
        RECT -37.435 90.525 -37.265 90.695 ;
        RECT -36.975 90.525 -36.805 90.695 ;
        RECT -29.815 90.525 -29.645 90.695 ;
        RECT -29.355 90.525 -29.185 90.695 ;
        RECT -28.895 90.525 -28.725 90.695 ;
        RECT -28.435 90.525 -28.265 90.695 ;
        RECT -27.975 90.525 -27.805 90.695 ;
        RECT -27.515 90.525 -27.345 90.695 ;
        RECT -27.055 90.525 -26.885 90.695 ;
        RECT -19.895 90.525 -19.725 90.695 ;
        RECT -19.435 90.525 -19.265 90.695 ;
        RECT -18.975 90.525 -18.805 90.695 ;
        RECT -18.515 90.525 -18.345 90.695 ;
        RECT -18.055 90.525 -17.885 90.695 ;
        RECT -17.595 90.525 -17.425 90.695 ;
        RECT -17.135 90.525 -16.965 90.695 ;
        RECT -9.975 90.525 -9.805 90.695 ;
        RECT -9.515 90.525 -9.345 90.695 ;
        RECT -9.055 90.525 -8.885 90.695 ;
        RECT -8.595 90.525 -8.425 90.695 ;
        RECT -8.135 90.525 -7.965 90.695 ;
        RECT -7.675 90.525 -7.505 90.695 ;
        RECT -7.215 90.525 -7.045 90.695 ;
        RECT -0.055 90.525 0.115 90.695 ;
        RECT 0.405 90.525 0.575 90.695 ;
        RECT 0.865 90.525 1.035 90.695 ;
        RECT 1.325 90.525 1.495 90.695 ;
        RECT 1.785 90.525 1.955 90.695 ;
        RECT 2.245 90.525 2.415 90.695 ;
        RECT 2.705 90.525 2.875 90.695 ;
        RECT 9.865 90.525 10.035 90.695 ;
        RECT 10.325 90.525 10.495 90.695 ;
        RECT 10.785 90.525 10.955 90.695 ;
        RECT 11.245 90.525 11.415 90.695 ;
        RECT 11.705 90.525 11.875 90.695 ;
        RECT 12.165 90.525 12.335 90.695 ;
        RECT 12.625 90.525 12.795 90.695 ;
        RECT 19.785 90.525 19.955 90.695 ;
        RECT 20.245 90.525 20.415 90.695 ;
        RECT 20.705 90.525 20.875 90.695 ;
        RECT 21.165 90.525 21.335 90.695 ;
        RECT 21.625 90.525 21.795 90.695 ;
        RECT 22.085 90.525 22.255 90.695 ;
        RECT 22.545 90.525 22.715 90.695 ;
        RECT -283.165 89.865 -282.995 90.035 ;
        RECT -283.165 89.405 -282.995 89.575 ;
        RECT -279.625 89.865 -279.455 90.035 ;
        RECT -273.245 89.865 -273.075 90.035 ;
        RECT -279.625 89.405 -279.455 89.575 ;
        RECT -273.245 89.405 -273.075 89.575 ;
        RECT -281.395 89.135 -281.225 89.305 ;
        RECT -283.165 88.945 -282.995 89.115 ;
        RECT -279.625 88.945 -279.455 89.115 ;
        RECT -269.705 89.865 -269.535 90.035 ;
        RECT -263.325 89.865 -263.155 90.035 ;
        RECT -269.705 89.405 -269.535 89.575 ;
        RECT -263.325 89.405 -263.155 89.575 ;
        RECT -271.475 89.135 -271.305 89.305 ;
        RECT -273.245 88.945 -273.075 89.115 ;
        RECT -269.705 88.945 -269.535 89.115 ;
        RECT -259.785 89.865 -259.615 90.035 ;
        RECT -253.405 89.865 -253.235 90.035 ;
        RECT -259.785 89.405 -259.615 89.575 ;
        RECT -253.405 89.405 -253.235 89.575 ;
        RECT -261.555 89.135 -261.385 89.305 ;
        RECT -263.325 88.945 -263.155 89.115 ;
        RECT -259.785 88.945 -259.615 89.115 ;
        RECT -249.865 89.865 -249.695 90.035 ;
        RECT -243.485 89.865 -243.315 90.035 ;
        RECT -249.865 89.405 -249.695 89.575 ;
        RECT -243.485 89.405 -243.315 89.575 ;
        RECT -251.635 89.135 -251.465 89.305 ;
        RECT -253.405 88.945 -253.235 89.115 ;
        RECT -249.865 88.945 -249.695 89.115 ;
        RECT -239.945 89.865 -239.775 90.035 ;
        RECT -233.565 89.865 -233.395 90.035 ;
        RECT -239.945 89.405 -239.775 89.575 ;
        RECT -233.565 89.405 -233.395 89.575 ;
        RECT -241.715 89.135 -241.545 89.305 ;
        RECT -243.485 88.945 -243.315 89.115 ;
        RECT -239.945 88.945 -239.775 89.115 ;
        RECT -230.025 89.865 -229.855 90.035 ;
        RECT -223.645 89.865 -223.475 90.035 ;
        RECT -230.025 89.405 -229.855 89.575 ;
        RECT -223.645 89.405 -223.475 89.575 ;
        RECT -231.795 89.135 -231.625 89.305 ;
        RECT -233.565 88.945 -233.395 89.115 ;
        RECT -230.025 88.945 -229.855 89.115 ;
        RECT -220.105 89.865 -219.935 90.035 ;
        RECT -213.725 89.865 -213.555 90.035 ;
        RECT -220.105 89.405 -219.935 89.575 ;
        RECT -213.725 89.405 -213.555 89.575 ;
        RECT -221.875 89.135 -221.705 89.305 ;
        RECT -223.645 88.945 -223.475 89.115 ;
        RECT -220.105 88.945 -219.935 89.115 ;
        RECT -210.185 89.865 -210.015 90.035 ;
        RECT -203.805 89.865 -203.635 90.035 ;
        RECT -210.185 89.405 -210.015 89.575 ;
        RECT -203.805 89.405 -203.635 89.575 ;
        RECT -211.955 89.135 -211.785 89.305 ;
        RECT -213.725 88.945 -213.555 89.115 ;
        RECT -210.185 88.945 -210.015 89.115 ;
        RECT -200.265 89.865 -200.095 90.035 ;
        RECT -193.885 89.865 -193.715 90.035 ;
        RECT -200.265 89.405 -200.095 89.575 ;
        RECT -193.885 89.405 -193.715 89.575 ;
        RECT -202.035 89.135 -201.865 89.305 ;
        RECT -203.805 88.945 -203.635 89.115 ;
        RECT -200.265 88.945 -200.095 89.115 ;
        RECT -190.345 89.865 -190.175 90.035 ;
        RECT -183.965 89.865 -183.795 90.035 ;
        RECT -190.345 89.405 -190.175 89.575 ;
        RECT -183.965 89.405 -183.795 89.575 ;
        RECT -192.115 89.135 -191.945 89.305 ;
        RECT -193.885 88.945 -193.715 89.115 ;
        RECT -190.345 88.945 -190.175 89.115 ;
        RECT -180.425 89.865 -180.255 90.035 ;
        RECT -174.045 89.865 -173.875 90.035 ;
        RECT -180.425 89.405 -180.255 89.575 ;
        RECT -174.045 89.405 -173.875 89.575 ;
        RECT -182.195 89.135 -182.025 89.305 ;
        RECT -183.965 88.945 -183.795 89.115 ;
        RECT -180.425 88.945 -180.255 89.115 ;
        RECT -170.505 89.865 -170.335 90.035 ;
        RECT -164.125 89.865 -163.955 90.035 ;
        RECT -170.505 89.405 -170.335 89.575 ;
        RECT -164.125 89.405 -163.955 89.575 ;
        RECT -172.275 89.135 -172.105 89.305 ;
        RECT -174.045 88.945 -173.875 89.115 ;
        RECT -170.505 88.945 -170.335 89.115 ;
        RECT -160.585 89.865 -160.415 90.035 ;
        RECT -154.205 89.865 -154.035 90.035 ;
        RECT -160.585 89.405 -160.415 89.575 ;
        RECT -154.205 89.405 -154.035 89.575 ;
        RECT -162.355 89.135 -162.185 89.305 ;
        RECT -164.125 88.945 -163.955 89.115 ;
        RECT -160.585 88.945 -160.415 89.115 ;
        RECT -150.665 89.865 -150.495 90.035 ;
        RECT -144.285 89.865 -144.115 90.035 ;
        RECT -150.665 89.405 -150.495 89.575 ;
        RECT -144.285 89.405 -144.115 89.575 ;
        RECT -152.435 89.135 -152.265 89.305 ;
        RECT -154.205 88.945 -154.035 89.115 ;
        RECT -150.665 88.945 -150.495 89.115 ;
        RECT -140.745 89.865 -140.575 90.035 ;
        RECT -134.365 89.865 -134.195 90.035 ;
        RECT -140.745 89.405 -140.575 89.575 ;
        RECT -134.365 89.405 -134.195 89.575 ;
        RECT -142.515 89.135 -142.345 89.305 ;
        RECT -144.285 88.945 -144.115 89.115 ;
        RECT -140.745 88.945 -140.575 89.115 ;
        RECT -130.825 89.865 -130.655 90.035 ;
        RECT -124.445 89.865 -124.275 90.035 ;
        RECT -130.825 89.405 -130.655 89.575 ;
        RECT -124.445 89.405 -124.275 89.575 ;
        RECT -132.595 89.135 -132.425 89.305 ;
        RECT -134.365 88.945 -134.195 89.115 ;
        RECT -130.825 88.945 -130.655 89.115 ;
        RECT -120.905 89.865 -120.735 90.035 ;
        RECT -114.525 89.865 -114.355 90.035 ;
        RECT -120.905 89.405 -120.735 89.575 ;
        RECT -114.525 89.405 -114.355 89.575 ;
        RECT -122.675 89.135 -122.505 89.305 ;
        RECT -124.445 88.945 -124.275 89.115 ;
        RECT -120.905 88.945 -120.735 89.115 ;
        RECT -110.985 89.865 -110.815 90.035 ;
        RECT -104.605 89.865 -104.435 90.035 ;
        RECT -110.985 89.405 -110.815 89.575 ;
        RECT -104.605 89.405 -104.435 89.575 ;
        RECT -112.755 89.135 -112.585 89.305 ;
        RECT -114.525 88.945 -114.355 89.115 ;
        RECT -110.985 88.945 -110.815 89.115 ;
        RECT -101.065 89.865 -100.895 90.035 ;
        RECT -94.685 89.865 -94.515 90.035 ;
        RECT -101.065 89.405 -100.895 89.575 ;
        RECT -94.685 89.405 -94.515 89.575 ;
        RECT -102.835 89.135 -102.665 89.305 ;
        RECT -104.605 88.945 -104.435 89.115 ;
        RECT -101.065 88.945 -100.895 89.115 ;
        RECT -91.145 89.865 -90.975 90.035 ;
        RECT -84.765 89.865 -84.595 90.035 ;
        RECT -91.145 89.405 -90.975 89.575 ;
        RECT -84.765 89.405 -84.595 89.575 ;
        RECT -92.915 89.135 -92.745 89.305 ;
        RECT -94.685 88.945 -94.515 89.115 ;
        RECT -91.145 88.945 -90.975 89.115 ;
        RECT -81.225 89.865 -81.055 90.035 ;
        RECT -74.845 89.865 -74.675 90.035 ;
        RECT -81.225 89.405 -81.055 89.575 ;
        RECT -74.845 89.405 -74.675 89.575 ;
        RECT -82.995 89.135 -82.825 89.305 ;
        RECT -84.765 88.945 -84.595 89.115 ;
        RECT -81.225 88.945 -81.055 89.115 ;
        RECT -71.305 89.865 -71.135 90.035 ;
        RECT -64.925 89.865 -64.755 90.035 ;
        RECT -71.305 89.405 -71.135 89.575 ;
        RECT -64.925 89.405 -64.755 89.575 ;
        RECT -73.075 89.135 -72.905 89.305 ;
        RECT -74.845 88.945 -74.675 89.115 ;
        RECT -71.305 88.945 -71.135 89.115 ;
        RECT -61.385 89.865 -61.215 90.035 ;
        RECT -55.005 89.865 -54.835 90.035 ;
        RECT -61.385 89.405 -61.215 89.575 ;
        RECT -55.005 89.405 -54.835 89.575 ;
        RECT -63.155 89.135 -62.985 89.305 ;
        RECT -64.925 88.945 -64.755 89.115 ;
        RECT -61.385 88.945 -61.215 89.115 ;
        RECT -51.465 89.865 -51.295 90.035 ;
        RECT -45.085 89.865 -44.915 90.035 ;
        RECT -51.465 89.405 -51.295 89.575 ;
        RECT -45.085 89.405 -44.915 89.575 ;
        RECT -53.235 89.135 -53.065 89.305 ;
        RECT -55.005 88.945 -54.835 89.115 ;
        RECT -51.465 88.945 -51.295 89.115 ;
        RECT -41.545 89.865 -41.375 90.035 ;
        RECT -35.165 89.865 -34.995 90.035 ;
        RECT -41.545 89.405 -41.375 89.575 ;
        RECT -35.165 89.405 -34.995 89.575 ;
        RECT -43.315 89.135 -43.145 89.305 ;
        RECT -45.085 88.945 -44.915 89.115 ;
        RECT -41.545 88.945 -41.375 89.115 ;
        RECT -31.625 89.865 -31.455 90.035 ;
        RECT -25.245 89.865 -25.075 90.035 ;
        RECT -31.625 89.405 -31.455 89.575 ;
        RECT -25.245 89.405 -25.075 89.575 ;
        RECT -33.395 89.135 -33.225 89.305 ;
        RECT -35.165 88.945 -34.995 89.115 ;
        RECT -31.625 88.945 -31.455 89.115 ;
        RECT -21.705 89.865 -21.535 90.035 ;
        RECT -15.325 89.865 -15.155 90.035 ;
        RECT -21.705 89.405 -21.535 89.575 ;
        RECT -15.325 89.405 -15.155 89.575 ;
        RECT -23.475 89.135 -23.305 89.305 ;
        RECT -25.245 88.945 -25.075 89.115 ;
        RECT -21.705 88.945 -21.535 89.115 ;
        RECT -11.785 89.865 -11.615 90.035 ;
        RECT -5.405 89.865 -5.235 90.035 ;
        RECT -11.785 89.405 -11.615 89.575 ;
        RECT -5.405 89.405 -5.235 89.575 ;
        RECT -13.555 89.135 -13.385 89.305 ;
        RECT -15.325 88.945 -15.155 89.115 ;
        RECT -11.785 88.945 -11.615 89.115 ;
        RECT -1.865 89.865 -1.695 90.035 ;
        RECT 4.515 89.865 4.685 90.035 ;
        RECT -1.865 89.405 -1.695 89.575 ;
        RECT 4.515 89.405 4.685 89.575 ;
        RECT -3.635 89.135 -3.465 89.305 ;
        RECT -5.405 88.945 -5.235 89.115 ;
        RECT -1.865 88.945 -1.695 89.115 ;
        RECT 8.055 89.865 8.225 90.035 ;
        RECT 14.435 89.865 14.605 90.035 ;
        RECT 8.055 89.405 8.225 89.575 ;
        RECT 14.435 89.405 14.605 89.575 ;
        RECT 6.285 89.135 6.455 89.305 ;
        RECT 4.515 88.945 4.685 89.115 ;
        RECT 8.055 88.945 8.225 89.115 ;
        RECT 17.975 89.865 18.145 90.035 ;
        RECT 17.975 89.405 18.145 89.575 ;
        RECT 16.205 89.135 16.375 89.305 ;
        RECT 14.435 88.945 14.605 89.115 ;
        RECT 17.975 88.945 18.145 89.115 ;
      LAYER met1 ;
        RECT -288.280 93.760 -284.260 95.140 ;
        RECT -278.360 93.760 -274.340 95.140 ;
        RECT -268.440 93.760 -264.420 95.140 ;
        RECT -258.520 93.760 -254.500 95.140 ;
        RECT -248.600 93.760 -244.580 95.140 ;
        RECT -238.680 93.760 -234.660 95.140 ;
        RECT -228.760 93.760 -224.740 95.140 ;
        RECT -218.840 93.760 -214.820 95.140 ;
        RECT -208.920 93.760 -204.900 95.140 ;
        RECT -199.000 93.760 -194.980 95.140 ;
        RECT -189.080 93.760 -185.060 95.140 ;
        RECT -179.160 93.760 -175.140 95.140 ;
        RECT -169.240 93.760 -165.220 95.140 ;
        RECT -159.320 93.760 -155.300 95.140 ;
        RECT -149.400 93.760 -145.380 95.140 ;
        RECT -139.480 93.760 -135.460 95.140 ;
        RECT -129.560 93.760 -125.540 95.140 ;
        RECT -119.640 93.760 -115.620 95.140 ;
        RECT -109.720 93.760 -105.700 95.140 ;
        RECT -99.800 93.760 -95.780 95.140 ;
        RECT -89.880 93.760 -85.860 95.140 ;
        RECT -79.960 93.760 -75.940 95.140 ;
        RECT -70.040 93.760 -66.020 95.140 ;
        RECT -60.120 93.760 -56.100 95.140 ;
        RECT -50.200 93.760 -46.180 95.140 ;
        RECT -40.280 93.760 -36.260 95.140 ;
        RECT -30.360 93.760 -26.340 95.140 ;
        RECT -20.440 93.760 -16.420 95.140 ;
        RECT -10.520 93.760 -6.500 95.140 ;
        RECT -0.600 93.760 3.420 95.140 ;
        RECT 9.320 93.760 13.340 95.140 ;
        RECT 19.240 93.760 23.260 95.140 ;
        RECT -282.920 93.090 -279.700 93.570 ;
        RECT -273.000 93.090 -269.780 93.570 ;
        RECT -263.080 93.090 -259.860 93.570 ;
        RECT -253.160 93.090 -249.940 93.570 ;
        RECT -243.240 93.090 -240.020 93.570 ;
        RECT -233.320 93.090 -230.100 93.570 ;
        RECT -223.400 93.090 -220.180 93.570 ;
        RECT -213.480 93.090 -210.260 93.570 ;
        RECT -203.560 93.090 -200.340 93.570 ;
        RECT -193.640 93.090 -190.420 93.570 ;
        RECT -183.720 93.090 -180.500 93.570 ;
        RECT -173.800 93.090 -170.580 93.570 ;
        RECT -163.880 93.090 -160.660 93.570 ;
        RECT -153.960 93.090 -150.740 93.570 ;
        RECT -144.040 93.090 -140.820 93.570 ;
        RECT -134.120 93.090 -130.900 93.570 ;
        RECT -124.200 93.090 -120.980 93.570 ;
        RECT -114.280 93.090 -111.060 93.570 ;
        RECT -104.360 93.090 -101.140 93.570 ;
        RECT -94.440 93.090 -91.220 93.570 ;
        RECT -84.520 93.090 -81.300 93.570 ;
        RECT -74.600 93.090 -71.380 93.570 ;
        RECT -64.680 93.090 -61.460 93.570 ;
        RECT -54.760 93.090 -51.540 93.570 ;
        RECT -44.840 93.090 -41.620 93.570 ;
        RECT -34.920 93.090 -31.700 93.570 ;
        RECT -25.000 93.090 -21.780 93.570 ;
        RECT -15.080 93.090 -11.860 93.570 ;
        RECT -5.160 93.090 -1.940 93.570 ;
        RECT 4.760 93.090 7.980 93.570 ;
        RECT 14.680 93.090 17.900 93.570 ;
        RECT -287.880 90.370 -284.660 90.850 ;
        RECT -277.960 90.370 -274.740 90.850 ;
        RECT -268.040 90.370 -264.820 90.850 ;
        RECT -258.120 90.370 -254.900 90.850 ;
        RECT -248.200 90.370 -244.980 90.850 ;
        RECT -238.280 90.370 -235.060 90.850 ;
        RECT -228.360 90.370 -225.140 90.850 ;
        RECT -218.440 90.370 -215.220 90.850 ;
        RECT -208.520 90.370 -205.300 90.850 ;
        RECT -198.600 90.370 -195.380 90.850 ;
        RECT -188.680 90.370 -185.460 90.850 ;
        RECT -178.760 90.370 -175.540 90.850 ;
        RECT -168.840 90.370 -165.620 90.850 ;
        RECT -158.920 90.370 -155.700 90.850 ;
        RECT -149.000 90.370 -145.780 90.850 ;
        RECT -139.080 90.370 -135.860 90.850 ;
        RECT -129.160 90.370 -125.940 90.850 ;
        RECT -119.240 90.370 -116.020 90.850 ;
        RECT -109.320 90.370 -106.100 90.850 ;
        RECT -99.400 90.370 -96.180 90.850 ;
        RECT -89.480 90.370 -86.260 90.850 ;
        RECT -79.560 90.370 -76.340 90.850 ;
        RECT -69.640 90.370 -66.420 90.850 ;
        RECT -59.720 90.370 -56.500 90.850 ;
        RECT -49.800 90.370 -46.580 90.850 ;
        RECT -39.880 90.370 -36.660 90.850 ;
        RECT -29.960 90.370 -26.740 90.850 ;
        RECT -20.040 90.370 -16.820 90.850 ;
        RECT -10.120 90.370 -6.900 90.850 ;
        RECT -0.200 90.370 3.020 90.850 ;
        RECT 9.720 90.370 12.940 90.850 ;
        RECT 19.640 90.370 22.860 90.850 ;
        RECT -283.320 88.800 -279.300 90.180 ;
        RECT -273.400 88.800 -269.380 90.180 ;
        RECT -263.480 88.800 -259.460 90.180 ;
        RECT -253.560 88.800 -249.540 90.180 ;
        RECT -243.640 88.800 -239.620 90.180 ;
        RECT -233.720 88.800 -229.700 90.180 ;
        RECT -223.800 88.800 -219.780 90.180 ;
        RECT -213.880 88.800 -209.860 90.180 ;
        RECT -203.960 88.800 -199.940 90.180 ;
        RECT -194.040 88.800 -190.020 90.180 ;
        RECT -184.120 88.800 -180.100 90.180 ;
        RECT -174.200 88.800 -170.180 90.180 ;
        RECT -164.280 88.800 -160.260 90.180 ;
        RECT -154.360 88.800 -150.340 90.180 ;
        RECT -144.440 88.800 -140.420 90.180 ;
        RECT -134.520 88.800 -130.500 90.180 ;
        RECT -124.600 88.800 -120.580 90.180 ;
        RECT -114.680 88.800 -110.660 90.180 ;
        RECT -104.760 88.800 -100.740 90.180 ;
        RECT -94.840 88.800 -90.820 90.180 ;
        RECT -84.920 88.800 -80.900 90.180 ;
        RECT -75.000 88.800 -70.980 90.180 ;
        RECT -65.080 88.800 -61.060 90.180 ;
        RECT -55.160 88.800 -51.140 90.180 ;
        RECT -45.240 88.800 -41.220 90.180 ;
        RECT -35.320 88.800 -31.300 90.180 ;
        RECT -25.400 88.800 -21.380 90.180 ;
        RECT -15.480 88.800 -11.460 90.180 ;
        RECT -5.560 88.800 -1.540 90.180 ;
        RECT 4.360 88.800 8.380 90.180 ;
        RECT 14.280 88.800 18.300 90.180 ;
      LAYER via ;
        RECT -287.700 94.070 -287.425 94.335 ;
        RECT -277.780 94.070 -277.505 94.335 ;
        RECT -267.860 94.070 -267.585 94.335 ;
        RECT -257.940 94.070 -257.665 94.335 ;
        RECT -248.020 94.070 -247.745 94.335 ;
        RECT -238.100 94.070 -237.825 94.335 ;
        RECT -228.180 94.070 -227.905 94.335 ;
        RECT -218.260 94.070 -217.985 94.335 ;
        RECT -208.340 94.070 -208.065 94.335 ;
        RECT -198.420 94.070 -198.145 94.335 ;
        RECT -188.500 94.070 -188.225 94.335 ;
        RECT -178.580 94.070 -178.305 94.335 ;
        RECT -168.660 94.070 -168.385 94.335 ;
        RECT -158.740 94.070 -158.465 94.335 ;
        RECT -148.820 94.070 -148.545 94.335 ;
        RECT -138.900 94.070 -138.625 94.335 ;
        RECT -128.980 94.070 -128.705 94.335 ;
        RECT -119.060 94.070 -118.785 94.335 ;
        RECT -109.140 94.070 -108.865 94.335 ;
        RECT -99.220 94.070 -98.945 94.335 ;
        RECT -89.300 94.070 -89.025 94.335 ;
        RECT -79.380 94.070 -79.105 94.335 ;
        RECT -69.460 94.070 -69.185 94.335 ;
        RECT -59.540 94.070 -59.265 94.335 ;
        RECT -49.620 94.070 -49.345 94.335 ;
        RECT -39.700 94.070 -39.425 94.335 ;
        RECT -29.780 94.070 -29.505 94.335 ;
        RECT -19.860 94.070 -19.585 94.335 ;
        RECT -9.940 94.070 -9.665 94.335 ;
        RECT -0.020 94.070 0.255 94.335 ;
        RECT 9.900 94.070 10.175 94.335 ;
        RECT 19.820 94.070 20.095 94.335 ;
        RECT -280.530 93.200 -280.255 93.465 ;
        RECT -280.060 93.200 -279.785 93.465 ;
        RECT -270.610 93.200 -270.335 93.465 ;
        RECT -270.140 93.200 -269.865 93.465 ;
        RECT -260.690 93.200 -260.415 93.465 ;
        RECT -260.220 93.200 -259.945 93.465 ;
        RECT -250.770 93.200 -250.495 93.465 ;
        RECT -250.300 93.200 -250.025 93.465 ;
        RECT -240.850 93.200 -240.575 93.465 ;
        RECT -240.380 93.200 -240.105 93.465 ;
        RECT -230.930 93.200 -230.655 93.465 ;
        RECT -230.460 93.200 -230.185 93.465 ;
        RECT -221.010 93.200 -220.735 93.465 ;
        RECT -220.540 93.200 -220.265 93.465 ;
        RECT -211.090 93.200 -210.815 93.465 ;
        RECT -210.620 93.200 -210.345 93.465 ;
        RECT -201.170 93.200 -200.895 93.465 ;
        RECT -200.700 93.200 -200.425 93.465 ;
        RECT -191.250 93.200 -190.975 93.465 ;
        RECT -190.780 93.200 -190.505 93.465 ;
        RECT -181.330 93.200 -181.055 93.465 ;
        RECT -180.860 93.200 -180.585 93.465 ;
        RECT -171.410 93.200 -171.135 93.465 ;
        RECT -170.940 93.200 -170.665 93.465 ;
        RECT -161.490 93.200 -161.215 93.465 ;
        RECT -161.020 93.200 -160.745 93.465 ;
        RECT -151.570 93.200 -151.295 93.465 ;
        RECT -151.100 93.200 -150.825 93.465 ;
        RECT -141.650 93.200 -141.375 93.465 ;
        RECT -141.180 93.200 -140.905 93.465 ;
        RECT -131.730 93.200 -131.455 93.465 ;
        RECT -131.260 93.200 -130.985 93.465 ;
        RECT -121.810 93.200 -121.535 93.465 ;
        RECT -121.340 93.200 -121.065 93.465 ;
        RECT -111.890 93.200 -111.615 93.465 ;
        RECT -111.420 93.200 -111.145 93.465 ;
        RECT -101.970 93.200 -101.695 93.465 ;
        RECT -101.500 93.200 -101.225 93.465 ;
        RECT -92.050 93.200 -91.775 93.465 ;
        RECT -91.580 93.200 -91.305 93.465 ;
        RECT -82.130 93.200 -81.855 93.465 ;
        RECT -81.660 93.200 -81.385 93.465 ;
        RECT -72.210 93.200 -71.935 93.465 ;
        RECT -71.740 93.200 -71.465 93.465 ;
        RECT -62.290 93.200 -62.015 93.465 ;
        RECT -61.820 93.200 -61.545 93.465 ;
        RECT -52.370 93.200 -52.095 93.465 ;
        RECT -51.900 93.200 -51.625 93.465 ;
        RECT -42.450 93.200 -42.175 93.465 ;
        RECT -41.980 93.200 -41.705 93.465 ;
        RECT -32.530 93.200 -32.255 93.465 ;
        RECT -32.060 93.200 -31.785 93.465 ;
        RECT -22.610 93.200 -22.335 93.465 ;
        RECT -22.140 93.200 -21.865 93.465 ;
        RECT -12.690 93.200 -12.415 93.465 ;
        RECT -12.220 93.200 -11.945 93.465 ;
        RECT -2.770 93.200 -2.495 93.465 ;
        RECT -2.300 93.200 -2.025 93.465 ;
        RECT 7.150 93.200 7.425 93.465 ;
        RECT 7.620 93.200 7.895 93.465 ;
        RECT 17.070 93.200 17.345 93.465 ;
        RECT 17.540 93.200 17.815 93.465 ;
        RECT -287.790 90.470 -287.515 90.735 ;
        RECT -287.330 90.480 -287.055 90.745 ;
        RECT -277.870 90.470 -277.595 90.735 ;
        RECT -277.410 90.480 -277.135 90.745 ;
        RECT -267.950 90.470 -267.675 90.735 ;
        RECT -267.490 90.480 -267.215 90.745 ;
        RECT -258.030 90.470 -257.755 90.735 ;
        RECT -257.570 90.480 -257.295 90.745 ;
        RECT -248.110 90.470 -247.835 90.735 ;
        RECT -247.650 90.480 -247.375 90.745 ;
        RECT -238.190 90.470 -237.915 90.735 ;
        RECT -237.730 90.480 -237.455 90.745 ;
        RECT -228.270 90.470 -227.995 90.735 ;
        RECT -227.810 90.480 -227.535 90.745 ;
        RECT -218.350 90.470 -218.075 90.735 ;
        RECT -217.890 90.480 -217.615 90.745 ;
        RECT -208.430 90.470 -208.155 90.735 ;
        RECT -207.970 90.480 -207.695 90.745 ;
        RECT -198.510 90.470 -198.235 90.735 ;
        RECT -198.050 90.480 -197.775 90.745 ;
        RECT -188.590 90.470 -188.315 90.735 ;
        RECT -188.130 90.480 -187.855 90.745 ;
        RECT -178.670 90.470 -178.395 90.735 ;
        RECT -178.210 90.480 -177.935 90.745 ;
        RECT -168.750 90.470 -168.475 90.735 ;
        RECT -168.290 90.480 -168.015 90.745 ;
        RECT -158.830 90.470 -158.555 90.735 ;
        RECT -158.370 90.480 -158.095 90.745 ;
        RECT -148.910 90.470 -148.635 90.735 ;
        RECT -148.450 90.480 -148.175 90.745 ;
        RECT -138.990 90.470 -138.715 90.735 ;
        RECT -138.530 90.480 -138.255 90.745 ;
        RECT -129.070 90.470 -128.795 90.735 ;
        RECT -128.610 90.480 -128.335 90.745 ;
        RECT -119.150 90.470 -118.875 90.735 ;
        RECT -118.690 90.480 -118.415 90.745 ;
        RECT -109.230 90.470 -108.955 90.735 ;
        RECT -108.770 90.480 -108.495 90.745 ;
        RECT -99.310 90.470 -99.035 90.735 ;
        RECT -98.850 90.480 -98.575 90.745 ;
        RECT -89.390 90.470 -89.115 90.735 ;
        RECT -88.930 90.480 -88.655 90.745 ;
        RECT -79.470 90.470 -79.195 90.735 ;
        RECT -79.010 90.480 -78.735 90.745 ;
        RECT -69.550 90.470 -69.275 90.735 ;
        RECT -69.090 90.480 -68.815 90.745 ;
        RECT -59.630 90.470 -59.355 90.735 ;
        RECT -59.170 90.480 -58.895 90.745 ;
        RECT -49.710 90.470 -49.435 90.735 ;
        RECT -49.250 90.480 -48.975 90.745 ;
        RECT -39.790 90.470 -39.515 90.735 ;
        RECT -39.330 90.480 -39.055 90.745 ;
        RECT -29.870 90.470 -29.595 90.735 ;
        RECT -29.410 90.480 -29.135 90.745 ;
        RECT -19.950 90.470 -19.675 90.735 ;
        RECT -19.490 90.480 -19.215 90.745 ;
        RECT -10.030 90.470 -9.755 90.735 ;
        RECT -9.570 90.480 -9.295 90.745 ;
        RECT -0.110 90.470 0.165 90.735 ;
        RECT 0.350 90.480 0.625 90.745 ;
        RECT 9.810 90.470 10.085 90.735 ;
        RECT 10.270 90.480 10.545 90.745 ;
        RECT 19.730 90.470 20.005 90.735 ;
        RECT 20.190 90.480 20.465 90.745 ;
        RECT -280.140 89.710 -279.865 89.975 ;
        RECT -270.220 89.710 -269.945 89.975 ;
        RECT -260.300 89.710 -260.025 89.975 ;
        RECT -250.380 89.710 -250.105 89.975 ;
        RECT -240.460 89.710 -240.185 89.975 ;
        RECT -230.540 89.710 -230.265 89.975 ;
        RECT -220.620 89.710 -220.345 89.975 ;
        RECT -210.700 89.710 -210.425 89.975 ;
        RECT -200.780 89.710 -200.505 89.975 ;
        RECT -190.860 89.710 -190.585 89.975 ;
        RECT -180.940 89.710 -180.665 89.975 ;
        RECT -171.020 89.710 -170.745 89.975 ;
        RECT -161.100 89.710 -160.825 89.975 ;
        RECT -151.180 89.710 -150.905 89.975 ;
        RECT -141.260 89.710 -140.985 89.975 ;
        RECT -131.340 89.710 -131.065 89.975 ;
        RECT -121.420 89.710 -121.145 89.975 ;
        RECT -111.500 89.710 -111.225 89.975 ;
        RECT -101.580 89.710 -101.305 89.975 ;
        RECT -91.660 89.710 -91.385 89.975 ;
        RECT -81.740 89.710 -81.465 89.975 ;
        RECT -71.820 89.710 -71.545 89.975 ;
        RECT -61.900 89.710 -61.625 89.975 ;
        RECT -51.980 89.710 -51.705 89.975 ;
        RECT -42.060 89.710 -41.785 89.975 ;
        RECT -32.140 89.710 -31.865 89.975 ;
        RECT -22.220 89.710 -21.945 89.975 ;
        RECT -12.300 89.710 -12.025 89.975 ;
        RECT -2.380 89.710 -2.105 89.975 ;
        RECT 7.540 89.710 7.815 89.975 ;
        RECT 17.460 89.710 17.735 89.975 ;
      LAYER met2 ;
        RECT -288.280 93.760 -287.110 94.560 ;
        RECT -278.360 93.760 -277.190 94.560 ;
        RECT -268.440 93.760 -267.270 94.560 ;
        RECT -258.520 93.760 -257.350 94.560 ;
        RECT -248.600 93.760 -247.430 94.560 ;
        RECT -238.680 93.760 -237.510 94.560 ;
        RECT -228.760 93.760 -227.590 94.560 ;
        RECT -218.840 93.760 -217.670 94.560 ;
        RECT -208.920 93.760 -207.750 94.560 ;
        RECT -199.000 93.760 -197.830 94.560 ;
        RECT -189.080 93.760 -187.910 94.560 ;
        RECT -179.160 93.760 -177.990 94.560 ;
        RECT -169.240 93.760 -168.070 94.560 ;
        RECT -159.320 93.760 -158.150 94.560 ;
        RECT -149.400 93.760 -148.230 94.560 ;
        RECT -139.480 93.760 -138.310 94.560 ;
        RECT -129.560 93.760 -128.390 94.560 ;
        RECT -119.640 93.760 -118.470 94.560 ;
        RECT -109.720 93.760 -108.550 94.560 ;
        RECT -99.800 93.760 -98.630 94.560 ;
        RECT -89.880 93.760 -88.710 94.560 ;
        RECT -79.960 93.760 -78.790 94.560 ;
        RECT -70.040 93.760 -68.870 94.560 ;
        RECT -60.120 93.760 -58.950 94.560 ;
        RECT -50.200 93.760 -49.030 94.560 ;
        RECT -40.280 93.760 -39.110 94.560 ;
        RECT -30.360 93.760 -29.190 94.560 ;
        RECT -20.440 93.760 -19.270 94.560 ;
        RECT -10.520 93.760 -9.350 94.560 ;
        RECT -0.600 93.760 0.570 94.560 ;
        RECT 9.320 93.760 10.490 94.560 ;
        RECT 19.240 93.760 20.410 94.560 ;
        RECT -280.620 93.090 -279.700 93.570 ;
        RECT -270.700 93.090 -269.780 93.570 ;
        RECT -260.780 93.090 -259.860 93.570 ;
        RECT -250.860 93.090 -249.940 93.570 ;
        RECT -240.940 93.090 -240.020 93.570 ;
        RECT -231.020 93.090 -230.100 93.570 ;
        RECT -221.100 93.090 -220.180 93.570 ;
        RECT -211.180 93.090 -210.260 93.570 ;
        RECT -201.260 93.090 -200.340 93.570 ;
        RECT -191.340 93.090 -190.420 93.570 ;
        RECT -181.420 93.090 -180.500 93.570 ;
        RECT -171.500 93.090 -170.580 93.570 ;
        RECT -161.580 93.090 -160.660 93.570 ;
        RECT -151.660 93.090 -150.740 93.570 ;
        RECT -141.740 93.090 -140.820 93.570 ;
        RECT -131.820 93.090 -130.900 93.570 ;
        RECT -121.900 93.090 -120.980 93.570 ;
        RECT -111.980 93.090 -111.060 93.570 ;
        RECT -102.060 93.090 -101.140 93.570 ;
        RECT -92.140 93.090 -91.220 93.570 ;
        RECT -82.220 93.090 -81.300 93.570 ;
        RECT -72.300 93.090 -71.380 93.570 ;
        RECT -62.380 93.090 -61.460 93.570 ;
        RECT -52.460 93.090 -51.540 93.570 ;
        RECT -42.540 93.090 -41.620 93.570 ;
        RECT -32.620 93.090 -31.700 93.570 ;
        RECT -22.700 93.090 -21.780 93.570 ;
        RECT -12.780 93.090 -11.860 93.570 ;
        RECT -2.860 93.090 -1.940 93.570 ;
        RECT 7.060 93.090 7.980 93.570 ;
        RECT 16.980 93.090 17.900 93.570 ;
        RECT -287.880 90.370 -286.960 90.850 ;
        RECT -277.960 90.370 -277.040 90.850 ;
        RECT -268.040 90.370 -267.120 90.850 ;
        RECT -258.120 90.370 -257.200 90.850 ;
        RECT -248.200 90.370 -247.280 90.850 ;
        RECT -238.280 90.370 -237.360 90.850 ;
        RECT -228.360 90.370 -227.440 90.850 ;
        RECT -218.440 90.370 -217.520 90.850 ;
        RECT -208.520 90.370 -207.600 90.850 ;
        RECT -198.600 90.370 -197.680 90.850 ;
        RECT -188.680 90.370 -187.760 90.850 ;
        RECT -178.760 90.370 -177.840 90.850 ;
        RECT -168.840 90.370 -167.920 90.850 ;
        RECT -158.920 90.370 -158.000 90.850 ;
        RECT -149.000 90.370 -148.080 90.850 ;
        RECT -139.080 90.370 -138.160 90.850 ;
        RECT -129.160 90.370 -128.240 90.850 ;
        RECT -119.240 90.370 -118.320 90.850 ;
        RECT -109.320 90.370 -108.400 90.850 ;
        RECT -99.400 90.370 -98.480 90.850 ;
        RECT -89.480 90.370 -88.560 90.850 ;
        RECT -79.560 90.370 -78.640 90.850 ;
        RECT -69.640 90.370 -68.720 90.850 ;
        RECT -59.720 90.370 -58.800 90.850 ;
        RECT -49.800 90.370 -48.880 90.850 ;
        RECT -39.880 90.370 -38.960 90.850 ;
        RECT -29.960 90.370 -29.040 90.850 ;
        RECT -20.040 90.370 -19.120 90.850 ;
        RECT -10.120 90.370 -9.200 90.850 ;
        RECT -0.200 90.370 0.720 90.850 ;
        RECT 9.720 90.370 10.640 90.850 ;
        RECT 19.640 90.370 20.560 90.850 ;
        RECT -280.460 89.390 -279.290 90.190 ;
        RECT -270.540 89.390 -269.370 90.190 ;
        RECT -260.620 89.390 -259.450 90.190 ;
        RECT -250.700 89.390 -249.530 90.190 ;
        RECT -240.780 89.390 -239.610 90.190 ;
        RECT -230.860 89.390 -229.690 90.190 ;
        RECT -220.940 89.390 -219.770 90.190 ;
        RECT -211.020 89.390 -209.850 90.190 ;
        RECT -201.100 89.390 -199.930 90.190 ;
        RECT -191.180 89.390 -190.010 90.190 ;
        RECT -181.260 89.390 -180.090 90.190 ;
        RECT -171.340 89.390 -170.170 90.190 ;
        RECT -161.420 89.390 -160.250 90.190 ;
        RECT -151.500 89.390 -150.330 90.190 ;
        RECT -141.580 89.390 -140.410 90.190 ;
        RECT -131.660 89.390 -130.490 90.190 ;
        RECT -121.740 89.390 -120.570 90.190 ;
        RECT -111.820 89.390 -110.650 90.190 ;
        RECT -101.900 89.390 -100.730 90.190 ;
        RECT -91.980 89.390 -90.810 90.190 ;
        RECT -82.060 89.390 -80.890 90.190 ;
        RECT -72.140 89.390 -70.970 90.190 ;
        RECT -62.220 89.390 -61.050 90.190 ;
        RECT -52.300 89.390 -51.130 90.190 ;
        RECT -42.380 89.390 -41.210 90.190 ;
        RECT -32.460 89.390 -31.290 90.190 ;
        RECT -22.540 89.390 -21.370 90.190 ;
        RECT -12.620 89.390 -11.450 90.190 ;
        RECT -2.700 89.390 -1.530 90.190 ;
        RECT 7.220 89.390 8.390 90.190 ;
        RECT 17.140 89.390 18.310 90.190 ;
      LAYER via2 ;
        RECT -287.710 94.060 -287.420 94.340 ;
        RECT -277.790 94.060 -277.500 94.340 ;
        RECT -267.870 94.060 -267.580 94.340 ;
        RECT -257.950 94.060 -257.660 94.340 ;
        RECT -248.030 94.060 -247.740 94.340 ;
        RECT -238.110 94.060 -237.820 94.340 ;
        RECT -228.190 94.060 -227.900 94.340 ;
        RECT -218.270 94.060 -217.980 94.340 ;
        RECT -208.350 94.060 -208.060 94.340 ;
        RECT -198.430 94.060 -198.140 94.340 ;
        RECT -188.510 94.060 -188.220 94.340 ;
        RECT -178.590 94.060 -178.300 94.340 ;
        RECT -168.670 94.060 -168.380 94.340 ;
        RECT -158.750 94.060 -158.460 94.340 ;
        RECT -148.830 94.060 -148.540 94.340 ;
        RECT -138.910 94.060 -138.620 94.340 ;
        RECT -128.990 94.060 -128.700 94.340 ;
        RECT -119.070 94.060 -118.780 94.340 ;
        RECT -109.150 94.060 -108.860 94.340 ;
        RECT -99.230 94.060 -98.940 94.340 ;
        RECT -89.310 94.060 -89.020 94.340 ;
        RECT -79.390 94.060 -79.100 94.340 ;
        RECT -69.470 94.060 -69.180 94.340 ;
        RECT -59.550 94.060 -59.260 94.340 ;
        RECT -49.630 94.060 -49.340 94.340 ;
        RECT -39.710 94.060 -39.420 94.340 ;
        RECT -29.790 94.060 -29.500 94.340 ;
        RECT -19.870 94.060 -19.580 94.340 ;
        RECT -9.950 94.060 -9.660 94.340 ;
        RECT -0.030 94.060 0.260 94.340 ;
        RECT 9.890 94.060 10.180 94.340 ;
        RECT 19.810 94.060 20.100 94.340 ;
        RECT -280.540 93.190 -280.250 93.470 ;
        RECT -280.070 93.190 -279.780 93.470 ;
        RECT -270.620 93.190 -270.330 93.470 ;
        RECT -270.150 93.190 -269.860 93.470 ;
        RECT -260.700 93.190 -260.410 93.470 ;
        RECT -260.230 93.190 -259.940 93.470 ;
        RECT -250.780 93.190 -250.490 93.470 ;
        RECT -250.310 93.190 -250.020 93.470 ;
        RECT -240.860 93.190 -240.570 93.470 ;
        RECT -240.390 93.190 -240.100 93.470 ;
        RECT -230.940 93.190 -230.650 93.470 ;
        RECT -230.470 93.190 -230.180 93.470 ;
        RECT -221.020 93.190 -220.730 93.470 ;
        RECT -220.550 93.190 -220.260 93.470 ;
        RECT -211.100 93.190 -210.810 93.470 ;
        RECT -210.630 93.190 -210.340 93.470 ;
        RECT -201.180 93.190 -200.890 93.470 ;
        RECT -200.710 93.190 -200.420 93.470 ;
        RECT -191.260 93.190 -190.970 93.470 ;
        RECT -190.790 93.190 -190.500 93.470 ;
        RECT -181.340 93.190 -181.050 93.470 ;
        RECT -180.870 93.190 -180.580 93.470 ;
        RECT -171.420 93.190 -171.130 93.470 ;
        RECT -170.950 93.190 -170.660 93.470 ;
        RECT -161.500 93.190 -161.210 93.470 ;
        RECT -161.030 93.190 -160.740 93.470 ;
        RECT -151.580 93.190 -151.290 93.470 ;
        RECT -151.110 93.190 -150.820 93.470 ;
        RECT -141.660 93.190 -141.370 93.470 ;
        RECT -141.190 93.190 -140.900 93.470 ;
        RECT -131.740 93.190 -131.450 93.470 ;
        RECT -131.270 93.190 -130.980 93.470 ;
        RECT -121.820 93.190 -121.530 93.470 ;
        RECT -121.350 93.190 -121.060 93.470 ;
        RECT -111.900 93.190 -111.610 93.470 ;
        RECT -111.430 93.190 -111.140 93.470 ;
        RECT -101.980 93.190 -101.690 93.470 ;
        RECT -101.510 93.190 -101.220 93.470 ;
        RECT -92.060 93.190 -91.770 93.470 ;
        RECT -91.590 93.190 -91.300 93.470 ;
        RECT -82.140 93.190 -81.850 93.470 ;
        RECT -81.670 93.190 -81.380 93.470 ;
        RECT -72.220 93.190 -71.930 93.470 ;
        RECT -71.750 93.190 -71.460 93.470 ;
        RECT -62.300 93.190 -62.010 93.470 ;
        RECT -61.830 93.190 -61.540 93.470 ;
        RECT -52.380 93.190 -52.090 93.470 ;
        RECT -51.910 93.190 -51.620 93.470 ;
        RECT -42.460 93.190 -42.170 93.470 ;
        RECT -41.990 93.190 -41.700 93.470 ;
        RECT -32.540 93.190 -32.250 93.470 ;
        RECT -32.070 93.190 -31.780 93.470 ;
        RECT -22.620 93.190 -22.330 93.470 ;
        RECT -22.150 93.190 -21.860 93.470 ;
        RECT -12.700 93.190 -12.410 93.470 ;
        RECT -12.230 93.190 -11.940 93.470 ;
        RECT -2.780 93.190 -2.490 93.470 ;
        RECT -2.310 93.190 -2.020 93.470 ;
        RECT 7.140 93.190 7.430 93.470 ;
        RECT 7.610 93.190 7.900 93.470 ;
        RECT 17.060 93.190 17.350 93.470 ;
        RECT 17.530 93.190 17.820 93.470 ;
        RECT -287.800 90.460 -287.510 90.740 ;
        RECT -287.340 90.470 -287.050 90.750 ;
        RECT -277.880 90.460 -277.590 90.740 ;
        RECT -277.420 90.470 -277.130 90.750 ;
        RECT -267.960 90.460 -267.670 90.740 ;
        RECT -267.500 90.470 -267.210 90.750 ;
        RECT -258.040 90.460 -257.750 90.740 ;
        RECT -257.580 90.470 -257.290 90.750 ;
        RECT -248.120 90.460 -247.830 90.740 ;
        RECT -247.660 90.470 -247.370 90.750 ;
        RECT -238.200 90.460 -237.910 90.740 ;
        RECT -237.740 90.470 -237.450 90.750 ;
        RECT -228.280 90.460 -227.990 90.740 ;
        RECT -227.820 90.470 -227.530 90.750 ;
        RECT -218.360 90.460 -218.070 90.740 ;
        RECT -217.900 90.470 -217.610 90.750 ;
        RECT -208.440 90.460 -208.150 90.740 ;
        RECT -207.980 90.470 -207.690 90.750 ;
        RECT -198.520 90.460 -198.230 90.740 ;
        RECT -198.060 90.470 -197.770 90.750 ;
        RECT -188.600 90.460 -188.310 90.740 ;
        RECT -188.140 90.470 -187.850 90.750 ;
        RECT -178.680 90.460 -178.390 90.740 ;
        RECT -178.220 90.470 -177.930 90.750 ;
        RECT -168.760 90.460 -168.470 90.740 ;
        RECT -168.300 90.470 -168.010 90.750 ;
        RECT -158.840 90.460 -158.550 90.740 ;
        RECT -158.380 90.470 -158.090 90.750 ;
        RECT -148.920 90.460 -148.630 90.740 ;
        RECT -148.460 90.470 -148.170 90.750 ;
        RECT -139.000 90.460 -138.710 90.740 ;
        RECT -138.540 90.470 -138.250 90.750 ;
        RECT -129.080 90.460 -128.790 90.740 ;
        RECT -128.620 90.470 -128.330 90.750 ;
        RECT -119.160 90.460 -118.870 90.740 ;
        RECT -118.700 90.470 -118.410 90.750 ;
        RECT -109.240 90.460 -108.950 90.740 ;
        RECT -108.780 90.470 -108.490 90.750 ;
        RECT -99.320 90.460 -99.030 90.740 ;
        RECT -98.860 90.470 -98.570 90.750 ;
        RECT -89.400 90.460 -89.110 90.740 ;
        RECT -88.940 90.470 -88.650 90.750 ;
        RECT -79.480 90.460 -79.190 90.740 ;
        RECT -79.020 90.470 -78.730 90.750 ;
        RECT -69.560 90.460 -69.270 90.740 ;
        RECT -69.100 90.470 -68.810 90.750 ;
        RECT -59.640 90.460 -59.350 90.740 ;
        RECT -59.180 90.470 -58.890 90.750 ;
        RECT -49.720 90.460 -49.430 90.740 ;
        RECT -49.260 90.470 -48.970 90.750 ;
        RECT -39.800 90.460 -39.510 90.740 ;
        RECT -39.340 90.470 -39.050 90.750 ;
        RECT -29.880 90.460 -29.590 90.740 ;
        RECT -29.420 90.470 -29.130 90.750 ;
        RECT -19.960 90.460 -19.670 90.740 ;
        RECT -19.500 90.470 -19.210 90.750 ;
        RECT -10.040 90.460 -9.750 90.740 ;
        RECT -9.580 90.470 -9.290 90.750 ;
        RECT -0.120 90.460 0.170 90.740 ;
        RECT 0.340 90.470 0.630 90.750 ;
        RECT 9.800 90.460 10.090 90.740 ;
        RECT 10.260 90.470 10.550 90.750 ;
        RECT 19.720 90.460 20.010 90.740 ;
        RECT 20.180 90.470 20.470 90.750 ;
        RECT -280.150 89.700 -279.860 89.980 ;
        RECT -270.230 89.700 -269.940 89.980 ;
        RECT -260.310 89.700 -260.020 89.980 ;
        RECT -250.390 89.700 -250.100 89.980 ;
        RECT -240.470 89.700 -240.180 89.980 ;
        RECT -230.550 89.700 -230.260 89.980 ;
        RECT -220.630 89.700 -220.340 89.980 ;
        RECT -210.710 89.700 -210.420 89.980 ;
        RECT -200.790 89.700 -200.500 89.980 ;
        RECT -190.870 89.700 -190.580 89.980 ;
        RECT -180.950 89.700 -180.660 89.980 ;
        RECT -171.030 89.700 -170.740 89.980 ;
        RECT -161.110 89.700 -160.820 89.980 ;
        RECT -151.190 89.700 -150.900 89.980 ;
        RECT -141.270 89.700 -140.980 89.980 ;
        RECT -131.350 89.700 -131.060 89.980 ;
        RECT -121.430 89.700 -121.140 89.980 ;
        RECT -111.510 89.700 -111.220 89.980 ;
        RECT -101.590 89.700 -101.300 89.980 ;
        RECT -91.670 89.700 -91.380 89.980 ;
        RECT -81.750 89.700 -81.460 89.980 ;
        RECT -71.830 89.700 -71.540 89.980 ;
        RECT -61.910 89.700 -61.620 89.980 ;
        RECT -51.990 89.700 -51.700 89.980 ;
        RECT -42.070 89.700 -41.780 89.980 ;
        RECT -32.150 89.700 -31.860 89.980 ;
        RECT -22.230 89.700 -21.940 89.980 ;
        RECT -12.310 89.700 -12.020 89.980 ;
        RECT -2.390 89.700 -2.100 89.980 ;
        RECT 7.530 89.700 7.820 89.980 ;
        RECT 17.450 89.700 17.740 89.980 ;
      LAYER met3 ;
        RECT -288.280 93.760 -287.110 94.560 ;
        RECT -278.360 93.760 -277.190 94.560 ;
        RECT -268.440 93.760 -267.270 94.560 ;
        RECT -258.520 93.760 -257.350 94.560 ;
        RECT -248.600 93.760 -247.430 94.560 ;
        RECT -238.680 93.760 -237.510 94.560 ;
        RECT -228.760 93.760 -227.590 94.560 ;
        RECT -218.840 93.760 -217.670 94.560 ;
        RECT -208.920 93.760 -207.750 94.560 ;
        RECT -199.000 93.760 -197.830 94.560 ;
        RECT -189.080 93.760 -187.910 94.560 ;
        RECT -179.160 93.760 -177.990 94.560 ;
        RECT -169.240 93.760 -168.070 94.560 ;
        RECT -159.320 93.760 -158.150 94.560 ;
        RECT -149.400 93.760 -148.230 94.560 ;
        RECT -139.480 93.760 -138.310 94.560 ;
        RECT -129.560 93.760 -128.390 94.560 ;
        RECT -119.640 93.760 -118.470 94.560 ;
        RECT -109.720 93.760 -108.550 94.560 ;
        RECT -99.800 93.760 -98.630 94.560 ;
        RECT -89.880 93.760 -88.710 94.560 ;
        RECT -79.960 93.760 -78.790 94.560 ;
        RECT -70.040 93.760 -68.870 94.560 ;
        RECT -60.120 93.760 -58.950 94.560 ;
        RECT -50.200 93.760 -49.030 94.560 ;
        RECT -40.280 93.760 -39.110 94.560 ;
        RECT -30.360 93.760 -29.190 94.560 ;
        RECT -20.440 93.760 -19.270 94.560 ;
        RECT -10.520 93.760 -9.350 94.560 ;
        RECT -0.600 93.760 0.570 94.560 ;
        RECT 9.320 93.760 10.490 94.560 ;
        RECT 19.240 93.760 20.410 94.560 ;
        RECT -280.620 93.090 -279.700 93.570 ;
        RECT -270.700 93.090 -269.780 93.570 ;
        RECT -260.780 93.090 -259.860 93.570 ;
        RECT -250.860 93.090 -249.940 93.570 ;
        RECT -240.940 93.090 -240.020 93.570 ;
        RECT -231.020 93.090 -230.100 93.570 ;
        RECT -221.100 93.090 -220.180 93.570 ;
        RECT -211.180 93.090 -210.260 93.570 ;
        RECT -201.260 93.090 -200.340 93.570 ;
        RECT -191.340 93.090 -190.420 93.570 ;
        RECT -181.420 93.090 -180.500 93.570 ;
        RECT -171.500 93.090 -170.580 93.570 ;
        RECT -161.580 93.090 -160.660 93.570 ;
        RECT -151.660 93.090 -150.740 93.570 ;
        RECT -141.740 93.090 -140.820 93.570 ;
        RECT -131.820 93.090 -130.900 93.570 ;
        RECT -121.900 93.090 -120.980 93.570 ;
        RECT -111.980 93.090 -111.060 93.570 ;
        RECT -102.060 93.090 -101.140 93.570 ;
        RECT -92.140 93.090 -91.220 93.570 ;
        RECT -82.220 93.090 -81.300 93.570 ;
        RECT -72.300 93.090 -71.380 93.570 ;
        RECT -62.380 93.090 -61.460 93.570 ;
        RECT -52.460 93.090 -51.540 93.570 ;
        RECT -42.540 93.090 -41.620 93.570 ;
        RECT -32.620 93.090 -31.700 93.570 ;
        RECT -22.700 93.090 -21.780 93.570 ;
        RECT -12.780 93.090 -11.860 93.570 ;
        RECT -2.860 93.090 -1.940 93.570 ;
        RECT 7.060 93.090 7.980 93.570 ;
        RECT 16.980 93.090 17.900 93.570 ;
        RECT -287.880 90.370 -286.960 90.850 ;
        RECT -277.960 90.370 -277.040 90.850 ;
        RECT -268.040 90.370 -267.120 90.850 ;
        RECT -258.120 90.370 -257.200 90.850 ;
        RECT -248.200 90.370 -247.280 90.850 ;
        RECT -238.280 90.370 -237.360 90.850 ;
        RECT -228.360 90.370 -227.440 90.850 ;
        RECT -218.440 90.370 -217.520 90.850 ;
        RECT -208.520 90.370 -207.600 90.850 ;
        RECT -198.600 90.370 -197.680 90.850 ;
        RECT -188.680 90.370 -187.760 90.850 ;
        RECT -178.760 90.370 -177.840 90.850 ;
        RECT -168.840 90.370 -167.920 90.850 ;
        RECT -158.920 90.370 -158.000 90.850 ;
        RECT -149.000 90.370 -148.080 90.850 ;
        RECT -139.080 90.370 -138.160 90.850 ;
        RECT -129.160 90.370 -128.240 90.850 ;
        RECT -119.240 90.370 -118.320 90.850 ;
        RECT -109.320 90.370 -108.400 90.850 ;
        RECT -99.400 90.370 -98.480 90.850 ;
        RECT -89.480 90.370 -88.560 90.850 ;
        RECT -79.560 90.370 -78.640 90.850 ;
        RECT -69.640 90.370 -68.720 90.850 ;
        RECT -59.720 90.370 -58.800 90.850 ;
        RECT -49.800 90.370 -48.880 90.850 ;
        RECT -39.880 90.370 -38.960 90.850 ;
        RECT -29.960 90.370 -29.040 90.850 ;
        RECT -20.040 90.370 -19.120 90.850 ;
        RECT -10.120 90.370 -9.200 90.850 ;
        RECT -0.200 90.370 0.720 90.850 ;
        RECT 9.720 90.370 10.640 90.850 ;
        RECT 19.640 90.370 20.560 90.850 ;
        RECT -280.460 89.390 -279.290 90.190 ;
        RECT -270.540 89.390 -269.370 90.190 ;
        RECT -260.620 89.390 -259.450 90.190 ;
        RECT -250.700 89.390 -249.530 90.190 ;
        RECT -240.780 89.390 -239.610 90.190 ;
        RECT -230.860 89.390 -229.690 90.190 ;
        RECT -220.940 89.390 -219.770 90.190 ;
        RECT -211.020 89.390 -209.850 90.190 ;
        RECT -201.100 89.390 -199.930 90.190 ;
        RECT -191.180 89.390 -190.010 90.190 ;
        RECT -181.260 89.390 -180.090 90.190 ;
        RECT -171.340 89.390 -170.170 90.190 ;
        RECT -161.420 89.390 -160.250 90.190 ;
        RECT -151.500 89.390 -150.330 90.190 ;
        RECT -141.580 89.390 -140.410 90.190 ;
        RECT -131.660 89.390 -130.490 90.190 ;
        RECT -121.740 89.390 -120.570 90.190 ;
        RECT -111.820 89.390 -110.650 90.190 ;
        RECT -101.900 89.390 -100.730 90.190 ;
        RECT -91.980 89.390 -90.810 90.190 ;
        RECT -82.060 89.390 -80.890 90.190 ;
        RECT -72.140 89.390 -70.970 90.190 ;
        RECT -62.220 89.390 -61.050 90.190 ;
        RECT -52.300 89.390 -51.130 90.190 ;
        RECT -42.380 89.390 -41.210 90.190 ;
        RECT -32.460 89.390 -31.290 90.190 ;
        RECT -22.540 89.390 -21.370 90.190 ;
        RECT -12.620 89.390 -11.450 90.190 ;
        RECT -2.700 89.390 -1.530 90.190 ;
        RECT 7.220 89.390 8.390 90.190 ;
        RECT 17.140 89.390 18.310 90.190 ;
      LAYER via3 ;
        RECT -287.740 94.030 -287.400 94.360 ;
        RECT -277.820 94.030 -277.480 94.360 ;
        RECT -267.900 94.030 -267.560 94.360 ;
        RECT -257.980 94.030 -257.640 94.360 ;
        RECT -248.060 94.030 -247.720 94.360 ;
        RECT -238.140 94.030 -237.800 94.360 ;
        RECT -228.220 94.030 -227.880 94.360 ;
        RECT -218.300 94.030 -217.960 94.360 ;
        RECT -208.380 94.030 -208.040 94.360 ;
        RECT -198.460 94.030 -198.120 94.360 ;
        RECT -188.540 94.030 -188.200 94.360 ;
        RECT -178.620 94.030 -178.280 94.360 ;
        RECT -168.700 94.030 -168.360 94.360 ;
        RECT -158.780 94.030 -158.440 94.360 ;
        RECT -148.860 94.030 -148.520 94.360 ;
        RECT -138.940 94.030 -138.600 94.360 ;
        RECT -129.020 94.030 -128.680 94.360 ;
        RECT -119.100 94.030 -118.760 94.360 ;
        RECT -109.180 94.030 -108.840 94.360 ;
        RECT -99.260 94.030 -98.920 94.360 ;
        RECT -89.340 94.030 -89.000 94.360 ;
        RECT -79.420 94.030 -79.080 94.360 ;
        RECT -69.500 94.030 -69.160 94.360 ;
        RECT -59.580 94.030 -59.240 94.360 ;
        RECT -49.660 94.030 -49.320 94.360 ;
        RECT -39.740 94.030 -39.400 94.360 ;
        RECT -29.820 94.030 -29.480 94.360 ;
        RECT -19.900 94.030 -19.560 94.360 ;
        RECT -9.980 94.030 -9.640 94.360 ;
        RECT -0.060 94.030 0.280 94.360 ;
        RECT 9.860 94.030 10.200 94.360 ;
        RECT 19.780 94.030 20.120 94.360 ;
        RECT -280.560 93.160 -280.220 93.490 ;
        RECT -280.090 93.160 -279.750 93.490 ;
        RECT -270.640 93.160 -270.300 93.490 ;
        RECT -270.170 93.160 -269.830 93.490 ;
        RECT -260.720 93.160 -260.380 93.490 ;
        RECT -260.250 93.160 -259.910 93.490 ;
        RECT -250.800 93.160 -250.460 93.490 ;
        RECT -250.330 93.160 -249.990 93.490 ;
        RECT -240.880 93.160 -240.540 93.490 ;
        RECT -240.410 93.160 -240.070 93.490 ;
        RECT -230.960 93.160 -230.620 93.490 ;
        RECT -230.490 93.160 -230.150 93.490 ;
        RECT -221.040 93.160 -220.700 93.490 ;
        RECT -220.570 93.160 -220.230 93.490 ;
        RECT -211.120 93.160 -210.780 93.490 ;
        RECT -210.650 93.160 -210.310 93.490 ;
        RECT -201.200 93.160 -200.860 93.490 ;
        RECT -200.730 93.160 -200.390 93.490 ;
        RECT -191.280 93.160 -190.940 93.490 ;
        RECT -190.810 93.160 -190.470 93.490 ;
        RECT -181.360 93.160 -181.020 93.490 ;
        RECT -180.890 93.160 -180.550 93.490 ;
        RECT -171.440 93.160 -171.100 93.490 ;
        RECT -170.970 93.160 -170.630 93.490 ;
        RECT -161.520 93.160 -161.180 93.490 ;
        RECT -161.050 93.160 -160.710 93.490 ;
        RECT -151.600 93.160 -151.260 93.490 ;
        RECT -151.130 93.160 -150.790 93.490 ;
        RECT -141.680 93.160 -141.340 93.490 ;
        RECT -141.210 93.160 -140.870 93.490 ;
        RECT -131.760 93.160 -131.420 93.490 ;
        RECT -131.290 93.160 -130.950 93.490 ;
        RECT -121.840 93.160 -121.500 93.490 ;
        RECT -121.370 93.160 -121.030 93.490 ;
        RECT -111.920 93.160 -111.580 93.490 ;
        RECT -111.450 93.160 -111.110 93.490 ;
        RECT -102.000 93.160 -101.660 93.490 ;
        RECT -101.530 93.160 -101.190 93.490 ;
        RECT -92.080 93.160 -91.740 93.490 ;
        RECT -91.610 93.160 -91.270 93.490 ;
        RECT -82.160 93.160 -81.820 93.490 ;
        RECT -81.690 93.160 -81.350 93.490 ;
        RECT -72.240 93.160 -71.900 93.490 ;
        RECT -71.770 93.160 -71.430 93.490 ;
        RECT -62.320 93.160 -61.980 93.490 ;
        RECT -61.850 93.160 -61.510 93.490 ;
        RECT -52.400 93.160 -52.060 93.490 ;
        RECT -51.930 93.160 -51.590 93.490 ;
        RECT -42.480 93.160 -42.140 93.490 ;
        RECT -42.010 93.160 -41.670 93.490 ;
        RECT -32.560 93.160 -32.220 93.490 ;
        RECT -32.090 93.160 -31.750 93.490 ;
        RECT -22.640 93.160 -22.300 93.490 ;
        RECT -22.170 93.160 -21.830 93.490 ;
        RECT -12.720 93.160 -12.380 93.490 ;
        RECT -12.250 93.160 -11.910 93.490 ;
        RECT -2.800 93.160 -2.460 93.490 ;
        RECT -2.330 93.160 -1.990 93.490 ;
        RECT 7.120 93.160 7.460 93.490 ;
        RECT 7.590 93.160 7.930 93.490 ;
        RECT 17.040 93.160 17.380 93.490 ;
        RECT 17.510 93.160 17.850 93.490 ;
        RECT -287.820 90.440 -287.480 90.770 ;
        RECT -287.360 90.440 -287.020 90.770 ;
        RECT -277.900 90.440 -277.560 90.770 ;
        RECT -277.440 90.440 -277.100 90.770 ;
        RECT -267.980 90.440 -267.640 90.770 ;
        RECT -267.520 90.440 -267.180 90.770 ;
        RECT -258.060 90.440 -257.720 90.770 ;
        RECT -257.600 90.440 -257.260 90.770 ;
        RECT -248.140 90.440 -247.800 90.770 ;
        RECT -247.680 90.440 -247.340 90.770 ;
        RECT -238.220 90.440 -237.880 90.770 ;
        RECT -237.760 90.440 -237.420 90.770 ;
        RECT -228.300 90.440 -227.960 90.770 ;
        RECT -227.840 90.440 -227.500 90.770 ;
        RECT -218.380 90.440 -218.040 90.770 ;
        RECT -217.920 90.440 -217.580 90.770 ;
        RECT -208.460 90.440 -208.120 90.770 ;
        RECT -208.000 90.440 -207.660 90.770 ;
        RECT -198.540 90.440 -198.200 90.770 ;
        RECT -198.080 90.440 -197.740 90.770 ;
        RECT -188.620 90.440 -188.280 90.770 ;
        RECT -188.160 90.440 -187.820 90.770 ;
        RECT -178.700 90.440 -178.360 90.770 ;
        RECT -178.240 90.440 -177.900 90.770 ;
        RECT -168.780 90.440 -168.440 90.770 ;
        RECT -168.320 90.440 -167.980 90.770 ;
        RECT -158.860 90.440 -158.520 90.770 ;
        RECT -158.400 90.440 -158.060 90.770 ;
        RECT -148.940 90.440 -148.600 90.770 ;
        RECT -148.480 90.440 -148.140 90.770 ;
        RECT -139.020 90.440 -138.680 90.770 ;
        RECT -138.560 90.440 -138.220 90.770 ;
        RECT -129.100 90.440 -128.760 90.770 ;
        RECT -128.640 90.440 -128.300 90.770 ;
        RECT -119.180 90.440 -118.840 90.770 ;
        RECT -118.720 90.440 -118.380 90.770 ;
        RECT -109.260 90.440 -108.920 90.770 ;
        RECT -108.800 90.440 -108.460 90.770 ;
        RECT -99.340 90.440 -99.000 90.770 ;
        RECT -98.880 90.440 -98.540 90.770 ;
        RECT -89.420 90.440 -89.080 90.770 ;
        RECT -88.960 90.440 -88.620 90.770 ;
        RECT -79.500 90.440 -79.160 90.770 ;
        RECT -79.040 90.440 -78.700 90.770 ;
        RECT -69.580 90.440 -69.240 90.770 ;
        RECT -69.120 90.440 -68.780 90.770 ;
        RECT -59.660 90.440 -59.320 90.770 ;
        RECT -59.200 90.440 -58.860 90.770 ;
        RECT -49.740 90.440 -49.400 90.770 ;
        RECT -49.280 90.440 -48.940 90.770 ;
        RECT -39.820 90.440 -39.480 90.770 ;
        RECT -39.360 90.440 -39.020 90.770 ;
        RECT -29.900 90.440 -29.560 90.770 ;
        RECT -29.440 90.440 -29.100 90.770 ;
        RECT -19.980 90.440 -19.640 90.770 ;
        RECT -19.520 90.440 -19.180 90.770 ;
        RECT -10.060 90.440 -9.720 90.770 ;
        RECT -9.600 90.440 -9.260 90.770 ;
        RECT -0.140 90.440 0.200 90.770 ;
        RECT 0.320 90.440 0.660 90.770 ;
        RECT 9.780 90.440 10.120 90.770 ;
        RECT 10.240 90.440 10.580 90.770 ;
        RECT 19.700 90.440 20.040 90.770 ;
        RECT 20.160 90.440 20.500 90.770 ;
        RECT -280.170 89.680 -279.830 90.010 ;
        RECT -270.250 89.680 -269.910 90.010 ;
        RECT -260.330 89.680 -259.990 90.010 ;
        RECT -250.410 89.680 -250.070 90.010 ;
        RECT -240.490 89.680 -240.150 90.010 ;
        RECT -230.570 89.680 -230.230 90.010 ;
        RECT -220.650 89.680 -220.310 90.010 ;
        RECT -210.730 89.680 -210.390 90.010 ;
        RECT -200.810 89.680 -200.470 90.010 ;
        RECT -190.890 89.680 -190.550 90.010 ;
        RECT -180.970 89.680 -180.630 90.010 ;
        RECT -171.050 89.680 -170.710 90.010 ;
        RECT -161.130 89.680 -160.790 90.010 ;
        RECT -151.210 89.680 -150.870 90.010 ;
        RECT -141.290 89.680 -140.950 90.010 ;
        RECT -131.370 89.680 -131.030 90.010 ;
        RECT -121.450 89.680 -121.110 90.010 ;
        RECT -111.530 89.680 -111.190 90.010 ;
        RECT -101.610 89.680 -101.270 90.010 ;
        RECT -91.690 89.680 -91.350 90.010 ;
        RECT -81.770 89.680 -81.430 90.010 ;
        RECT -71.850 89.680 -71.510 90.010 ;
        RECT -61.930 89.680 -61.590 90.010 ;
        RECT -52.010 89.680 -51.670 90.010 ;
        RECT -42.090 89.680 -41.750 90.010 ;
        RECT -32.170 89.680 -31.830 90.010 ;
        RECT -22.250 89.680 -21.910 90.010 ;
        RECT -12.330 89.680 -11.990 90.010 ;
        RECT -2.410 89.680 -2.070 90.010 ;
        RECT 7.510 89.680 7.850 90.010 ;
        RECT 17.430 89.680 17.770 90.010 ;
      LAYER met4 ;
        RECT 68.120 94.560 119.650 94.590 ;
        RECT -301.240 90.960 119.650 94.560 ;
        RECT -310.220 89.420 119.650 90.960 ;
        RECT -310.220 89.390 72.030 89.420 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -283.195 93.570 -279.425 95.330 ;
        RECT -273.275 93.570 -269.505 95.330 ;
        RECT -263.355 93.570 -259.585 95.330 ;
        RECT -253.435 93.570 -249.665 95.330 ;
        RECT -243.515 93.570 -239.745 95.330 ;
        RECT -233.595 93.570 -229.825 95.330 ;
        RECT -223.675 93.570 -219.905 95.330 ;
        RECT -213.755 93.570 -209.985 95.330 ;
        RECT -203.835 93.570 -200.065 95.330 ;
        RECT -193.915 93.570 -190.145 95.330 ;
        RECT -183.995 93.570 -180.225 95.330 ;
        RECT -174.075 93.570 -170.305 95.330 ;
        RECT -164.155 93.570 -160.385 95.330 ;
        RECT -154.235 93.570 -150.465 95.330 ;
        RECT -144.315 93.570 -140.545 95.330 ;
        RECT -134.395 93.570 -130.625 95.330 ;
        RECT -124.475 93.570 -120.705 95.330 ;
        RECT -114.555 93.570 -110.785 95.330 ;
        RECT -104.635 93.570 -100.865 95.330 ;
        RECT -94.715 93.570 -90.945 95.330 ;
        RECT -84.795 93.570 -81.025 95.330 ;
        RECT -74.875 93.570 -71.105 95.330 ;
        RECT -64.955 93.570 -61.185 95.330 ;
        RECT -55.035 93.570 -51.265 95.330 ;
        RECT -45.115 93.570 -41.345 95.330 ;
        RECT -35.195 93.570 -31.425 95.330 ;
        RECT -25.275 93.570 -21.505 95.330 ;
        RECT -15.355 93.570 -11.585 95.330 ;
        RECT -5.435 93.570 -1.665 95.330 ;
        RECT 4.485 93.570 8.255 95.330 ;
        RECT 14.405 93.570 18.175 95.330 ;
        RECT 24.325 95.095 25.930 95.330 ;
        RECT 24.325 95.090 26.440 95.095 ;
        RECT 24.325 93.570 26.630 95.090 ;
        RECT -281.730 93.520 -280.890 93.570 ;
        RECT -288.070 91.915 -284.470 93.520 ;
        RECT -283.110 90.420 -279.510 92.025 ;
        RECT -278.150 91.915 -274.550 93.520 ;
        RECT -271.810 93.510 -270.970 93.570 ;
        RECT -261.890 93.520 -261.050 93.570 ;
        RECT -273.190 90.420 -269.590 92.025 ;
        RECT -268.230 91.915 -264.630 93.520 ;
        RECT -263.270 90.420 -259.670 92.025 ;
        RECT -258.310 91.915 -254.710 93.520 ;
        RECT -251.970 93.510 -251.130 93.570 ;
        RECT -242.050 93.520 -241.210 93.570 ;
        RECT -253.350 90.420 -249.750 92.025 ;
        RECT -248.390 91.915 -244.790 93.520 ;
        RECT -243.430 90.420 -239.830 92.025 ;
        RECT -238.470 91.915 -234.870 93.520 ;
        RECT -232.130 93.510 -231.290 93.570 ;
        RECT -222.210 93.520 -221.370 93.570 ;
        RECT -233.510 90.420 -229.910 92.025 ;
        RECT -228.550 91.915 -224.950 93.520 ;
        RECT -223.590 90.420 -219.990 92.025 ;
        RECT -218.630 91.915 -215.030 93.520 ;
        RECT -212.290 93.510 -211.450 93.570 ;
        RECT -202.370 93.520 -201.530 93.570 ;
        RECT -213.670 90.420 -210.070 92.025 ;
        RECT -208.710 91.915 -205.110 93.520 ;
        RECT -203.750 90.420 -200.150 92.025 ;
        RECT -198.790 91.915 -195.190 93.520 ;
        RECT -192.450 93.510 -191.610 93.570 ;
        RECT -182.530 93.520 -181.690 93.570 ;
        RECT -193.830 90.420 -190.230 92.025 ;
        RECT -188.870 91.915 -185.270 93.520 ;
        RECT -183.910 90.420 -180.310 92.025 ;
        RECT -178.950 91.915 -175.350 93.520 ;
        RECT -172.610 93.510 -171.770 93.570 ;
        RECT -162.690 93.520 -161.850 93.570 ;
        RECT -173.990 90.420 -170.390 92.025 ;
        RECT -169.030 91.915 -165.430 93.520 ;
        RECT -164.070 90.420 -160.470 92.025 ;
        RECT -159.110 91.915 -155.510 93.520 ;
        RECT -152.770 93.510 -151.930 93.570 ;
        RECT -142.850 93.520 -142.010 93.570 ;
        RECT -154.150 90.420 -150.550 92.025 ;
        RECT -149.190 91.915 -145.590 93.520 ;
        RECT -144.230 90.420 -140.630 92.025 ;
        RECT -139.270 91.915 -135.670 93.520 ;
        RECT -132.930 93.510 -132.090 93.570 ;
        RECT -123.010 93.520 -122.170 93.570 ;
        RECT -134.310 90.420 -130.710 92.025 ;
        RECT -129.350 91.915 -125.750 93.520 ;
        RECT -124.390 90.420 -120.790 92.025 ;
        RECT -119.430 91.915 -115.830 93.520 ;
        RECT -113.090 93.510 -112.250 93.570 ;
        RECT -103.170 93.520 -102.330 93.570 ;
        RECT -114.470 90.420 -110.870 92.025 ;
        RECT -109.510 91.915 -105.910 93.520 ;
        RECT -104.550 90.420 -100.950 92.025 ;
        RECT -99.590 91.915 -95.990 93.520 ;
        RECT -93.250 93.510 -92.410 93.570 ;
        RECT -83.330 93.520 -82.490 93.570 ;
        RECT -94.630 90.420 -91.030 92.025 ;
        RECT -89.670 91.915 -86.070 93.520 ;
        RECT -84.710 90.420 -81.110 92.025 ;
        RECT -79.750 91.915 -76.150 93.520 ;
        RECT -73.410 93.510 -72.570 93.570 ;
        RECT -63.490 93.520 -62.650 93.570 ;
        RECT -74.790 90.420 -71.190 92.025 ;
        RECT -69.830 91.915 -66.230 93.520 ;
        RECT -64.870 90.420 -61.270 92.025 ;
        RECT -59.910 91.915 -56.310 93.520 ;
        RECT -53.570 93.510 -52.730 93.570 ;
        RECT -43.650 93.520 -42.810 93.570 ;
        RECT -54.950 90.420 -51.350 92.025 ;
        RECT -49.990 91.915 -46.390 93.520 ;
        RECT -45.030 90.420 -41.430 92.025 ;
        RECT -40.070 91.915 -36.470 93.520 ;
        RECT -33.730 93.510 -32.890 93.570 ;
        RECT -23.810 93.520 -22.970 93.570 ;
        RECT -35.110 90.420 -31.510 92.025 ;
        RECT -30.150 91.915 -26.550 93.520 ;
        RECT -25.190 90.420 -21.590 92.025 ;
        RECT -20.230 91.915 -16.630 93.520 ;
        RECT -13.890 93.510 -13.050 93.570 ;
        RECT -3.970 93.520 -3.130 93.570 ;
        RECT -15.270 90.420 -11.670 92.025 ;
        RECT -10.310 91.915 -6.710 93.520 ;
        RECT -5.350 90.420 -1.750 92.025 ;
        RECT -0.390 91.915 3.210 93.520 ;
        RECT 5.950 93.510 6.790 93.570 ;
        RECT 15.870 93.520 16.710 93.570 ;
        RECT 25.790 93.520 26.630 93.570 ;
        RECT 4.570 90.420 8.170 92.025 ;
        RECT 9.530 91.915 13.130 93.520 ;
        RECT 14.490 90.420 18.090 92.025 ;
        RECT 19.450 91.915 23.050 93.520 ;
        RECT 24.410 90.420 26.630 92.025 ;
        RECT -288.155 88.610 -284.385 90.370 ;
        RECT -278.235 88.610 -274.465 90.370 ;
        RECT -268.315 88.610 -264.545 90.370 ;
        RECT -258.395 88.610 -254.625 90.370 ;
        RECT -248.475 88.610 -244.705 90.370 ;
        RECT -238.555 88.610 -234.785 90.370 ;
        RECT -228.635 88.610 -224.865 90.370 ;
        RECT -218.715 88.610 -214.945 90.370 ;
        RECT -208.795 88.610 -205.025 90.370 ;
        RECT -198.875 88.610 -195.105 90.370 ;
        RECT -188.955 88.610 -185.185 90.370 ;
        RECT -179.035 88.610 -175.265 90.370 ;
        RECT -169.115 88.610 -165.345 90.370 ;
        RECT -159.195 88.610 -155.425 90.370 ;
        RECT -149.275 88.610 -145.505 90.370 ;
        RECT -139.355 88.610 -135.585 90.370 ;
        RECT -129.435 88.610 -125.665 90.370 ;
        RECT -119.515 88.610 -115.745 90.370 ;
        RECT -109.595 88.610 -105.825 90.370 ;
        RECT -99.675 88.610 -95.905 90.370 ;
        RECT -89.755 88.610 -85.985 90.370 ;
        RECT -79.835 88.610 -76.065 90.370 ;
        RECT -69.915 88.610 -66.145 90.370 ;
        RECT -59.995 88.610 -56.225 90.370 ;
        RECT -50.075 88.610 -46.305 90.370 ;
        RECT -40.155 88.610 -36.385 90.370 ;
        RECT -30.235 88.610 -26.465 90.370 ;
        RECT -20.315 88.610 -16.545 90.370 ;
        RECT -10.395 88.610 -6.625 90.370 ;
        RECT -0.475 88.610 3.295 90.370 ;
        RECT 9.445 88.610 13.215 90.370 ;
        RECT 19.365 88.610 23.135 90.370 ;
      LAYER li1 ;
        RECT -281.865 94.990 -281.695 95.140 ;
        RECT -280.925 94.990 -280.755 95.140 ;
        RECT -281.865 94.820 -280.755 94.990 ;
        RECT -281.865 94.615 -281.695 94.820 ;
        RECT -282.625 94.285 -281.695 94.615 ;
        RECT -281.865 93.760 -281.695 94.285 ;
        RECT -281.455 93.655 -281.165 94.820 ;
        RECT -280.925 94.615 -280.755 94.820 ;
        RECT -271.945 94.990 -271.775 95.140 ;
        RECT -271.005 94.990 -270.835 95.140 ;
        RECT -271.945 94.820 -270.835 94.990 ;
        RECT -271.945 94.615 -271.775 94.820 ;
        RECT -280.925 94.285 -279.995 94.615 ;
        RECT -272.705 94.285 -271.775 94.615 ;
        RECT -280.925 93.760 -280.755 94.285 ;
        RECT -271.945 93.760 -271.775 94.285 ;
        RECT -271.535 93.655 -271.245 94.820 ;
        RECT -271.005 94.615 -270.835 94.820 ;
        RECT -262.025 94.990 -261.855 95.140 ;
        RECT -261.085 94.990 -260.915 95.140 ;
        RECT -262.025 94.820 -260.915 94.990 ;
        RECT -262.025 94.615 -261.855 94.820 ;
        RECT -271.005 94.285 -270.075 94.615 ;
        RECT -262.785 94.285 -261.855 94.615 ;
        RECT -271.005 93.760 -270.835 94.285 ;
        RECT -262.025 93.760 -261.855 94.285 ;
        RECT -261.615 93.655 -261.325 94.820 ;
        RECT -261.085 94.615 -260.915 94.820 ;
        RECT -252.105 94.990 -251.935 95.140 ;
        RECT -251.165 94.990 -250.995 95.140 ;
        RECT -252.105 94.820 -250.995 94.990 ;
        RECT -252.105 94.615 -251.935 94.820 ;
        RECT -261.085 94.285 -260.155 94.615 ;
        RECT -252.865 94.285 -251.935 94.615 ;
        RECT -261.085 93.760 -260.915 94.285 ;
        RECT -252.105 93.760 -251.935 94.285 ;
        RECT -251.695 93.655 -251.405 94.820 ;
        RECT -251.165 94.615 -250.995 94.820 ;
        RECT -242.185 94.990 -242.015 95.140 ;
        RECT -241.245 94.990 -241.075 95.140 ;
        RECT -242.185 94.820 -241.075 94.990 ;
        RECT -242.185 94.615 -242.015 94.820 ;
        RECT -251.165 94.285 -250.235 94.615 ;
        RECT -242.945 94.285 -242.015 94.615 ;
        RECT -251.165 93.760 -250.995 94.285 ;
        RECT -242.185 93.760 -242.015 94.285 ;
        RECT -241.775 93.655 -241.485 94.820 ;
        RECT -241.245 94.615 -241.075 94.820 ;
        RECT -232.265 94.990 -232.095 95.140 ;
        RECT -231.325 94.990 -231.155 95.140 ;
        RECT -232.265 94.820 -231.155 94.990 ;
        RECT -232.265 94.615 -232.095 94.820 ;
        RECT -241.245 94.285 -240.315 94.615 ;
        RECT -233.025 94.285 -232.095 94.615 ;
        RECT -241.245 93.760 -241.075 94.285 ;
        RECT -232.265 93.760 -232.095 94.285 ;
        RECT -231.855 93.655 -231.565 94.820 ;
        RECT -231.325 94.615 -231.155 94.820 ;
        RECT -222.345 94.990 -222.175 95.140 ;
        RECT -221.405 94.990 -221.235 95.140 ;
        RECT -222.345 94.820 -221.235 94.990 ;
        RECT -222.345 94.615 -222.175 94.820 ;
        RECT -231.325 94.285 -230.395 94.615 ;
        RECT -223.105 94.285 -222.175 94.615 ;
        RECT -231.325 93.760 -231.155 94.285 ;
        RECT -222.345 93.760 -222.175 94.285 ;
        RECT -221.935 93.655 -221.645 94.820 ;
        RECT -221.405 94.615 -221.235 94.820 ;
        RECT -212.425 94.990 -212.255 95.140 ;
        RECT -211.485 94.990 -211.315 95.140 ;
        RECT -212.425 94.820 -211.315 94.990 ;
        RECT -212.425 94.615 -212.255 94.820 ;
        RECT -221.405 94.285 -220.475 94.615 ;
        RECT -213.185 94.285 -212.255 94.615 ;
        RECT -221.405 93.760 -221.235 94.285 ;
        RECT -212.425 93.760 -212.255 94.285 ;
        RECT -212.015 93.655 -211.725 94.820 ;
        RECT -211.485 94.615 -211.315 94.820 ;
        RECT -202.505 94.990 -202.335 95.140 ;
        RECT -201.565 94.990 -201.395 95.140 ;
        RECT -202.505 94.820 -201.395 94.990 ;
        RECT -202.505 94.615 -202.335 94.820 ;
        RECT -211.485 94.285 -210.555 94.615 ;
        RECT -203.265 94.285 -202.335 94.615 ;
        RECT -211.485 93.760 -211.315 94.285 ;
        RECT -202.505 93.760 -202.335 94.285 ;
        RECT -202.095 93.655 -201.805 94.820 ;
        RECT -201.565 94.615 -201.395 94.820 ;
        RECT -192.585 94.990 -192.415 95.140 ;
        RECT -191.645 94.990 -191.475 95.140 ;
        RECT -192.585 94.820 -191.475 94.990 ;
        RECT -192.585 94.615 -192.415 94.820 ;
        RECT -201.565 94.285 -200.635 94.615 ;
        RECT -193.345 94.285 -192.415 94.615 ;
        RECT -201.565 93.760 -201.395 94.285 ;
        RECT -192.585 93.760 -192.415 94.285 ;
        RECT -192.175 93.655 -191.885 94.820 ;
        RECT -191.645 94.615 -191.475 94.820 ;
        RECT -182.665 94.990 -182.495 95.140 ;
        RECT -181.725 94.990 -181.555 95.140 ;
        RECT -182.665 94.820 -181.555 94.990 ;
        RECT -182.665 94.615 -182.495 94.820 ;
        RECT -191.645 94.285 -190.715 94.615 ;
        RECT -183.425 94.285 -182.495 94.615 ;
        RECT -191.645 93.760 -191.475 94.285 ;
        RECT -182.665 93.760 -182.495 94.285 ;
        RECT -182.255 93.655 -181.965 94.820 ;
        RECT -181.725 94.615 -181.555 94.820 ;
        RECT -172.745 94.990 -172.575 95.140 ;
        RECT -171.805 94.990 -171.635 95.140 ;
        RECT -172.745 94.820 -171.635 94.990 ;
        RECT -172.745 94.615 -172.575 94.820 ;
        RECT -181.725 94.285 -180.795 94.615 ;
        RECT -173.505 94.285 -172.575 94.615 ;
        RECT -181.725 93.760 -181.555 94.285 ;
        RECT -172.745 93.760 -172.575 94.285 ;
        RECT -172.335 93.655 -172.045 94.820 ;
        RECT -171.805 94.615 -171.635 94.820 ;
        RECT -162.825 94.990 -162.655 95.140 ;
        RECT -161.885 94.990 -161.715 95.140 ;
        RECT -162.825 94.820 -161.715 94.990 ;
        RECT -162.825 94.615 -162.655 94.820 ;
        RECT -171.805 94.285 -170.875 94.615 ;
        RECT -163.585 94.285 -162.655 94.615 ;
        RECT -171.805 93.760 -171.635 94.285 ;
        RECT -162.825 93.760 -162.655 94.285 ;
        RECT -162.415 93.655 -162.125 94.820 ;
        RECT -161.885 94.615 -161.715 94.820 ;
        RECT -152.905 94.990 -152.735 95.140 ;
        RECT -151.965 94.990 -151.795 95.140 ;
        RECT -152.905 94.820 -151.795 94.990 ;
        RECT -152.905 94.615 -152.735 94.820 ;
        RECT -161.885 94.285 -160.955 94.615 ;
        RECT -153.665 94.285 -152.735 94.615 ;
        RECT -161.885 93.760 -161.715 94.285 ;
        RECT -152.905 93.760 -152.735 94.285 ;
        RECT -152.495 93.655 -152.205 94.820 ;
        RECT -151.965 94.615 -151.795 94.820 ;
        RECT -142.985 94.990 -142.815 95.140 ;
        RECT -142.045 94.990 -141.875 95.140 ;
        RECT -142.985 94.820 -141.875 94.990 ;
        RECT -142.985 94.615 -142.815 94.820 ;
        RECT -151.965 94.285 -151.035 94.615 ;
        RECT -143.745 94.285 -142.815 94.615 ;
        RECT -151.965 93.760 -151.795 94.285 ;
        RECT -142.985 93.760 -142.815 94.285 ;
        RECT -142.575 93.655 -142.285 94.820 ;
        RECT -142.045 94.615 -141.875 94.820 ;
        RECT -133.065 94.990 -132.895 95.140 ;
        RECT -132.125 94.990 -131.955 95.140 ;
        RECT -133.065 94.820 -131.955 94.990 ;
        RECT -133.065 94.615 -132.895 94.820 ;
        RECT -142.045 94.285 -141.115 94.615 ;
        RECT -133.825 94.285 -132.895 94.615 ;
        RECT -142.045 93.760 -141.875 94.285 ;
        RECT -133.065 93.760 -132.895 94.285 ;
        RECT -132.655 93.655 -132.365 94.820 ;
        RECT -132.125 94.615 -131.955 94.820 ;
        RECT -123.145 94.990 -122.975 95.140 ;
        RECT -122.205 94.990 -122.035 95.140 ;
        RECT -123.145 94.820 -122.035 94.990 ;
        RECT -123.145 94.615 -122.975 94.820 ;
        RECT -132.125 94.285 -131.195 94.615 ;
        RECT -123.905 94.285 -122.975 94.615 ;
        RECT -132.125 93.760 -131.955 94.285 ;
        RECT -123.145 93.760 -122.975 94.285 ;
        RECT -122.735 93.655 -122.445 94.820 ;
        RECT -122.205 94.615 -122.035 94.820 ;
        RECT -113.225 94.990 -113.055 95.140 ;
        RECT -112.285 94.990 -112.115 95.140 ;
        RECT -113.225 94.820 -112.115 94.990 ;
        RECT -113.225 94.615 -113.055 94.820 ;
        RECT -122.205 94.285 -121.275 94.615 ;
        RECT -113.985 94.285 -113.055 94.615 ;
        RECT -122.205 93.760 -122.035 94.285 ;
        RECT -113.225 93.760 -113.055 94.285 ;
        RECT -112.815 93.655 -112.525 94.820 ;
        RECT -112.285 94.615 -112.115 94.820 ;
        RECT -103.305 94.990 -103.135 95.140 ;
        RECT -102.365 94.990 -102.195 95.140 ;
        RECT -103.305 94.820 -102.195 94.990 ;
        RECT -103.305 94.615 -103.135 94.820 ;
        RECT -112.285 94.285 -111.355 94.615 ;
        RECT -104.065 94.285 -103.135 94.615 ;
        RECT -112.285 93.760 -112.115 94.285 ;
        RECT -103.305 93.760 -103.135 94.285 ;
        RECT -102.895 93.655 -102.605 94.820 ;
        RECT -102.365 94.615 -102.195 94.820 ;
        RECT -93.385 94.990 -93.215 95.140 ;
        RECT -92.445 94.990 -92.275 95.140 ;
        RECT -93.385 94.820 -92.275 94.990 ;
        RECT -93.385 94.615 -93.215 94.820 ;
        RECT -102.365 94.285 -101.435 94.615 ;
        RECT -94.145 94.285 -93.215 94.615 ;
        RECT -102.365 93.760 -102.195 94.285 ;
        RECT -93.385 93.760 -93.215 94.285 ;
        RECT -92.975 93.655 -92.685 94.820 ;
        RECT -92.445 94.615 -92.275 94.820 ;
        RECT -83.465 94.990 -83.295 95.140 ;
        RECT -82.525 94.990 -82.355 95.140 ;
        RECT -83.465 94.820 -82.355 94.990 ;
        RECT -83.465 94.615 -83.295 94.820 ;
        RECT -92.445 94.285 -91.515 94.615 ;
        RECT -84.225 94.285 -83.295 94.615 ;
        RECT -92.445 93.760 -92.275 94.285 ;
        RECT -83.465 93.760 -83.295 94.285 ;
        RECT -83.055 93.655 -82.765 94.820 ;
        RECT -82.525 94.615 -82.355 94.820 ;
        RECT -73.545 94.990 -73.375 95.140 ;
        RECT -72.605 94.990 -72.435 95.140 ;
        RECT -73.545 94.820 -72.435 94.990 ;
        RECT -73.545 94.615 -73.375 94.820 ;
        RECT -82.525 94.285 -81.595 94.615 ;
        RECT -74.305 94.285 -73.375 94.615 ;
        RECT -82.525 93.760 -82.355 94.285 ;
        RECT -73.545 93.760 -73.375 94.285 ;
        RECT -73.135 93.655 -72.845 94.820 ;
        RECT -72.605 94.615 -72.435 94.820 ;
        RECT -63.625 94.990 -63.455 95.140 ;
        RECT -62.685 94.990 -62.515 95.140 ;
        RECT -63.625 94.820 -62.515 94.990 ;
        RECT -63.625 94.615 -63.455 94.820 ;
        RECT -72.605 94.285 -71.675 94.615 ;
        RECT -64.385 94.285 -63.455 94.615 ;
        RECT -72.605 93.760 -72.435 94.285 ;
        RECT -63.625 93.760 -63.455 94.285 ;
        RECT -63.215 93.655 -62.925 94.820 ;
        RECT -62.685 94.615 -62.515 94.820 ;
        RECT -53.705 94.990 -53.535 95.140 ;
        RECT -52.765 94.990 -52.595 95.140 ;
        RECT -53.705 94.820 -52.595 94.990 ;
        RECT -53.705 94.615 -53.535 94.820 ;
        RECT -62.685 94.285 -61.755 94.615 ;
        RECT -54.465 94.285 -53.535 94.615 ;
        RECT -62.685 93.760 -62.515 94.285 ;
        RECT -53.705 93.760 -53.535 94.285 ;
        RECT -53.295 93.655 -53.005 94.820 ;
        RECT -52.765 94.615 -52.595 94.820 ;
        RECT -43.785 94.990 -43.615 95.140 ;
        RECT -42.845 94.990 -42.675 95.140 ;
        RECT -43.785 94.820 -42.675 94.990 ;
        RECT -43.785 94.615 -43.615 94.820 ;
        RECT -52.765 94.285 -51.835 94.615 ;
        RECT -44.545 94.285 -43.615 94.615 ;
        RECT -52.765 93.760 -52.595 94.285 ;
        RECT -43.785 93.760 -43.615 94.285 ;
        RECT -43.375 93.655 -43.085 94.820 ;
        RECT -42.845 94.615 -42.675 94.820 ;
        RECT -33.865 94.990 -33.695 95.140 ;
        RECT -32.925 94.990 -32.755 95.140 ;
        RECT -33.865 94.820 -32.755 94.990 ;
        RECT -33.865 94.615 -33.695 94.820 ;
        RECT -42.845 94.285 -41.915 94.615 ;
        RECT -34.625 94.285 -33.695 94.615 ;
        RECT -42.845 93.760 -42.675 94.285 ;
        RECT -33.865 93.760 -33.695 94.285 ;
        RECT -33.455 93.655 -33.165 94.820 ;
        RECT -32.925 94.615 -32.755 94.820 ;
        RECT -23.945 94.990 -23.775 95.140 ;
        RECT -23.005 94.990 -22.835 95.140 ;
        RECT -23.945 94.820 -22.835 94.990 ;
        RECT -23.945 94.615 -23.775 94.820 ;
        RECT -32.925 94.285 -31.995 94.615 ;
        RECT -24.705 94.285 -23.775 94.615 ;
        RECT -32.925 93.760 -32.755 94.285 ;
        RECT -23.945 93.760 -23.775 94.285 ;
        RECT -23.535 93.655 -23.245 94.820 ;
        RECT -23.005 94.615 -22.835 94.820 ;
        RECT -14.025 94.990 -13.855 95.140 ;
        RECT -13.085 94.990 -12.915 95.140 ;
        RECT -14.025 94.820 -12.915 94.990 ;
        RECT -14.025 94.615 -13.855 94.820 ;
        RECT -23.005 94.285 -22.075 94.615 ;
        RECT -14.785 94.285 -13.855 94.615 ;
        RECT -23.005 93.760 -22.835 94.285 ;
        RECT -14.025 93.760 -13.855 94.285 ;
        RECT -13.615 93.655 -13.325 94.820 ;
        RECT -13.085 94.615 -12.915 94.820 ;
        RECT -4.105 94.990 -3.935 95.140 ;
        RECT -3.165 94.990 -2.995 95.140 ;
        RECT -4.105 94.820 -2.995 94.990 ;
        RECT -4.105 94.615 -3.935 94.820 ;
        RECT -13.085 94.285 -12.155 94.615 ;
        RECT -4.865 94.285 -3.935 94.615 ;
        RECT -13.085 93.760 -12.915 94.285 ;
        RECT -4.105 93.760 -3.935 94.285 ;
        RECT -3.695 93.655 -3.405 94.820 ;
        RECT -3.165 94.615 -2.995 94.820 ;
        RECT 5.815 94.990 5.985 95.140 ;
        RECT 6.755 94.990 6.925 95.140 ;
        RECT 5.815 94.820 6.925 94.990 ;
        RECT 5.815 94.615 5.985 94.820 ;
        RECT -3.165 94.285 -2.235 94.615 ;
        RECT 5.055 94.285 5.985 94.615 ;
        RECT -3.165 93.760 -2.995 94.285 ;
        RECT 5.815 93.760 5.985 94.285 ;
        RECT 6.225 93.655 6.515 94.820 ;
        RECT 6.755 94.615 6.925 94.820 ;
        RECT 15.735 94.990 15.905 95.140 ;
        RECT 16.675 94.990 16.845 95.140 ;
        RECT 15.735 94.820 16.845 94.990 ;
        RECT 15.735 94.615 15.905 94.820 ;
        RECT 6.755 94.285 7.685 94.615 ;
        RECT 14.975 94.285 15.905 94.615 ;
        RECT 6.755 93.760 6.925 94.285 ;
        RECT 15.735 93.760 15.905 94.285 ;
        RECT 16.145 93.655 16.435 94.820 ;
        RECT 16.675 94.615 16.845 94.820 ;
        RECT 25.655 94.990 25.825 95.140 ;
        RECT 25.655 94.820 26.440 94.990 ;
        RECT 25.655 94.615 25.825 94.820 ;
        RECT 16.675 94.285 17.605 94.615 ;
        RECT 24.895 94.285 25.825 94.615 ;
        RECT 16.675 93.760 16.845 94.285 ;
        RECT 25.655 93.760 25.825 94.285 ;
        RECT 26.065 93.655 26.355 94.820 ;
        RECT -287.880 93.245 -284.660 93.415 ;
        RECT -277.960 93.245 -274.740 93.415 ;
        RECT -268.040 93.245 -264.820 93.415 ;
        RECT -258.120 93.245 -254.900 93.415 ;
        RECT -248.200 93.245 -244.980 93.415 ;
        RECT -238.280 93.245 -235.060 93.415 ;
        RECT -228.360 93.245 -225.140 93.415 ;
        RECT -218.440 93.245 -215.220 93.415 ;
        RECT -208.520 93.245 -205.300 93.415 ;
        RECT -198.600 93.245 -195.380 93.415 ;
        RECT -188.680 93.245 -185.460 93.415 ;
        RECT -178.760 93.245 -175.540 93.415 ;
        RECT -168.840 93.245 -165.620 93.415 ;
        RECT -158.920 93.245 -155.700 93.415 ;
        RECT -149.000 93.245 -145.780 93.415 ;
        RECT -139.080 93.245 -135.860 93.415 ;
        RECT -129.160 93.245 -125.940 93.415 ;
        RECT -119.240 93.245 -116.020 93.415 ;
        RECT -109.320 93.245 -106.100 93.415 ;
        RECT -99.400 93.245 -96.180 93.415 ;
        RECT -89.480 93.245 -86.260 93.415 ;
        RECT -79.560 93.245 -76.340 93.415 ;
        RECT -69.640 93.245 -66.420 93.415 ;
        RECT -59.720 93.245 -56.500 93.415 ;
        RECT -49.800 93.245 -46.580 93.415 ;
        RECT -39.880 93.245 -36.660 93.415 ;
        RECT -29.960 93.245 -26.740 93.415 ;
        RECT -20.040 93.245 -16.820 93.415 ;
        RECT -10.120 93.245 -6.900 93.415 ;
        RECT -0.200 93.245 3.020 93.415 ;
        RECT 9.720 93.245 12.940 93.415 ;
        RECT 19.640 93.245 22.860 93.415 ;
        RECT -287.795 92.105 -287.535 93.245 ;
        RECT -286.865 92.105 -286.585 93.245 ;
        RECT -286.415 92.080 -286.125 93.245 ;
        RECT -285.955 92.105 -285.675 93.245 ;
        RECT -285.005 92.105 -284.745 93.245 ;
        RECT -277.875 92.105 -277.615 93.245 ;
        RECT -276.945 92.105 -276.665 93.245 ;
        RECT -276.495 92.080 -276.205 93.245 ;
        RECT -276.035 92.105 -275.755 93.245 ;
        RECT -275.085 92.105 -274.825 93.245 ;
        RECT -267.955 92.105 -267.695 93.245 ;
        RECT -267.025 92.105 -266.745 93.245 ;
        RECT -266.575 92.080 -266.285 93.245 ;
        RECT -266.115 92.105 -265.835 93.245 ;
        RECT -265.165 92.105 -264.905 93.245 ;
        RECT -258.035 92.105 -257.775 93.245 ;
        RECT -257.105 92.105 -256.825 93.245 ;
        RECT -256.655 92.080 -256.365 93.245 ;
        RECT -256.195 92.105 -255.915 93.245 ;
        RECT -255.245 92.105 -254.985 93.245 ;
        RECT -248.115 92.105 -247.855 93.245 ;
        RECT -247.185 92.105 -246.905 93.245 ;
        RECT -246.735 92.080 -246.445 93.245 ;
        RECT -246.275 92.105 -245.995 93.245 ;
        RECT -245.325 92.105 -245.065 93.245 ;
        RECT -238.195 92.105 -237.935 93.245 ;
        RECT -237.265 92.105 -236.985 93.245 ;
        RECT -236.815 92.080 -236.525 93.245 ;
        RECT -236.355 92.105 -236.075 93.245 ;
        RECT -235.405 92.105 -235.145 93.245 ;
        RECT -228.275 92.105 -228.015 93.245 ;
        RECT -227.345 92.105 -227.065 93.245 ;
        RECT -226.895 92.080 -226.605 93.245 ;
        RECT -226.435 92.105 -226.155 93.245 ;
        RECT -225.485 92.105 -225.225 93.245 ;
        RECT -218.355 92.105 -218.095 93.245 ;
        RECT -217.425 92.105 -217.145 93.245 ;
        RECT -216.975 92.080 -216.685 93.245 ;
        RECT -216.515 92.105 -216.235 93.245 ;
        RECT -215.565 92.105 -215.305 93.245 ;
        RECT -208.435 92.105 -208.175 93.245 ;
        RECT -207.505 92.105 -207.225 93.245 ;
        RECT -207.055 92.080 -206.765 93.245 ;
        RECT -206.595 92.105 -206.315 93.245 ;
        RECT -205.645 92.105 -205.385 93.245 ;
        RECT -198.515 92.105 -198.255 93.245 ;
        RECT -197.585 92.105 -197.305 93.245 ;
        RECT -197.135 92.080 -196.845 93.245 ;
        RECT -196.675 92.105 -196.395 93.245 ;
        RECT -195.725 92.105 -195.465 93.245 ;
        RECT -188.595 92.105 -188.335 93.245 ;
        RECT -187.665 92.105 -187.385 93.245 ;
        RECT -187.215 92.080 -186.925 93.245 ;
        RECT -186.755 92.105 -186.475 93.245 ;
        RECT -185.805 92.105 -185.545 93.245 ;
        RECT -178.675 92.105 -178.415 93.245 ;
        RECT -177.745 92.105 -177.465 93.245 ;
        RECT -177.295 92.080 -177.005 93.245 ;
        RECT -176.835 92.105 -176.555 93.245 ;
        RECT -175.885 92.105 -175.625 93.245 ;
        RECT -168.755 92.105 -168.495 93.245 ;
        RECT -167.825 92.105 -167.545 93.245 ;
        RECT -167.375 92.080 -167.085 93.245 ;
        RECT -166.915 92.105 -166.635 93.245 ;
        RECT -165.965 92.105 -165.705 93.245 ;
        RECT -158.835 92.105 -158.575 93.245 ;
        RECT -157.905 92.105 -157.625 93.245 ;
        RECT -157.455 92.080 -157.165 93.245 ;
        RECT -156.995 92.105 -156.715 93.245 ;
        RECT -156.045 92.105 -155.785 93.245 ;
        RECT -148.915 92.105 -148.655 93.245 ;
        RECT -147.985 92.105 -147.705 93.245 ;
        RECT -147.535 92.080 -147.245 93.245 ;
        RECT -147.075 92.105 -146.795 93.245 ;
        RECT -146.125 92.105 -145.865 93.245 ;
        RECT -138.995 92.105 -138.735 93.245 ;
        RECT -138.065 92.105 -137.785 93.245 ;
        RECT -137.615 92.080 -137.325 93.245 ;
        RECT -137.155 92.105 -136.875 93.245 ;
        RECT -136.205 92.105 -135.945 93.245 ;
        RECT -129.075 92.105 -128.815 93.245 ;
        RECT -128.145 92.105 -127.865 93.245 ;
        RECT -127.695 92.080 -127.405 93.245 ;
        RECT -127.235 92.105 -126.955 93.245 ;
        RECT -126.285 92.105 -126.025 93.245 ;
        RECT -119.155 92.105 -118.895 93.245 ;
        RECT -118.225 92.105 -117.945 93.245 ;
        RECT -117.775 92.080 -117.485 93.245 ;
        RECT -117.315 92.105 -117.035 93.245 ;
        RECT -116.365 92.105 -116.105 93.245 ;
        RECT -109.235 92.105 -108.975 93.245 ;
        RECT -108.305 92.105 -108.025 93.245 ;
        RECT -107.855 92.080 -107.565 93.245 ;
        RECT -107.395 92.105 -107.115 93.245 ;
        RECT -106.445 92.105 -106.185 93.245 ;
        RECT -99.315 92.105 -99.055 93.245 ;
        RECT -98.385 92.105 -98.105 93.245 ;
        RECT -97.935 92.080 -97.645 93.245 ;
        RECT -97.475 92.105 -97.195 93.245 ;
        RECT -96.525 92.105 -96.265 93.245 ;
        RECT -89.395 92.105 -89.135 93.245 ;
        RECT -88.465 92.105 -88.185 93.245 ;
        RECT -88.015 92.080 -87.725 93.245 ;
        RECT -87.555 92.105 -87.275 93.245 ;
        RECT -86.605 92.105 -86.345 93.245 ;
        RECT -79.475 92.105 -79.215 93.245 ;
        RECT -78.545 92.105 -78.265 93.245 ;
        RECT -78.095 92.080 -77.805 93.245 ;
        RECT -77.635 92.105 -77.355 93.245 ;
        RECT -76.685 92.105 -76.425 93.245 ;
        RECT -69.555 92.105 -69.295 93.245 ;
        RECT -68.625 92.105 -68.345 93.245 ;
        RECT -68.175 92.080 -67.885 93.245 ;
        RECT -67.715 92.105 -67.435 93.245 ;
        RECT -66.765 92.105 -66.505 93.245 ;
        RECT -59.635 92.105 -59.375 93.245 ;
        RECT -58.705 92.105 -58.425 93.245 ;
        RECT -58.255 92.080 -57.965 93.245 ;
        RECT -57.795 92.105 -57.515 93.245 ;
        RECT -56.845 92.105 -56.585 93.245 ;
        RECT -49.715 92.105 -49.455 93.245 ;
        RECT -48.785 92.105 -48.505 93.245 ;
        RECT -48.335 92.080 -48.045 93.245 ;
        RECT -47.875 92.105 -47.595 93.245 ;
        RECT -46.925 92.105 -46.665 93.245 ;
        RECT -39.795 92.105 -39.535 93.245 ;
        RECT -38.865 92.105 -38.585 93.245 ;
        RECT -38.415 92.080 -38.125 93.245 ;
        RECT -37.955 92.105 -37.675 93.245 ;
        RECT -37.005 92.105 -36.745 93.245 ;
        RECT -29.875 92.105 -29.615 93.245 ;
        RECT -28.945 92.105 -28.665 93.245 ;
        RECT -28.495 92.080 -28.205 93.245 ;
        RECT -28.035 92.105 -27.755 93.245 ;
        RECT -27.085 92.105 -26.825 93.245 ;
        RECT -19.955 92.105 -19.695 93.245 ;
        RECT -19.025 92.105 -18.745 93.245 ;
        RECT -18.575 92.080 -18.285 93.245 ;
        RECT -18.115 92.105 -17.835 93.245 ;
        RECT -17.165 92.105 -16.905 93.245 ;
        RECT -10.035 92.105 -9.775 93.245 ;
        RECT -9.105 92.105 -8.825 93.245 ;
        RECT -8.655 92.080 -8.365 93.245 ;
        RECT -8.195 92.105 -7.915 93.245 ;
        RECT -7.245 92.105 -6.985 93.245 ;
        RECT -0.115 92.105 0.145 93.245 ;
        RECT 0.815 92.105 1.095 93.245 ;
        RECT 1.265 92.080 1.555 93.245 ;
        RECT 1.725 92.105 2.005 93.245 ;
        RECT 2.675 92.105 2.935 93.245 ;
        RECT 9.805 92.105 10.065 93.245 ;
        RECT 10.735 92.105 11.015 93.245 ;
        RECT 11.185 92.080 11.475 93.245 ;
        RECT 11.645 92.105 11.925 93.245 ;
        RECT 12.595 92.105 12.855 93.245 ;
        RECT 19.725 92.105 19.985 93.245 ;
        RECT 20.655 92.105 20.935 93.245 ;
        RECT 21.105 92.080 21.395 93.245 ;
        RECT 21.565 92.105 21.845 93.245 ;
        RECT 22.515 92.105 22.775 93.245 ;
        RECT -282.835 90.695 -282.575 91.835 ;
        RECT -281.905 90.695 -281.625 91.835 ;
        RECT -281.455 90.695 -281.165 91.860 ;
        RECT -280.995 90.695 -280.715 91.835 ;
        RECT -280.045 90.695 -279.785 91.835 ;
        RECT -272.915 90.695 -272.655 91.835 ;
        RECT -271.985 90.695 -271.705 91.835 ;
        RECT -271.535 90.695 -271.245 91.860 ;
        RECT -271.075 90.695 -270.795 91.835 ;
        RECT -270.125 90.695 -269.865 91.835 ;
        RECT -262.995 90.695 -262.735 91.835 ;
        RECT -262.065 90.695 -261.785 91.835 ;
        RECT -261.615 90.695 -261.325 91.860 ;
        RECT -261.155 90.695 -260.875 91.835 ;
        RECT -260.205 90.695 -259.945 91.835 ;
        RECT -253.075 90.695 -252.815 91.835 ;
        RECT -252.145 90.695 -251.865 91.835 ;
        RECT -251.695 90.695 -251.405 91.860 ;
        RECT -251.235 90.695 -250.955 91.835 ;
        RECT -250.285 90.695 -250.025 91.835 ;
        RECT -243.155 90.695 -242.895 91.835 ;
        RECT -242.225 90.695 -241.945 91.835 ;
        RECT -241.775 90.695 -241.485 91.860 ;
        RECT -241.315 90.695 -241.035 91.835 ;
        RECT -240.365 90.695 -240.105 91.835 ;
        RECT -233.235 90.695 -232.975 91.835 ;
        RECT -232.305 90.695 -232.025 91.835 ;
        RECT -231.855 90.695 -231.565 91.860 ;
        RECT -231.395 90.695 -231.115 91.835 ;
        RECT -230.445 90.695 -230.185 91.835 ;
        RECT -223.315 90.695 -223.055 91.835 ;
        RECT -222.385 90.695 -222.105 91.835 ;
        RECT -221.935 90.695 -221.645 91.860 ;
        RECT -221.475 90.695 -221.195 91.835 ;
        RECT -220.525 90.695 -220.265 91.835 ;
        RECT -213.395 90.695 -213.135 91.835 ;
        RECT -212.465 90.695 -212.185 91.835 ;
        RECT -212.015 90.695 -211.725 91.860 ;
        RECT -211.555 90.695 -211.275 91.835 ;
        RECT -210.605 90.695 -210.345 91.835 ;
        RECT -203.475 90.695 -203.215 91.835 ;
        RECT -202.545 90.695 -202.265 91.835 ;
        RECT -202.095 90.695 -201.805 91.860 ;
        RECT -201.635 90.695 -201.355 91.835 ;
        RECT -200.685 90.695 -200.425 91.835 ;
        RECT -193.555 90.695 -193.295 91.835 ;
        RECT -192.625 90.695 -192.345 91.835 ;
        RECT -192.175 90.695 -191.885 91.860 ;
        RECT -191.715 90.695 -191.435 91.835 ;
        RECT -190.765 90.695 -190.505 91.835 ;
        RECT -183.635 90.695 -183.375 91.835 ;
        RECT -182.705 90.695 -182.425 91.835 ;
        RECT -182.255 90.695 -181.965 91.860 ;
        RECT -181.795 90.695 -181.515 91.835 ;
        RECT -180.845 90.695 -180.585 91.835 ;
        RECT -173.715 90.695 -173.455 91.835 ;
        RECT -172.785 90.695 -172.505 91.835 ;
        RECT -172.335 90.695 -172.045 91.860 ;
        RECT -171.875 90.695 -171.595 91.835 ;
        RECT -170.925 90.695 -170.665 91.835 ;
        RECT -163.795 90.695 -163.535 91.835 ;
        RECT -162.865 90.695 -162.585 91.835 ;
        RECT -162.415 90.695 -162.125 91.860 ;
        RECT -161.955 90.695 -161.675 91.835 ;
        RECT -161.005 90.695 -160.745 91.835 ;
        RECT -153.875 90.695 -153.615 91.835 ;
        RECT -152.945 90.695 -152.665 91.835 ;
        RECT -152.495 90.695 -152.205 91.860 ;
        RECT -152.035 90.695 -151.755 91.835 ;
        RECT -151.085 90.695 -150.825 91.835 ;
        RECT -143.955 90.695 -143.695 91.835 ;
        RECT -143.025 90.695 -142.745 91.835 ;
        RECT -142.575 90.695 -142.285 91.860 ;
        RECT -142.115 90.695 -141.835 91.835 ;
        RECT -141.165 90.695 -140.905 91.835 ;
        RECT -134.035 90.695 -133.775 91.835 ;
        RECT -133.105 90.695 -132.825 91.835 ;
        RECT -132.655 90.695 -132.365 91.860 ;
        RECT -132.195 90.695 -131.915 91.835 ;
        RECT -131.245 90.695 -130.985 91.835 ;
        RECT -124.115 90.695 -123.855 91.835 ;
        RECT -123.185 90.695 -122.905 91.835 ;
        RECT -122.735 90.695 -122.445 91.860 ;
        RECT -122.275 90.695 -121.995 91.835 ;
        RECT -121.325 90.695 -121.065 91.835 ;
        RECT -114.195 90.695 -113.935 91.835 ;
        RECT -113.265 90.695 -112.985 91.835 ;
        RECT -112.815 90.695 -112.525 91.860 ;
        RECT -112.355 90.695 -112.075 91.835 ;
        RECT -111.405 90.695 -111.145 91.835 ;
        RECT -104.275 90.695 -104.015 91.835 ;
        RECT -103.345 90.695 -103.065 91.835 ;
        RECT -102.895 90.695 -102.605 91.860 ;
        RECT -102.435 90.695 -102.155 91.835 ;
        RECT -101.485 90.695 -101.225 91.835 ;
        RECT -94.355 90.695 -94.095 91.835 ;
        RECT -93.425 90.695 -93.145 91.835 ;
        RECT -92.975 90.695 -92.685 91.860 ;
        RECT -92.515 90.695 -92.235 91.835 ;
        RECT -91.565 90.695 -91.305 91.835 ;
        RECT -84.435 90.695 -84.175 91.835 ;
        RECT -83.505 90.695 -83.225 91.835 ;
        RECT -83.055 90.695 -82.765 91.860 ;
        RECT -82.595 90.695 -82.315 91.835 ;
        RECT -81.645 90.695 -81.385 91.835 ;
        RECT -74.515 90.695 -74.255 91.835 ;
        RECT -73.585 90.695 -73.305 91.835 ;
        RECT -73.135 90.695 -72.845 91.860 ;
        RECT -72.675 90.695 -72.395 91.835 ;
        RECT -71.725 90.695 -71.465 91.835 ;
        RECT -64.595 90.695 -64.335 91.835 ;
        RECT -63.665 90.695 -63.385 91.835 ;
        RECT -63.215 90.695 -62.925 91.860 ;
        RECT -62.755 90.695 -62.475 91.835 ;
        RECT -61.805 90.695 -61.545 91.835 ;
        RECT -54.675 90.695 -54.415 91.835 ;
        RECT -53.745 90.695 -53.465 91.835 ;
        RECT -53.295 90.695 -53.005 91.860 ;
        RECT -52.835 90.695 -52.555 91.835 ;
        RECT -51.885 90.695 -51.625 91.835 ;
        RECT -44.755 90.695 -44.495 91.835 ;
        RECT -43.825 90.695 -43.545 91.835 ;
        RECT -43.375 90.695 -43.085 91.860 ;
        RECT -42.915 90.695 -42.635 91.835 ;
        RECT -41.965 90.695 -41.705 91.835 ;
        RECT -34.835 90.695 -34.575 91.835 ;
        RECT -33.905 90.695 -33.625 91.835 ;
        RECT -33.455 90.695 -33.165 91.860 ;
        RECT -32.995 90.695 -32.715 91.835 ;
        RECT -32.045 90.695 -31.785 91.835 ;
        RECT -24.915 90.695 -24.655 91.835 ;
        RECT -23.985 90.695 -23.705 91.835 ;
        RECT -23.535 90.695 -23.245 91.860 ;
        RECT -23.075 90.695 -22.795 91.835 ;
        RECT -22.125 90.695 -21.865 91.835 ;
        RECT -14.995 90.695 -14.735 91.835 ;
        RECT -14.065 90.695 -13.785 91.835 ;
        RECT -13.615 90.695 -13.325 91.860 ;
        RECT -13.155 90.695 -12.875 91.835 ;
        RECT -12.205 90.695 -11.945 91.835 ;
        RECT -5.075 90.695 -4.815 91.835 ;
        RECT -4.145 90.695 -3.865 91.835 ;
        RECT -3.695 90.695 -3.405 91.860 ;
        RECT -3.235 90.695 -2.955 91.835 ;
        RECT -2.285 90.695 -2.025 91.835 ;
        RECT 4.845 90.695 5.105 91.835 ;
        RECT 5.775 90.695 6.055 91.835 ;
        RECT 6.225 90.695 6.515 91.860 ;
        RECT 6.685 90.695 6.965 91.835 ;
        RECT 7.635 90.695 7.895 91.835 ;
        RECT 14.765 90.695 15.025 91.835 ;
        RECT 15.695 90.695 15.975 91.835 ;
        RECT 16.145 90.695 16.435 91.860 ;
        RECT 16.605 90.695 16.885 91.835 ;
        RECT 17.555 90.695 17.815 91.835 ;
        RECT 24.685 90.695 24.945 91.835 ;
        RECT 25.615 90.695 25.895 91.835 ;
        RECT 26.065 90.695 26.355 91.860 ;
        RECT -282.920 90.525 -279.700 90.695 ;
        RECT -273.000 90.525 -269.780 90.695 ;
        RECT -263.080 90.525 -259.860 90.695 ;
        RECT -253.160 90.525 -249.940 90.695 ;
        RECT -243.240 90.525 -240.020 90.695 ;
        RECT -233.320 90.525 -230.100 90.695 ;
        RECT -223.400 90.525 -220.180 90.695 ;
        RECT -213.480 90.525 -210.260 90.695 ;
        RECT -203.560 90.525 -200.340 90.695 ;
        RECT -193.640 90.525 -190.420 90.695 ;
        RECT -183.720 90.525 -180.500 90.695 ;
        RECT -173.800 90.525 -170.580 90.695 ;
        RECT -163.880 90.525 -160.660 90.695 ;
        RECT -153.960 90.525 -150.740 90.695 ;
        RECT -144.040 90.525 -140.820 90.695 ;
        RECT -134.120 90.525 -130.900 90.695 ;
        RECT -124.200 90.525 -120.980 90.695 ;
        RECT -114.280 90.525 -111.060 90.695 ;
        RECT -104.360 90.525 -101.140 90.695 ;
        RECT -94.440 90.525 -91.220 90.695 ;
        RECT -84.520 90.525 -81.300 90.695 ;
        RECT -74.600 90.525 -71.380 90.695 ;
        RECT -64.680 90.525 -61.460 90.695 ;
        RECT -54.760 90.525 -51.540 90.695 ;
        RECT -44.840 90.525 -41.620 90.695 ;
        RECT -34.920 90.525 -31.700 90.695 ;
        RECT -25.000 90.525 -21.780 90.695 ;
        RECT -15.080 90.525 -11.860 90.695 ;
        RECT -5.160 90.525 -1.940 90.695 ;
        RECT 4.760 90.525 7.980 90.695 ;
        RECT 14.680 90.525 17.900 90.695 ;
        RECT 24.600 90.525 26.440 90.695 ;
        RECT -286.825 90.110 -286.655 90.180 ;
        RECT -285.885 90.110 -285.715 90.180 ;
        RECT -286.825 89.940 -285.715 90.110 ;
        RECT -286.825 89.655 -286.655 89.940 ;
        RECT -287.585 89.325 -286.655 89.655 ;
        RECT -286.825 88.800 -286.655 89.325 ;
        RECT -286.415 88.775 -286.125 89.940 ;
        RECT -285.885 89.655 -285.715 89.940 ;
        RECT -276.905 90.110 -276.735 90.180 ;
        RECT -275.965 90.110 -275.795 90.180 ;
        RECT -276.905 89.940 -275.795 90.110 ;
        RECT -276.905 89.655 -276.735 89.940 ;
        RECT -285.885 89.325 -284.955 89.655 ;
        RECT -277.665 89.325 -276.735 89.655 ;
        RECT -285.885 88.800 -285.715 89.325 ;
        RECT -276.905 88.800 -276.735 89.325 ;
        RECT -276.495 88.775 -276.205 89.940 ;
        RECT -275.965 89.655 -275.795 89.940 ;
        RECT -266.985 90.110 -266.815 90.180 ;
        RECT -266.045 90.110 -265.875 90.180 ;
        RECT -266.985 89.940 -265.875 90.110 ;
        RECT -266.985 89.655 -266.815 89.940 ;
        RECT -275.965 89.325 -275.035 89.655 ;
        RECT -267.745 89.325 -266.815 89.655 ;
        RECT -275.965 88.800 -275.795 89.325 ;
        RECT -266.985 88.800 -266.815 89.325 ;
        RECT -266.575 88.775 -266.285 89.940 ;
        RECT -266.045 89.655 -265.875 89.940 ;
        RECT -257.065 90.110 -256.895 90.180 ;
        RECT -256.125 90.110 -255.955 90.180 ;
        RECT -257.065 89.940 -255.955 90.110 ;
        RECT -257.065 89.655 -256.895 89.940 ;
        RECT -266.045 89.325 -265.115 89.655 ;
        RECT -257.825 89.325 -256.895 89.655 ;
        RECT -266.045 88.800 -265.875 89.325 ;
        RECT -257.065 88.800 -256.895 89.325 ;
        RECT -256.655 88.775 -256.365 89.940 ;
        RECT -256.125 89.655 -255.955 89.940 ;
        RECT -247.145 90.110 -246.975 90.180 ;
        RECT -246.205 90.110 -246.035 90.180 ;
        RECT -247.145 89.940 -246.035 90.110 ;
        RECT -247.145 89.655 -246.975 89.940 ;
        RECT -256.125 89.325 -255.195 89.655 ;
        RECT -247.905 89.325 -246.975 89.655 ;
        RECT -256.125 88.800 -255.955 89.325 ;
        RECT -247.145 88.800 -246.975 89.325 ;
        RECT -246.735 88.775 -246.445 89.940 ;
        RECT -246.205 89.655 -246.035 89.940 ;
        RECT -237.225 90.110 -237.055 90.180 ;
        RECT -236.285 90.110 -236.115 90.180 ;
        RECT -237.225 89.940 -236.115 90.110 ;
        RECT -237.225 89.655 -237.055 89.940 ;
        RECT -246.205 89.325 -245.275 89.655 ;
        RECT -237.985 89.325 -237.055 89.655 ;
        RECT -246.205 88.800 -246.035 89.325 ;
        RECT -237.225 88.800 -237.055 89.325 ;
        RECT -236.815 88.775 -236.525 89.940 ;
        RECT -236.285 89.655 -236.115 89.940 ;
        RECT -227.305 90.110 -227.135 90.180 ;
        RECT -226.365 90.110 -226.195 90.180 ;
        RECT -227.305 89.940 -226.195 90.110 ;
        RECT -227.305 89.655 -227.135 89.940 ;
        RECT -236.285 89.325 -235.355 89.655 ;
        RECT -228.065 89.325 -227.135 89.655 ;
        RECT -236.285 88.800 -236.115 89.325 ;
        RECT -227.305 88.800 -227.135 89.325 ;
        RECT -226.895 88.775 -226.605 89.940 ;
        RECT -226.365 89.655 -226.195 89.940 ;
        RECT -217.385 90.110 -217.215 90.180 ;
        RECT -216.445 90.110 -216.275 90.180 ;
        RECT -217.385 89.940 -216.275 90.110 ;
        RECT -217.385 89.655 -217.215 89.940 ;
        RECT -226.365 89.325 -225.435 89.655 ;
        RECT -218.145 89.325 -217.215 89.655 ;
        RECT -226.365 88.800 -226.195 89.325 ;
        RECT -217.385 88.800 -217.215 89.325 ;
        RECT -216.975 88.775 -216.685 89.940 ;
        RECT -216.445 89.655 -216.275 89.940 ;
        RECT -207.465 90.110 -207.295 90.180 ;
        RECT -206.525 90.110 -206.355 90.180 ;
        RECT -207.465 89.940 -206.355 90.110 ;
        RECT -207.465 89.655 -207.295 89.940 ;
        RECT -216.445 89.325 -215.515 89.655 ;
        RECT -208.225 89.325 -207.295 89.655 ;
        RECT -216.445 88.800 -216.275 89.325 ;
        RECT -207.465 88.800 -207.295 89.325 ;
        RECT -207.055 88.775 -206.765 89.940 ;
        RECT -206.525 89.655 -206.355 89.940 ;
        RECT -197.545 90.110 -197.375 90.180 ;
        RECT -196.605 90.110 -196.435 90.180 ;
        RECT -197.545 89.940 -196.435 90.110 ;
        RECT -197.545 89.655 -197.375 89.940 ;
        RECT -206.525 89.325 -205.595 89.655 ;
        RECT -198.305 89.325 -197.375 89.655 ;
        RECT -206.525 88.800 -206.355 89.325 ;
        RECT -197.545 88.800 -197.375 89.325 ;
        RECT -197.135 88.775 -196.845 89.940 ;
        RECT -196.605 89.655 -196.435 89.940 ;
        RECT -187.625 90.110 -187.455 90.180 ;
        RECT -186.685 90.110 -186.515 90.180 ;
        RECT -187.625 89.940 -186.515 90.110 ;
        RECT -187.625 89.655 -187.455 89.940 ;
        RECT -196.605 89.325 -195.675 89.655 ;
        RECT -188.385 89.325 -187.455 89.655 ;
        RECT -196.605 88.800 -196.435 89.325 ;
        RECT -187.625 88.800 -187.455 89.325 ;
        RECT -187.215 88.775 -186.925 89.940 ;
        RECT -186.685 89.655 -186.515 89.940 ;
        RECT -177.705 90.110 -177.535 90.180 ;
        RECT -176.765 90.110 -176.595 90.180 ;
        RECT -177.705 89.940 -176.595 90.110 ;
        RECT -177.705 89.655 -177.535 89.940 ;
        RECT -186.685 89.325 -185.755 89.655 ;
        RECT -178.465 89.325 -177.535 89.655 ;
        RECT -186.685 88.800 -186.515 89.325 ;
        RECT -177.705 88.800 -177.535 89.325 ;
        RECT -177.295 88.775 -177.005 89.940 ;
        RECT -176.765 89.655 -176.595 89.940 ;
        RECT -167.785 90.110 -167.615 90.180 ;
        RECT -166.845 90.110 -166.675 90.180 ;
        RECT -167.785 89.940 -166.675 90.110 ;
        RECT -167.785 89.655 -167.615 89.940 ;
        RECT -176.765 89.325 -175.835 89.655 ;
        RECT -168.545 89.325 -167.615 89.655 ;
        RECT -176.765 88.800 -176.595 89.325 ;
        RECT -167.785 88.800 -167.615 89.325 ;
        RECT -167.375 88.775 -167.085 89.940 ;
        RECT -166.845 89.655 -166.675 89.940 ;
        RECT -157.865 90.110 -157.695 90.180 ;
        RECT -156.925 90.110 -156.755 90.180 ;
        RECT -157.865 89.940 -156.755 90.110 ;
        RECT -157.865 89.655 -157.695 89.940 ;
        RECT -166.845 89.325 -165.915 89.655 ;
        RECT -158.625 89.325 -157.695 89.655 ;
        RECT -166.845 88.800 -166.675 89.325 ;
        RECT -157.865 88.800 -157.695 89.325 ;
        RECT -157.455 88.775 -157.165 89.940 ;
        RECT -156.925 89.655 -156.755 89.940 ;
        RECT -147.945 90.110 -147.775 90.180 ;
        RECT -147.005 90.110 -146.835 90.180 ;
        RECT -147.945 89.940 -146.835 90.110 ;
        RECT -147.945 89.655 -147.775 89.940 ;
        RECT -156.925 89.325 -155.995 89.655 ;
        RECT -148.705 89.325 -147.775 89.655 ;
        RECT -156.925 88.800 -156.755 89.325 ;
        RECT -147.945 88.800 -147.775 89.325 ;
        RECT -147.535 88.775 -147.245 89.940 ;
        RECT -147.005 89.655 -146.835 89.940 ;
        RECT -138.025 90.110 -137.855 90.180 ;
        RECT -137.085 90.110 -136.915 90.180 ;
        RECT -138.025 89.940 -136.915 90.110 ;
        RECT -138.025 89.655 -137.855 89.940 ;
        RECT -147.005 89.325 -146.075 89.655 ;
        RECT -138.785 89.325 -137.855 89.655 ;
        RECT -147.005 88.800 -146.835 89.325 ;
        RECT -138.025 88.800 -137.855 89.325 ;
        RECT -137.615 88.775 -137.325 89.940 ;
        RECT -137.085 89.655 -136.915 89.940 ;
        RECT -128.105 90.110 -127.935 90.180 ;
        RECT -127.165 90.110 -126.995 90.180 ;
        RECT -128.105 89.940 -126.995 90.110 ;
        RECT -128.105 89.655 -127.935 89.940 ;
        RECT -137.085 89.325 -136.155 89.655 ;
        RECT -128.865 89.325 -127.935 89.655 ;
        RECT -137.085 88.800 -136.915 89.325 ;
        RECT -128.105 88.800 -127.935 89.325 ;
        RECT -127.695 88.775 -127.405 89.940 ;
        RECT -127.165 89.655 -126.995 89.940 ;
        RECT -118.185 90.110 -118.015 90.180 ;
        RECT -117.245 90.110 -117.075 90.180 ;
        RECT -118.185 89.940 -117.075 90.110 ;
        RECT -118.185 89.655 -118.015 89.940 ;
        RECT -127.165 89.325 -126.235 89.655 ;
        RECT -118.945 89.325 -118.015 89.655 ;
        RECT -127.165 88.800 -126.995 89.325 ;
        RECT -118.185 88.800 -118.015 89.325 ;
        RECT -117.775 88.775 -117.485 89.940 ;
        RECT -117.245 89.655 -117.075 89.940 ;
        RECT -108.265 90.110 -108.095 90.180 ;
        RECT -107.325 90.110 -107.155 90.180 ;
        RECT -108.265 89.940 -107.155 90.110 ;
        RECT -108.265 89.655 -108.095 89.940 ;
        RECT -117.245 89.325 -116.315 89.655 ;
        RECT -109.025 89.325 -108.095 89.655 ;
        RECT -117.245 88.800 -117.075 89.325 ;
        RECT -108.265 88.800 -108.095 89.325 ;
        RECT -107.855 88.775 -107.565 89.940 ;
        RECT -107.325 89.655 -107.155 89.940 ;
        RECT -98.345 90.110 -98.175 90.180 ;
        RECT -97.405 90.110 -97.235 90.180 ;
        RECT -98.345 89.940 -97.235 90.110 ;
        RECT -98.345 89.655 -98.175 89.940 ;
        RECT -107.325 89.325 -106.395 89.655 ;
        RECT -99.105 89.325 -98.175 89.655 ;
        RECT -107.325 88.800 -107.155 89.325 ;
        RECT -98.345 88.800 -98.175 89.325 ;
        RECT -97.935 88.775 -97.645 89.940 ;
        RECT -97.405 89.655 -97.235 89.940 ;
        RECT -88.425 90.110 -88.255 90.180 ;
        RECT -87.485 90.110 -87.315 90.180 ;
        RECT -88.425 89.940 -87.315 90.110 ;
        RECT -88.425 89.655 -88.255 89.940 ;
        RECT -97.405 89.325 -96.475 89.655 ;
        RECT -89.185 89.325 -88.255 89.655 ;
        RECT -97.405 88.800 -97.235 89.325 ;
        RECT -88.425 88.800 -88.255 89.325 ;
        RECT -88.015 88.775 -87.725 89.940 ;
        RECT -87.485 89.655 -87.315 89.940 ;
        RECT -78.505 90.110 -78.335 90.180 ;
        RECT -77.565 90.110 -77.395 90.180 ;
        RECT -78.505 89.940 -77.395 90.110 ;
        RECT -78.505 89.655 -78.335 89.940 ;
        RECT -87.485 89.325 -86.555 89.655 ;
        RECT -79.265 89.325 -78.335 89.655 ;
        RECT -87.485 88.800 -87.315 89.325 ;
        RECT -78.505 88.800 -78.335 89.325 ;
        RECT -78.095 88.775 -77.805 89.940 ;
        RECT -77.565 89.655 -77.395 89.940 ;
        RECT -68.585 90.110 -68.415 90.180 ;
        RECT -67.645 90.110 -67.475 90.180 ;
        RECT -68.585 89.940 -67.475 90.110 ;
        RECT -68.585 89.655 -68.415 89.940 ;
        RECT -77.565 89.325 -76.635 89.655 ;
        RECT -69.345 89.325 -68.415 89.655 ;
        RECT -77.565 88.800 -77.395 89.325 ;
        RECT -68.585 88.800 -68.415 89.325 ;
        RECT -68.175 88.775 -67.885 89.940 ;
        RECT -67.645 89.655 -67.475 89.940 ;
        RECT -58.665 90.110 -58.495 90.180 ;
        RECT -57.725 90.110 -57.555 90.180 ;
        RECT -58.665 89.940 -57.555 90.110 ;
        RECT -58.665 89.655 -58.495 89.940 ;
        RECT -67.645 89.325 -66.715 89.655 ;
        RECT -59.425 89.325 -58.495 89.655 ;
        RECT -67.645 88.800 -67.475 89.325 ;
        RECT -58.665 88.800 -58.495 89.325 ;
        RECT -58.255 88.775 -57.965 89.940 ;
        RECT -57.725 89.655 -57.555 89.940 ;
        RECT -48.745 90.110 -48.575 90.180 ;
        RECT -47.805 90.110 -47.635 90.180 ;
        RECT -48.745 89.940 -47.635 90.110 ;
        RECT -48.745 89.655 -48.575 89.940 ;
        RECT -57.725 89.325 -56.795 89.655 ;
        RECT -49.505 89.325 -48.575 89.655 ;
        RECT -57.725 88.800 -57.555 89.325 ;
        RECT -48.745 88.800 -48.575 89.325 ;
        RECT -48.335 88.775 -48.045 89.940 ;
        RECT -47.805 89.655 -47.635 89.940 ;
        RECT -38.825 90.110 -38.655 90.180 ;
        RECT -37.885 90.110 -37.715 90.180 ;
        RECT -38.825 89.940 -37.715 90.110 ;
        RECT -38.825 89.655 -38.655 89.940 ;
        RECT -47.805 89.325 -46.875 89.655 ;
        RECT -39.585 89.325 -38.655 89.655 ;
        RECT -47.805 88.800 -47.635 89.325 ;
        RECT -38.825 88.800 -38.655 89.325 ;
        RECT -38.415 88.775 -38.125 89.940 ;
        RECT -37.885 89.655 -37.715 89.940 ;
        RECT -28.905 90.110 -28.735 90.180 ;
        RECT -27.965 90.110 -27.795 90.180 ;
        RECT -28.905 89.940 -27.795 90.110 ;
        RECT -28.905 89.655 -28.735 89.940 ;
        RECT -37.885 89.325 -36.955 89.655 ;
        RECT -29.665 89.325 -28.735 89.655 ;
        RECT -37.885 88.800 -37.715 89.325 ;
        RECT -28.905 88.800 -28.735 89.325 ;
        RECT -28.495 88.775 -28.205 89.940 ;
        RECT -27.965 89.655 -27.795 89.940 ;
        RECT -18.985 90.110 -18.815 90.180 ;
        RECT -18.045 90.110 -17.875 90.180 ;
        RECT -18.985 89.940 -17.875 90.110 ;
        RECT -18.985 89.655 -18.815 89.940 ;
        RECT -27.965 89.325 -27.035 89.655 ;
        RECT -19.745 89.325 -18.815 89.655 ;
        RECT -27.965 88.800 -27.795 89.325 ;
        RECT -18.985 88.800 -18.815 89.325 ;
        RECT -18.575 88.775 -18.285 89.940 ;
        RECT -18.045 89.655 -17.875 89.940 ;
        RECT -9.065 90.110 -8.895 90.180 ;
        RECT -8.125 90.110 -7.955 90.180 ;
        RECT -9.065 89.940 -7.955 90.110 ;
        RECT -9.065 89.655 -8.895 89.940 ;
        RECT -18.045 89.325 -17.115 89.655 ;
        RECT -9.825 89.325 -8.895 89.655 ;
        RECT -18.045 88.800 -17.875 89.325 ;
        RECT -9.065 88.800 -8.895 89.325 ;
        RECT -8.655 88.775 -8.365 89.940 ;
        RECT -8.125 89.655 -7.955 89.940 ;
        RECT 0.855 90.110 1.025 90.180 ;
        RECT 1.795 90.110 1.965 90.180 ;
        RECT 0.855 89.940 1.965 90.110 ;
        RECT 0.855 89.655 1.025 89.940 ;
        RECT -8.125 89.325 -7.195 89.655 ;
        RECT 0.095 89.325 1.025 89.655 ;
        RECT -8.125 88.800 -7.955 89.325 ;
        RECT 0.855 88.800 1.025 89.325 ;
        RECT 1.265 88.775 1.555 89.940 ;
        RECT 1.795 89.655 1.965 89.940 ;
        RECT 10.775 90.110 10.945 90.180 ;
        RECT 11.715 90.110 11.885 90.180 ;
        RECT 10.775 89.940 11.885 90.110 ;
        RECT 10.775 89.655 10.945 89.940 ;
        RECT 1.795 89.325 2.725 89.655 ;
        RECT 10.015 89.325 10.945 89.655 ;
        RECT 1.795 88.800 1.965 89.325 ;
        RECT 10.775 88.800 10.945 89.325 ;
        RECT 11.185 88.775 11.475 89.940 ;
        RECT 11.715 89.655 11.885 89.940 ;
        RECT 20.695 90.110 20.865 90.180 ;
        RECT 21.635 90.110 21.805 90.180 ;
        RECT 20.695 89.940 21.805 90.110 ;
        RECT 20.695 89.655 20.865 89.940 ;
        RECT 11.715 89.325 12.645 89.655 ;
        RECT 19.935 89.325 20.865 89.655 ;
        RECT 11.715 88.800 11.885 89.325 ;
        RECT 20.695 88.800 20.865 89.325 ;
        RECT 21.105 88.775 21.395 89.940 ;
        RECT 21.635 89.655 21.805 89.940 ;
        RECT 21.635 89.325 22.565 89.655 ;
        RECT 21.635 88.800 21.805 89.325 ;
      LAYER mcon ;
        RECT -281.865 94.825 -281.695 94.995 ;
        RECT -281.395 94.820 -281.225 94.990 ;
        RECT -280.925 94.825 -280.755 94.995 ;
        RECT -281.865 94.365 -281.695 94.535 ;
        RECT -281.865 93.905 -281.695 94.075 ;
        RECT -271.945 94.825 -271.775 94.995 ;
        RECT -271.475 94.820 -271.305 94.990 ;
        RECT -271.005 94.825 -270.835 94.995 ;
        RECT -280.925 94.365 -280.755 94.535 ;
        RECT -271.945 94.365 -271.775 94.535 ;
        RECT -280.925 93.905 -280.755 94.075 ;
        RECT -271.945 93.905 -271.775 94.075 ;
        RECT -262.025 94.825 -261.855 94.995 ;
        RECT -261.555 94.820 -261.385 94.990 ;
        RECT -261.085 94.825 -260.915 94.995 ;
        RECT -271.005 94.365 -270.835 94.535 ;
        RECT -262.025 94.365 -261.855 94.535 ;
        RECT -271.005 93.905 -270.835 94.075 ;
        RECT -262.025 93.905 -261.855 94.075 ;
        RECT -252.105 94.825 -251.935 94.995 ;
        RECT -251.635 94.820 -251.465 94.990 ;
        RECT -251.165 94.825 -250.995 94.995 ;
        RECT -261.085 94.365 -260.915 94.535 ;
        RECT -252.105 94.365 -251.935 94.535 ;
        RECT -261.085 93.905 -260.915 94.075 ;
        RECT -252.105 93.905 -251.935 94.075 ;
        RECT -242.185 94.825 -242.015 94.995 ;
        RECT -241.715 94.820 -241.545 94.990 ;
        RECT -241.245 94.825 -241.075 94.995 ;
        RECT -251.165 94.365 -250.995 94.535 ;
        RECT -242.185 94.365 -242.015 94.535 ;
        RECT -251.165 93.905 -250.995 94.075 ;
        RECT -242.185 93.905 -242.015 94.075 ;
        RECT -232.265 94.825 -232.095 94.995 ;
        RECT -231.795 94.820 -231.625 94.990 ;
        RECT -231.325 94.825 -231.155 94.995 ;
        RECT -241.245 94.365 -241.075 94.535 ;
        RECT -232.265 94.365 -232.095 94.535 ;
        RECT -241.245 93.905 -241.075 94.075 ;
        RECT -232.265 93.905 -232.095 94.075 ;
        RECT -222.345 94.825 -222.175 94.995 ;
        RECT -221.875 94.820 -221.705 94.990 ;
        RECT -221.405 94.825 -221.235 94.995 ;
        RECT -231.325 94.365 -231.155 94.535 ;
        RECT -222.345 94.365 -222.175 94.535 ;
        RECT -231.325 93.905 -231.155 94.075 ;
        RECT -222.345 93.905 -222.175 94.075 ;
        RECT -212.425 94.825 -212.255 94.995 ;
        RECT -211.955 94.820 -211.785 94.990 ;
        RECT -211.485 94.825 -211.315 94.995 ;
        RECT -221.405 94.365 -221.235 94.535 ;
        RECT -212.425 94.365 -212.255 94.535 ;
        RECT -221.405 93.905 -221.235 94.075 ;
        RECT -212.425 93.905 -212.255 94.075 ;
        RECT -202.505 94.825 -202.335 94.995 ;
        RECT -202.035 94.820 -201.865 94.990 ;
        RECT -201.565 94.825 -201.395 94.995 ;
        RECT -211.485 94.365 -211.315 94.535 ;
        RECT -202.505 94.365 -202.335 94.535 ;
        RECT -211.485 93.905 -211.315 94.075 ;
        RECT -202.505 93.905 -202.335 94.075 ;
        RECT -192.585 94.825 -192.415 94.995 ;
        RECT -192.115 94.820 -191.945 94.990 ;
        RECT -191.645 94.825 -191.475 94.995 ;
        RECT -201.565 94.365 -201.395 94.535 ;
        RECT -192.585 94.365 -192.415 94.535 ;
        RECT -201.565 93.905 -201.395 94.075 ;
        RECT -192.585 93.905 -192.415 94.075 ;
        RECT -182.665 94.825 -182.495 94.995 ;
        RECT -182.195 94.820 -182.025 94.990 ;
        RECT -181.725 94.825 -181.555 94.995 ;
        RECT -191.645 94.365 -191.475 94.535 ;
        RECT -182.665 94.365 -182.495 94.535 ;
        RECT -191.645 93.905 -191.475 94.075 ;
        RECT -182.665 93.905 -182.495 94.075 ;
        RECT -172.745 94.825 -172.575 94.995 ;
        RECT -172.275 94.820 -172.105 94.990 ;
        RECT -171.805 94.825 -171.635 94.995 ;
        RECT -181.725 94.365 -181.555 94.535 ;
        RECT -172.745 94.365 -172.575 94.535 ;
        RECT -181.725 93.905 -181.555 94.075 ;
        RECT -172.745 93.905 -172.575 94.075 ;
        RECT -162.825 94.825 -162.655 94.995 ;
        RECT -162.355 94.820 -162.185 94.990 ;
        RECT -161.885 94.825 -161.715 94.995 ;
        RECT -171.805 94.365 -171.635 94.535 ;
        RECT -162.825 94.365 -162.655 94.535 ;
        RECT -171.805 93.905 -171.635 94.075 ;
        RECT -162.825 93.905 -162.655 94.075 ;
        RECT -152.905 94.825 -152.735 94.995 ;
        RECT -152.435 94.820 -152.265 94.990 ;
        RECT -151.965 94.825 -151.795 94.995 ;
        RECT -161.885 94.365 -161.715 94.535 ;
        RECT -152.905 94.365 -152.735 94.535 ;
        RECT -161.885 93.905 -161.715 94.075 ;
        RECT -152.905 93.905 -152.735 94.075 ;
        RECT -142.985 94.825 -142.815 94.995 ;
        RECT -142.515 94.820 -142.345 94.990 ;
        RECT -142.045 94.825 -141.875 94.995 ;
        RECT -151.965 94.365 -151.795 94.535 ;
        RECT -142.985 94.365 -142.815 94.535 ;
        RECT -151.965 93.905 -151.795 94.075 ;
        RECT -142.985 93.905 -142.815 94.075 ;
        RECT -133.065 94.825 -132.895 94.995 ;
        RECT -132.595 94.820 -132.425 94.990 ;
        RECT -132.125 94.825 -131.955 94.995 ;
        RECT -142.045 94.365 -141.875 94.535 ;
        RECT -133.065 94.365 -132.895 94.535 ;
        RECT -142.045 93.905 -141.875 94.075 ;
        RECT -133.065 93.905 -132.895 94.075 ;
        RECT -123.145 94.825 -122.975 94.995 ;
        RECT -122.675 94.820 -122.505 94.990 ;
        RECT -122.205 94.825 -122.035 94.995 ;
        RECT -132.125 94.365 -131.955 94.535 ;
        RECT -123.145 94.365 -122.975 94.535 ;
        RECT -132.125 93.905 -131.955 94.075 ;
        RECT -123.145 93.905 -122.975 94.075 ;
        RECT -113.225 94.825 -113.055 94.995 ;
        RECT -112.755 94.820 -112.585 94.990 ;
        RECT -112.285 94.825 -112.115 94.995 ;
        RECT -122.205 94.365 -122.035 94.535 ;
        RECT -113.225 94.365 -113.055 94.535 ;
        RECT -122.205 93.905 -122.035 94.075 ;
        RECT -113.225 93.905 -113.055 94.075 ;
        RECT -103.305 94.825 -103.135 94.995 ;
        RECT -102.835 94.820 -102.665 94.990 ;
        RECT -102.365 94.825 -102.195 94.995 ;
        RECT -112.285 94.365 -112.115 94.535 ;
        RECT -103.305 94.365 -103.135 94.535 ;
        RECT -112.285 93.905 -112.115 94.075 ;
        RECT -103.305 93.905 -103.135 94.075 ;
        RECT -93.385 94.825 -93.215 94.995 ;
        RECT -92.915 94.820 -92.745 94.990 ;
        RECT -92.445 94.825 -92.275 94.995 ;
        RECT -102.365 94.365 -102.195 94.535 ;
        RECT -93.385 94.365 -93.215 94.535 ;
        RECT -102.365 93.905 -102.195 94.075 ;
        RECT -93.385 93.905 -93.215 94.075 ;
        RECT -83.465 94.825 -83.295 94.995 ;
        RECT -82.995 94.820 -82.825 94.990 ;
        RECT -82.525 94.825 -82.355 94.995 ;
        RECT -92.445 94.365 -92.275 94.535 ;
        RECT -83.465 94.365 -83.295 94.535 ;
        RECT -92.445 93.905 -92.275 94.075 ;
        RECT -83.465 93.905 -83.295 94.075 ;
        RECT -73.545 94.825 -73.375 94.995 ;
        RECT -73.075 94.820 -72.905 94.990 ;
        RECT -72.605 94.825 -72.435 94.995 ;
        RECT -82.525 94.365 -82.355 94.535 ;
        RECT -73.545 94.365 -73.375 94.535 ;
        RECT -82.525 93.905 -82.355 94.075 ;
        RECT -73.545 93.905 -73.375 94.075 ;
        RECT -63.625 94.825 -63.455 94.995 ;
        RECT -63.155 94.820 -62.985 94.990 ;
        RECT -62.685 94.825 -62.515 94.995 ;
        RECT -72.605 94.365 -72.435 94.535 ;
        RECT -63.625 94.365 -63.455 94.535 ;
        RECT -72.605 93.905 -72.435 94.075 ;
        RECT -63.625 93.905 -63.455 94.075 ;
        RECT -53.705 94.825 -53.535 94.995 ;
        RECT -53.235 94.820 -53.065 94.990 ;
        RECT -52.765 94.825 -52.595 94.995 ;
        RECT -62.685 94.365 -62.515 94.535 ;
        RECT -53.705 94.365 -53.535 94.535 ;
        RECT -62.685 93.905 -62.515 94.075 ;
        RECT -53.705 93.905 -53.535 94.075 ;
        RECT -43.785 94.825 -43.615 94.995 ;
        RECT -43.315 94.820 -43.145 94.990 ;
        RECT -42.845 94.825 -42.675 94.995 ;
        RECT -52.765 94.365 -52.595 94.535 ;
        RECT -43.785 94.365 -43.615 94.535 ;
        RECT -52.765 93.905 -52.595 94.075 ;
        RECT -43.785 93.905 -43.615 94.075 ;
        RECT -33.865 94.825 -33.695 94.995 ;
        RECT -33.395 94.820 -33.225 94.990 ;
        RECT -32.925 94.825 -32.755 94.995 ;
        RECT -42.845 94.365 -42.675 94.535 ;
        RECT -33.865 94.365 -33.695 94.535 ;
        RECT -42.845 93.905 -42.675 94.075 ;
        RECT -33.865 93.905 -33.695 94.075 ;
        RECT -23.945 94.825 -23.775 94.995 ;
        RECT -23.475 94.820 -23.305 94.990 ;
        RECT -23.005 94.825 -22.835 94.995 ;
        RECT -32.925 94.365 -32.755 94.535 ;
        RECT -23.945 94.365 -23.775 94.535 ;
        RECT -32.925 93.905 -32.755 94.075 ;
        RECT -23.945 93.905 -23.775 94.075 ;
        RECT -14.025 94.825 -13.855 94.995 ;
        RECT -13.555 94.820 -13.385 94.990 ;
        RECT -13.085 94.825 -12.915 94.995 ;
        RECT -23.005 94.365 -22.835 94.535 ;
        RECT -14.025 94.365 -13.855 94.535 ;
        RECT -23.005 93.905 -22.835 94.075 ;
        RECT -14.025 93.905 -13.855 94.075 ;
        RECT -4.105 94.825 -3.935 94.995 ;
        RECT -3.635 94.820 -3.465 94.990 ;
        RECT -3.165 94.825 -2.995 94.995 ;
        RECT -13.085 94.365 -12.915 94.535 ;
        RECT -4.105 94.365 -3.935 94.535 ;
        RECT -13.085 93.905 -12.915 94.075 ;
        RECT -4.105 93.905 -3.935 94.075 ;
        RECT 5.815 94.825 5.985 94.995 ;
        RECT 6.285 94.820 6.455 94.990 ;
        RECT 6.755 94.825 6.925 94.995 ;
        RECT -3.165 94.365 -2.995 94.535 ;
        RECT 5.815 94.365 5.985 94.535 ;
        RECT -3.165 93.905 -2.995 94.075 ;
        RECT 5.815 93.905 5.985 94.075 ;
        RECT 15.735 94.825 15.905 94.995 ;
        RECT 16.205 94.820 16.375 94.990 ;
        RECT 16.675 94.825 16.845 94.995 ;
        RECT 6.755 94.365 6.925 94.535 ;
        RECT 15.735 94.365 15.905 94.535 ;
        RECT 6.755 93.905 6.925 94.075 ;
        RECT 15.735 93.905 15.905 94.075 ;
        RECT 25.655 94.825 25.825 94.995 ;
        RECT 26.125 94.820 26.295 94.990 ;
        RECT 16.675 94.365 16.845 94.535 ;
        RECT 25.655 94.365 25.825 94.535 ;
        RECT 16.675 93.905 16.845 94.075 ;
        RECT 25.655 93.905 25.825 94.075 ;
        RECT -287.735 93.245 -287.565 93.415 ;
        RECT -287.275 93.245 -287.105 93.415 ;
        RECT -286.815 93.245 -286.645 93.415 ;
        RECT -286.355 93.245 -286.185 93.415 ;
        RECT -285.895 93.245 -285.725 93.415 ;
        RECT -285.435 93.245 -285.265 93.415 ;
        RECT -284.975 93.245 -284.805 93.415 ;
        RECT -277.815 93.245 -277.645 93.415 ;
        RECT -277.355 93.245 -277.185 93.415 ;
        RECT -276.895 93.245 -276.725 93.415 ;
        RECT -276.435 93.245 -276.265 93.415 ;
        RECT -275.975 93.245 -275.805 93.415 ;
        RECT -275.515 93.245 -275.345 93.415 ;
        RECT -275.055 93.245 -274.885 93.415 ;
        RECT -267.895 93.245 -267.725 93.415 ;
        RECT -267.435 93.245 -267.265 93.415 ;
        RECT -266.975 93.245 -266.805 93.415 ;
        RECT -266.515 93.245 -266.345 93.415 ;
        RECT -266.055 93.245 -265.885 93.415 ;
        RECT -265.595 93.245 -265.425 93.415 ;
        RECT -265.135 93.245 -264.965 93.415 ;
        RECT -257.975 93.245 -257.805 93.415 ;
        RECT -257.515 93.245 -257.345 93.415 ;
        RECT -257.055 93.245 -256.885 93.415 ;
        RECT -256.595 93.245 -256.425 93.415 ;
        RECT -256.135 93.245 -255.965 93.415 ;
        RECT -255.675 93.245 -255.505 93.415 ;
        RECT -255.215 93.245 -255.045 93.415 ;
        RECT -248.055 93.245 -247.885 93.415 ;
        RECT -247.595 93.245 -247.425 93.415 ;
        RECT -247.135 93.245 -246.965 93.415 ;
        RECT -246.675 93.245 -246.505 93.415 ;
        RECT -246.215 93.245 -246.045 93.415 ;
        RECT -245.755 93.245 -245.585 93.415 ;
        RECT -245.295 93.245 -245.125 93.415 ;
        RECT -238.135 93.245 -237.965 93.415 ;
        RECT -237.675 93.245 -237.505 93.415 ;
        RECT -237.215 93.245 -237.045 93.415 ;
        RECT -236.755 93.245 -236.585 93.415 ;
        RECT -236.295 93.245 -236.125 93.415 ;
        RECT -235.835 93.245 -235.665 93.415 ;
        RECT -235.375 93.245 -235.205 93.415 ;
        RECT -228.215 93.245 -228.045 93.415 ;
        RECT -227.755 93.245 -227.585 93.415 ;
        RECT -227.295 93.245 -227.125 93.415 ;
        RECT -226.835 93.245 -226.665 93.415 ;
        RECT -226.375 93.245 -226.205 93.415 ;
        RECT -225.915 93.245 -225.745 93.415 ;
        RECT -225.455 93.245 -225.285 93.415 ;
        RECT -218.295 93.245 -218.125 93.415 ;
        RECT -217.835 93.245 -217.665 93.415 ;
        RECT -217.375 93.245 -217.205 93.415 ;
        RECT -216.915 93.245 -216.745 93.415 ;
        RECT -216.455 93.245 -216.285 93.415 ;
        RECT -215.995 93.245 -215.825 93.415 ;
        RECT -215.535 93.245 -215.365 93.415 ;
        RECT -208.375 93.245 -208.205 93.415 ;
        RECT -207.915 93.245 -207.745 93.415 ;
        RECT -207.455 93.245 -207.285 93.415 ;
        RECT -206.995 93.245 -206.825 93.415 ;
        RECT -206.535 93.245 -206.365 93.415 ;
        RECT -206.075 93.245 -205.905 93.415 ;
        RECT -205.615 93.245 -205.445 93.415 ;
        RECT -198.455 93.245 -198.285 93.415 ;
        RECT -197.995 93.245 -197.825 93.415 ;
        RECT -197.535 93.245 -197.365 93.415 ;
        RECT -197.075 93.245 -196.905 93.415 ;
        RECT -196.615 93.245 -196.445 93.415 ;
        RECT -196.155 93.245 -195.985 93.415 ;
        RECT -195.695 93.245 -195.525 93.415 ;
        RECT -188.535 93.245 -188.365 93.415 ;
        RECT -188.075 93.245 -187.905 93.415 ;
        RECT -187.615 93.245 -187.445 93.415 ;
        RECT -187.155 93.245 -186.985 93.415 ;
        RECT -186.695 93.245 -186.525 93.415 ;
        RECT -186.235 93.245 -186.065 93.415 ;
        RECT -185.775 93.245 -185.605 93.415 ;
        RECT -178.615 93.245 -178.445 93.415 ;
        RECT -178.155 93.245 -177.985 93.415 ;
        RECT -177.695 93.245 -177.525 93.415 ;
        RECT -177.235 93.245 -177.065 93.415 ;
        RECT -176.775 93.245 -176.605 93.415 ;
        RECT -176.315 93.245 -176.145 93.415 ;
        RECT -175.855 93.245 -175.685 93.415 ;
        RECT -168.695 93.245 -168.525 93.415 ;
        RECT -168.235 93.245 -168.065 93.415 ;
        RECT -167.775 93.245 -167.605 93.415 ;
        RECT -167.315 93.245 -167.145 93.415 ;
        RECT -166.855 93.245 -166.685 93.415 ;
        RECT -166.395 93.245 -166.225 93.415 ;
        RECT -165.935 93.245 -165.765 93.415 ;
        RECT -158.775 93.245 -158.605 93.415 ;
        RECT -158.315 93.245 -158.145 93.415 ;
        RECT -157.855 93.245 -157.685 93.415 ;
        RECT -157.395 93.245 -157.225 93.415 ;
        RECT -156.935 93.245 -156.765 93.415 ;
        RECT -156.475 93.245 -156.305 93.415 ;
        RECT -156.015 93.245 -155.845 93.415 ;
        RECT -148.855 93.245 -148.685 93.415 ;
        RECT -148.395 93.245 -148.225 93.415 ;
        RECT -147.935 93.245 -147.765 93.415 ;
        RECT -147.475 93.245 -147.305 93.415 ;
        RECT -147.015 93.245 -146.845 93.415 ;
        RECT -146.555 93.245 -146.385 93.415 ;
        RECT -146.095 93.245 -145.925 93.415 ;
        RECT -138.935 93.245 -138.765 93.415 ;
        RECT -138.475 93.245 -138.305 93.415 ;
        RECT -138.015 93.245 -137.845 93.415 ;
        RECT -137.555 93.245 -137.385 93.415 ;
        RECT -137.095 93.245 -136.925 93.415 ;
        RECT -136.635 93.245 -136.465 93.415 ;
        RECT -136.175 93.245 -136.005 93.415 ;
        RECT -129.015 93.245 -128.845 93.415 ;
        RECT -128.555 93.245 -128.385 93.415 ;
        RECT -128.095 93.245 -127.925 93.415 ;
        RECT -127.635 93.245 -127.465 93.415 ;
        RECT -127.175 93.245 -127.005 93.415 ;
        RECT -126.715 93.245 -126.545 93.415 ;
        RECT -126.255 93.245 -126.085 93.415 ;
        RECT -119.095 93.245 -118.925 93.415 ;
        RECT -118.635 93.245 -118.465 93.415 ;
        RECT -118.175 93.245 -118.005 93.415 ;
        RECT -117.715 93.245 -117.545 93.415 ;
        RECT -117.255 93.245 -117.085 93.415 ;
        RECT -116.795 93.245 -116.625 93.415 ;
        RECT -116.335 93.245 -116.165 93.415 ;
        RECT -109.175 93.245 -109.005 93.415 ;
        RECT -108.715 93.245 -108.545 93.415 ;
        RECT -108.255 93.245 -108.085 93.415 ;
        RECT -107.795 93.245 -107.625 93.415 ;
        RECT -107.335 93.245 -107.165 93.415 ;
        RECT -106.875 93.245 -106.705 93.415 ;
        RECT -106.415 93.245 -106.245 93.415 ;
        RECT -99.255 93.245 -99.085 93.415 ;
        RECT -98.795 93.245 -98.625 93.415 ;
        RECT -98.335 93.245 -98.165 93.415 ;
        RECT -97.875 93.245 -97.705 93.415 ;
        RECT -97.415 93.245 -97.245 93.415 ;
        RECT -96.955 93.245 -96.785 93.415 ;
        RECT -96.495 93.245 -96.325 93.415 ;
        RECT -89.335 93.245 -89.165 93.415 ;
        RECT -88.875 93.245 -88.705 93.415 ;
        RECT -88.415 93.245 -88.245 93.415 ;
        RECT -87.955 93.245 -87.785 93.415 ;
        RECT -87.495 93.245 -87.325 93.415 ;
        RECT -87.035 93.245 -86.865 93.415 ;
        RECT -86.575 93.245 -86.405 93.415 ;
        RECT -79.415 93.245 -79.245 93.415 ;
        RECT -78.955 93.245 -78.785 93.415 ;
        RECT -78.495 93.245 -78.325 93.415 ;
        RECT -78.035 93.245 -77.865 93.415 ;
        RECT -77.575 93.245 -77.405 93.415 ;
        RECT -77.115 93.245 -76.945 93.415 ;
        RECT -76.655 93.245 -76.485 93.415 ;
        RECT -69.495 93.245 -69.325 93.415 ;
        RECT -69.035 93.245 -68.865 93.415 ;
        RECT -68.575 93.245 -68.405 93.415 ;
        RECT -68.115 93.245 -67.945 93.415 ;
        RECT -67.655 93.245 -67.485 93.415 ;
        RECT -67.195 93.245 -67.025 93.415 ;
        RECT -66.735 93.245 -66.565 93.415 ;
        RECT -59.575 93.245 -59.405 93.415 ;
        RECT -59.115 93.245 -58.945 93.415 ;
        RECT -58.655 93.245 -58.485 93.415 ;
        RECT -58.195 93.245 -58.025 93.415 ;
        RECT -57.735 93.245 -57.565 93.415 ;
        RECT -57.275 93.245 -57.105 93.415 ;
        RECT -56.815 93.245 -56.645 93.415 ;
        RECT -49.655 93.245 -49.485 93.415 ;
        RECT -49.195 93.245 -49.025 93.415 ;
        RECT -48.735 93.245 -48.565 93.415 ;
        RECT -48.275 93.245 -48.105 93.415 ;
        RECT -47.815 93.245 -47.645 93.415 ;
        RECT -47.355 93.245 -47.185 93.415 ;
        RECT -46.895 93.245 -46.725 93.415 ;
        RECT -39.735 93.245 -39.565 93.415 ;
        RECT -39.275 93.245 -39.105 93.415 ;
        RECT -38.815 93.245 -38.645 93.415 ;
        RECT -38.355 93.245 -38.185 93.415 ;
        RECT -37.895 93.245 -37.725 93.415 ;
        RECT -37.435 93.245 -37.265 93.415 ;
        RECT -36.975 93.245 -36.805 93.415 ;
        RECT -29.815 93.245 -29.645 93.415 ;
        RECT -29.355 93.245 -29.185 93.415 ;
        RECT -28.895 93.245 -28.725 93.415 ;
        RECT -28.435 93.245 -28.265 93.415 ;
        RECT -27.975 93.245 -27.805 93.415 ;
        RECT -27.515 93.245 -27.345 93.415 ;
        RECT -27.055 93.245 -26.885 93.415 ;
        RECT -19.895 93.245 -19.725 93.415 ;
        RECT -19.435 93.245 -19.265 93.415 ;
        RECT -18.975 93.245 -18.805 93.415 ;
        RECT -18.515 93.245 -18.345 93.415 ;
        RECT -18.055 93.245 -17.885 93.415 ;
        RECT -17.595 93.245 -17.425 93.415 ;
        RECT -17.135 93.245 -16.965 93.415 ;
        RECT -9.975 93.245 -9.805 93.415 ;
        RECT -9.515 93.245 -9.345 93.415 ;
        RECT -9.055 93.245 -8.885 93.415 ;
        RECT -8.595 93.245 -8.425 93.415 ;
        RECT -8.135 93.245 -7.965 93.415 ;
        RECT -7.675 93.245 -7.505 93.415 ;
        RECT -7.215 93.245 -7.045 93.415 ;
        RECT -0.055 93.245 0.115 93.415 ;
        RECT 0.405 93.245 0.575 93.415 ;
        RECT 0.865 93.245 1.035 93.415 ;
        RECT 1.325 93.245 1.495 93.415 ;
        RECT 1.785 93.245 1.955 93.415 ;
        RECT 2.245 93.245 2.415 93.415 ;
        RECT 2.705 93.245 2.875 93.415 ;
        RECT 9.865 93.245 10.035 93.415 ;
        RECT 10.325 93.245 10.495 93.415 ;
        RECT 10.785 93.245 10.955 93.415 ;
        RECT 11.245 93.245 11.415 93.415 ;
        RECT 11.705 93.245 11.875 93.415 ;
        RECT 12.165 93.245 12.335 93.415 ;
        RECT 12.625 93.245 12.795 93.415 ;
        RECT 19.785 93.245 19.955 93.415 ;
        RECT 20.245 93.245 20.415 93.415 ;
        RECT 20.705 93.245 20.875 93.415 ;
        RECT 21.165 93.245 21.335 93.415 ;
        RECT 21.625 93.245 21.795 93.415 ;
        RECT 22.085 93.245 22.255 93.415 ;
        RECT 22.545 93.245 22.715 93.415 ;
        RECT -282.775 90.525 -282.605 90.695 ;
        RECT -282.315 90.525 -282.145 90.695 ;
        RECT -281.855 90.525 -281.685 90.695 ;
        RECT -281.395 90.525 -281.225 90.695 ;
        RECT -280.935 90.525 -280.765 90.695 ;
        RECT -280.475 90.525 -280.305 90.695 ;
        RECT -280.015 90.525 -279.845 90.695 ;
        RECT -272.855 90.525 -272.685 90.695 ;
        RECT -272.395 90.525 -272.225 90.695 ;
        RECT -271.935 90.525 -271.765 90.695 ;
        RECT -271.475 90.525 -271.305 90.695 ;
        RECT -271.015 90.525 -270.845 90.695 ;
        RECT -270.555 90.525 -270.385 90.695 ;
        RECT -270.095 90.525 -269.925 90.695 ;
        RECT -262.935 90.525 -262.765 90.695 ;
        RECT -262.475 90.525 -262.305 90.695 ;
        RECT -262.015 90.525 -261.845 90.695 ;
        RECT -261.555 90.525 -261.385 90.695 ;
        RECT -261.095 90.525 -260.925 90.695 ;
        RECT -260.635 90.525 -260.465 90.695 ;
        RECT -260.175 90.525 -260.005 90.695 ;
        RECT -253.015 90.525 -252.845 90.695 ;
        RECT -252.555 90.525 -252.385 90.695 ;
        RECT -252.095 90.525 -251.925 90.695 ;
        RECT -251.635 90.525 -251.465 90.695 ;
        RECT -251.175 90.525 -251.005 90.695 ;
        RECT -250.715 90.525 -250.545 90.695 ;
        RECT -250.255 90.525 -250.085 90.695 ;
        RECT -243.095 90.525 -242.925 90.695 ;
        RECT -242.635 90.525 -242.465 90.695 ;
        RECT -242.175 90.525 -242.005 90.695 ;
        RECT -241.715 90.525 -241.545 90.695 ;
        RECT -241.255 90.525 -241.085 90.695 ;
        RECT -240.795 90.525 -240.625 90.695 ;
        RECT -240.335 90.525 -240.165 90.695 ;
        RECT -233.175 90.525 -233.005 90.695 ;
        RECT -232.715 90.525 -232.545 90.695 ;
        RECT -232.255 90.525 -232.085 90.695 ;
        RECT -231.795 90.525 -231.625 90.695 ;
        RECT -231.335 90.525 -231.165 90.695 ;
        RECT -230.875 90.525 -230.705 90.695 ;
        RECT -230.415 90.525 -230.245 90.695 ;
        RECT -223.255 90.525 -223.085 90.695 ;
        RECT -222.795 90.525 -222.625 90.695 ;
        RECT -222.335 90.525 -222.165 90.695 ;
        RECT -221.875 90.525 -221.705 90.695 ;
        RECT -221.415 90.525 -221.245 90.695 ;
        RECT -220.955 90.525 -220.785 90.695 ;
        RECT -220.495 90.525 -220.325 90.695 ;
        RECT -213.335 90.525 -213.165 90.695 ;
        RECT -212.875 90.525 -212.705 90.695 ;
        RECT -212.415 90.525 -212.245 90.695 ;
        RECT -211.955 90.525 -211.785 90.695 ;
        RECT -211.495 90.525 -211.325 90.695 ;
        RECT -211.035 90.525 -210.865 90.695 ;
        RECT -210.575 90.525 -210.405 90.695 ;
        RECT -203.415 90.525 -203.245 90.695 ;
        RECT -202.955 90.525 -202.785 90.695 ;
        RECT -202.495 90.525 -202.325 90.695 ;
        RECT -202.035 90.525 -201.865 90.695 ;
        RECT -201.575 90.525 -201.405 90.695 ;
        RECT -201.115 90.525 -200.945 90.695 ;
        RECT -200.655 90.525 -200.485 90.695 ;
        RECT -193.495 90.525 -193.325 90.695 ;
        RECT -193.035 90.525 -192.865 90.695 ;
        RECT -192.575 90.525 -192.405 90.695 ;
        RECT -192.115 90.525 -191.945 90.695 ;
        RECT -191.655 90.525 -191.485 90.695 ;
        RECT -191.195 90.525 -191.025 90.695 ;
        RECT -190.735 90.525 -190.565 90.695 ;
        RECT -183.575 90.525 -183.405 90.695 ;
        RECT -183.115 90.525 -182.945 90.695 ;
        RECT -182.655 90.525 -182.485 90.695 ;
        RECT -182.195 90.525 -182.025 90.695 ;
        RECT -181.735 90.525 -181.565 90.695 ;
        RECT -181.275 90.525 -181.105 90.695 ;
        RECT -180.815 90.525 -180.645 90.695 ;
        RECT -173.655 90.525 -173.485 90.695 ;
        RECT -173.195 90.525 -173.025 90.695 ;
        RECT -172.735 90.525 -172.565 90.695 ;
        RECT -172.275 90.525 -172.105 90.695 ;
        RECT -171.815 90.525 -171.645 90.695 ;
        RECT -171.355 90.525 -171.185 90.695 ;
        RECT -170.895 90.525 -170.725 90.695 ;
        RECT -163.735 90.525 -163.565 90.695 ;
        RECT -163.275 90.525 -163.105 90.695 ;
        RECT -162.815 90.525 -162.645 90.695 ;
        RECT -162.355 90.525 -162.185 90.695 ;
        RECT -161.895 90.525 -161.725 90.695 ;
        RECT -161.435 90.525 -161.265 90.695 ;
        RECT -160.975 90.525 -160.805 90.695 ;
        RECT -153.815 90.525 -153.645 90.695 ;
        RECT -153.355 90.525 -153.185 90.695 ;
        RECT -152.895 90.525 -152.725 90.695 ;
        RECT -152.435 90.525 -152.265 90.695 ;
        RECT -151.975 90.525 -151.805 90.695 ;
        RECT -151.515 90.525 -151.345 90.695 ;
        RECT -151.055 90.525 -150.885 90.695 ;
        RECT -143.895 90.525 -143.725 90.695 ;
        RECT -143.435 90.525 -143.265 90.695 ;
        RECT -142.975 90.525 -142.805 90.695 ;
        RECT -142.515 90.525 -142.345 90.695 ;
        RECT -142.055 90.525 -141.885 90.695 ;
        RECT -141.595 90.525 -141.425 90.695 ;
        RECT -141.135 90.525 -140.965 90.695 ;
        RECT -133.975 90.525 -133.805 90.695 ;
        RECT -133.515 90.525 -133.345 90.695 ;
        RECT -133.055 90.525 -132.885 90.695 ;
        RECT -132.595 90.525 -132.425 90.695 ;
        RECT -132.135 90.525 -131.965 90.695 ;
        RECT -131.675 90.525 -131.505 90.695 ;
        RECT -131.215 90.525 -131.045 90.695 ;
        RECT -124.055 90.525 -123.885 90.695 ;
        RECT -123.595 90.525 -123.425 90.695 ;
        RECT -123.135 90.525 -122.965 90.695 ;
        RECT -122.675 90.525 -122.505 90.695 ;
        RECT -122.215 90.525 -122.045 90.695 ;
        RECT -121.755 90.525 -121.585 90.695 ;
        RECT -121.295 90.525 -121.125 90.695 ;
        RECT -114.135 90.525 -113.965 90.695 ;
        RECT -113.675 90.525 -113.505 90.695 ;
        RECT -113.215 90.525 -113.045 90.695 ;
        RECT -112.755 90.525 -112.585 90.695 ;
        RECT -112.295 90.525 -112.125 90.695 ;
        RECT -111.835 90.525 -111.665 90.695 ;
        RECT -111.375 90.525 -111.205 90.695 ;
        RECT -104.215 90.525 -104.045 90.695 ;
        RECT -103.755 90.525 -103.585 90.695 ;
        RECT -103.295 90.525 -103.125 90.695 ;
        RECT -102.835 90.525 -102.665 90.695 ;
        RECT -102.375 90.525 -102.205 90.695 ;
        RECT -101.915 90.525 -101.745 90.695 ;
        RECT -101.455 90.525 -101.285 90.695 ;
        RECT -94.295 90.525 -94.125 90.695 ;
        RECT -93.835 90.525 -93.665 90.695 ;
        RECT -93.375 90.525 -93.205 90.695 ;
        RECT -92.915 90.525 -92.745 90.695 ;
        RECT -92.455 90.525 -92.285 90.695 ;
        RECT -91.995 90.525 -91.825 90.695 ;
        RECT -91.535 90.525 -91.365 90.695 ;
        RECT -84.375 90.525 -84.205 90.695 ;
        RECT -83.915 90.525 -83.745 90.695 ;
        RECT -83.455 90.525 -83.285 90.695 ;
        RECT -82.995 90.525 -82.825 90.695 ;
        RECT -82.535 90.525 -82.365 90.695 ;
        RECT -82.075 90.525 -81.905 90.695 ;
        RECT -81.615 90.525 -81.445 90.695 ;
        RECT -74.455 90.525 -74.285 90.695 ;
        RECT -73.995 90.525 -73.825 90.695 ;
        RECT -73.535 90.525 -73.365 90.695 ;
        RECT -73.075 90.525 -72.905 90.695 ;
        RECT -72.615 90.525 -72.445 90.695 ;
        RECT -72.155 90.525 -71.985 90.695 ;
        RECT -71.695 90.525 -71.525 90.695 ;
        RECT -64.535 90.525 -64.365 90.695 ;
        RECT -64.075 90.525 -63.905 90.695 ;
        RECT -63.615 90.525 -63.445 90.695 ;
        RECT -63.155 90.525 -62.985 90.695 ;
        RECT -62.695 90.525 -62.525 90.695 ;
        RECT -62.235 90.525 -62.065 90.695 ;
        RECT -61.775 90.525 -61.605 90.695 ;
        RECT -54.615 90.525 -54.445 90.695 ;
        RECT -54.155 90.525 -53.985 90.695 ;
        RECT -53.695 90.525 -53.525 90.695 ;
        RECT -53.235 90.525 -53.065 90.695 ;
        RECT -52.775 90.525 -52.605 90.695 ;
        RECT -52.315 90.525 -52.145 90.695 ;
        RECT -51.855 90.525 -51.685 90.695 ;
        RECT -44.695 90.525 -44.525 90.695 ;
        RECT -44.235 90.525 -44.065 90.695 ;
        RECT -43.775 90.525 -43.605 90.695 ;
        RECT -43.315 90.525 -43.145 90.695 ;
        RECT -42.855 90.525 -42.685 90.695 ;
        RECT -42.395 90.525 -42.225 90.695 ;
        RECT -41.935 90.525 -41.765 90.695 ;
        RECT -34.775 90.525 -34.605 90.695 ;
        RECT -34.315 90.525 -34.145 90.695 ;
        RECT -33.855 90.525 -33.685 90.695 ;
        RECT -33.395 90.525 -33.225 90.695 ;
        RECT -32.935 90.525 -32.765 90.695 ;
        RECT -32.475 90.525 -32.305 90.695 ;
        RECT -32.015 90.525 -31.845 90.695 ;
        RECT -24.855 90.525 -24.685 90.695 ;
        RECT -24.395 90.525 -24.225 90.695 ;
        RECT -23.935 90.525 -23.765 90.695 ;
        RECT -23.475 90.525 -23.305 90.695 ;
        RECT -23.015 90.525 -22.845 90.695 ;
        RECT -22.555 90.525 -22.385 90.695 ;
        RECT -22.095 90.525 -21.925 90.695 ;
        RECT -14.935 90.525 -14.765 90.695 ;
        RECT -14.475 90.525 -14.305 90.695 ;
        RECT -14.015 90.525 -13.845 90.695 ;
        RECT -13.555 90.525 -13.385 90.695 ;
        RECT -13.095 90.525 -12.925 90.695 ;
        RECT -12.635 90.525 -12.465 90.695 ;
        RECT -12.175 90.525 -12.005 90.695 ;
        RECT -5.015 90.525 -4.845 90.695 ;
        RECT -4.555 90.525 -4.385 90.695 ;
        RECT -4.095 90.525 -3.925 90.695 ;
        RECT -3.635 90.525 -3.465 90.695 ;
        RECT -3.175 90.525 -3.005 90.695 ;
        RECT -2.715 90.525 -2.545 90.695 ;
        RECT -2.255 90.525 -2.085 90.695 ;
        RECT 4.905 90.525 5.075 90.695 ;
        RECT 5.365 90.525 5.535 90.695 ;
        RECT 5.825 90.525 5.995 90.695 ;
        RECT 6.285 90.525 6.455 90.695 ;
        RECT 6.745 90.525 6.915 90.695 ;
        RECT 7.205 90.525 7.375 90.695 ;
        RECT 7.665 90.525 7.835 90.695 ;
        RECT 14.825 90.525 14.995 90.695 ;
        RECT 15.285 90.525 15.455 90.695 ;
        RECT 15.745 90.525 15.915 90.695 ;
        RECT 16.205 90.525 16.375 90.695 ;
        RECT 16.665 90.525 16.835 90.695 ;
        RECT 17.125 90.525 17.295 90.695 ;
        RECT 17.585 90.525 17.755 90.695 ;
        RECT 24.745 90.525 24.915 90.695 ;
        RECT 25.205 90.525 25.375 90.695 ;
        RECT 25.665 90.525 25.835 90.695 ;
        RECT 26.125 90.525 26.295 90.695 ;
        RECT -286.825 89.865 -286.655 90.035 ;
        RECT -286.355 89.940 -286.185 90.110 ;
        RECT -286.825 89.405 -286.655 89.575 ;
        RECT -286.825 88.945 -286.655 89.115 ;
        RECT -285.885 89.865 -285.715 90.035 ;
        RECT -276.905 89.865 -276.735 90.035 ;
        RECT -276.435 89.940 -276.265 90.110 ;
        RECT -285.885 89.405 -285.715 89.575 ;
        RECT -276.905 89.405 -276.735 89.575 ;
        RECT -285.885 88.945 -285.715 89.115 ;
        RECT -276.905 88.945 -276.735 89.115 ;
        RECT -275.965 89.865 -275.795 90.035 ;
        RECT -266.985 89.865 -266.815 90.035 ;
        RECT -266.515 89.940 -266.345 90.110 ;
        RECT -275.965 89.405 -275.795 89.575 ;
        RECT -266.985 89.405 -266.815 89.575 ;
        RECT -275.965 88.945 -275.795 89.115 ;
        RECT -266.985 88.945 -266.815 89.115 ;
        RECT -266.045 89.865 -265.875 90.035 ;
        RECT -257.065 89.865 -256.895 90.035 ;
        RECT -256.595 89.940 -256.425 90.110 ;
        RECT -266.045 89.405 -265.875 89.575 ;
        RECT -257.065 89.405 -256.895 89.575 ;
        RECT -266.045 88.945 -265.875 89.115 ;
        RECT -257.065 88.945 -256.895 89.115 ;
        RECT -256.125 89.865 -255.955 90.035 ;
        RECT -247.145 89.865 -246.975 90.035 ;
        RECT -246.675 89.940 -246.505 90.110 ;
        RECT -256.125 89.405 -255.955 89.575 ;
        RECT -247.145 89.405 -246.975 89.575 ;
        RECT -256.125 88.945 -255.955 89.115 ;
        RECT -247.145 88.945 -246.975 89.115 ;
        RECT -246.205 89.865 -246.035 90.035 ;
        RECT -237.225 89.865 -237.055 90.035 ;
        RECT -236.755 89.940 -236.585 90.110 ;
        RECT -246.205 89.405 -246.035 89.575 ;
        RECT -237.225 89.405 -237.055 89.575 ;
        RECT -246.205 88.945 -246.035 89.115 ;
        RECT -237.225 88.945 -237.055 89.115 ;
        RECT -236.285 89.865 -236.115 90.035 ;
        RECT -227.305 89.865 -227.135 90.035 ;
        RECT -226.835 89.940 -226.665 90.110 ;
        RECT -236.285 89.405 -236.115 89.575 ;
        RECT -227.305 89.405 -227.135 89.575 ;
        RECT -236.285 88.945 -236.115 89.115 ;
        RECT -227.305 88.945 -227.135 89.115 ;
        RECT -226.365 89.865 -226.195 90.035 ;
        RECT -217.385 89.865 -217.215 90.035 ;
        RECT -216.915 89.940 -216.745 90.110 ;
        RECT -226.365 89.405 -226.195 89.575 ;
        RECT -217.385 89.405 -217.215 89.575 ;
        RECT -226.365 88.945 -226.195 89.115 ;
        RECT -217.385 88.945 -217.215 89.115 ;
        RECT -216.445 89.865 -216.275 90.035 ;
        RECT -207.465 89.865 -207.295 90.035 ;
        RECT -206.995 89.940 -206.825 90.110 ;
        RECT -216.445 89.405 -216.275 89.575 ;
        RECT -207.465 89.405 -207.295 89.575 ;
        RECT -216.445 88.945 -216.275 89.115 ;
        RECT -207.465 88.945 -207.295 89.115 ;
        RECT -206.525 89.865 -206.355 90.035 ;
        RECT -197.545 89.865 -197.375 90.035 ;
        RECT -197.075 89.940 -196.905 90.110 ;
        RECT -206.525 89.405 -206.355 89.575 ;
        RECT -197.545 89.405 -197.375 89.575 ;
        RECT -206.525 88.945 -206.355 89.115 ;
        RECT -197.545 88.945 -197.375 89.115 ;
        RECT -196.605 89.865 -196.435 90.035 ;
        RECT -187.625 89.865 -187.455 90.035 ;
        RECT -187.155 89.940 -186.985 90.110 ;
        RECT -196.605 89.405 -196.435 89.575 ;
        RECT -187.625 89.405 -187.455 89.575 ;
        RECT -196.605 88.945 -196.435 89.115 ;
        RECT -187.625 88.945 -187.455 89.115 ;
        RECT -186.685 89.865 -186.515 90.035 ;
        RECT -177.705 89.865 -177.535 90.035 ;
        RECT -177.235 89.940 -177.065 90.110 ;
        RECT -186.685 89.405 -186.515 89.575 ;
        RECT -177.705 89.405 -177.535 89.575 ;
        RECT -186.685 88.945 -186.515 89.115 ;
        RECT -177.705 88.945 -177.535 89.115 ;
        RECT -176.765 89.865 -176.595 90.035 ;
        RECT -167.785 89.865 -167.615 90.035 ;
        RECT -167.315 89.940 -167.145 90.110 ;
        RECT -176.765 89.405 -176.595 89.575 ;
        RECT -167.785 89.405 -167.615 89.575 ;
        RECT -176.765 88.945 -176.595 89.115 ;
        RECT -167.785 88.945 -167.615 89.115 ;
        RECT -166.845 89.865 -166.675 90.035 ;
        RECT -157.865 89.865 -157.695 90.035 ;
        RECT -157.395 89.940 -157.225 90.110 ;
        RECT -166.845 89.405 -166.675 89.575 ;
        RECT -157.865 89.405 -157.695 89.575 ;
        RECT -166.845 88.945 -166.675 89.115 ;
        RECT -157.865 88.945 -157.695 89.115 ;
        RECT -156.925 89.865 -156.755 90.035 ;
        RECT -147.945 89.865 -147.775 90.035 ;
        RECT -147.475 89.940 -147.305 90.110 ;
        RECT -156.925 89.405 -156.755 89.575 ;
        RECT -147.945 89.405 -147.775 89.575 ;
        RECT -156.925 88.945 -156.755 89.115 ;
        RECT -147.945 88.945 -147.775 89.115 ;
        RECT -147.005 89.865 -146.835 90.035 ;
        RECT -138.025 89.865 -137.855 90.035 ;
        RECT -137.555 89.940 -137.385 90.110 ;
        RECT -147.005 89.405 -146.835 89.575 ;
        RECT -138.025 89.405 -137.855 89.575 ;
        RECT -147.005 88.945 -146.835 89.115 ;
        RECT -138.025 88.945 -137.855 89.115 ;
        RECT -137.085 89.865 -136.915 90.035 ;
        RECT -128.105 89.865 -127.935 90.035 ;
        RECT -127.635 89.940 -127.465 90.110 ;
        RECT -137.085 89.405 -136.915 89.575 ;
        RECT -128.105 89.405 -127.935 89.575 ;
        RECT -137.085 88.945 -136.915 89.115 ;
        RECT -128.105 88.945 -127.935 89.115 ;
        RECT -127.165 89.865 -126.995 90.035 ;
        RECT -118.185 89.865 -118.015 90.035 ;
        RECT -117.715 89.940 -117.545 90.110 ;
        RECT -127.165 89.405 -126.995 89.575 ;
        RECT -118.185 89.405 -118.015 89.575 ;
        RECT -127.165 88.945 -126.995 89.115 ;
        RECT -118.185 88.945 -118.015 89.115 ;
        RECT -117.245 89.865 -117.075 90.035 ;
        RECT -108.265 89.865 -108.095 90.035 ;
        RECT -107.795 89.940 -107.625 90.110 ;
        RECT -117.245 89.405 -117.075 89.575 ;
        RECT -108.265 89.405 -108.095 89.575 ;
        RECT -117.245 88.945 -117.075 89.115 ;
        RECT -108.265 88.945 -108.095 89.115 ;
        RECT -107.325 89.865 -107.155 90.035 ;
        RECT -98.345 89.865 -98.175 90.035 ;
        RECT -97.875 89.940 -97.705 90.110 ;
        RECT -107.325 89.405 -107.155 89.575 ;
        RECT -98.345 89.405 -98.175 89.575 ;
        RECT -107.325 88.945 -107.155 89.115 ;
        RECT -98.345 88.945 -98.175 89.115 ;
        RECT -97.405 89.865 -97.235 90.035 ;
        RECT -88.425 89.865 -88.255 90.035 ;
        RECT -87.955 89.940 -87.785 90.110 ;
        RECT -97.405 89.405 -97.235 89.575 ;
        RECT -88.425 89.405 -88.255 89.575 ;
        RECT -97.405 88.945 -97.235 89.115 ;
        RECT -88.425 88.945 -88.255 89.115 ;
        RECT -87.485 89.865 -87.315 90.035 ;
        RECT -78.505 89.865 -78.335 90.035 ;
        RECT -78.035 89.940 -77.865 90.110 ;
        RECT -87.485 89.405 -87.315 89.575 ;
        RECT -78.505 89.405 -78.335 89.575 ;
        RECT -87.485 88.945 -87.315 89.115 ;
        RECT -78.505 88.945 -78.335 89.115 ;
        RECT -77.565 89.865 -77.395 90.035 ;
        RECT -68.585 89.865 -68.415 90.035 ;
        RECT -68.115 89.940 -67.945 90.110 ;
        RECT -77.565 89.405 -77.395 89.575 ;
        RECT -68.585 89.405 -68.415 89.575 ;
        RECT -77.565 88.945 -77.395 89.115 ;
        RECT -68.585 88.945 -68.415 89.115 ;
        RECT -67.645 89.865 -67.475 90.035 ;
        RECT -58.665 89.865 -58.495 90.035 ;
        RECT -58.195 89.940 -58.025 90.110 ;
        RECT -67.645 89.405 -67.475 89.575 ;
        RECT -58.665 89.405 -58.495 89.575 ;
        RECT -67.645 88.945 -67.475 89.115 ;
        RECT -58.665 88.945 -58.495 89.115 ;
        RECT -57.725 89.865 -57.555 90.035 ;
        RECT -48.745 89.865 -48.575 90.035 ;
        RECT -48.275 89.940 -48.105 90.110 ;
        RECT -57.725 89.405 -57.555 89.575 ;
        RECT -48.745 89.405 -48.575 89.575 ;
        RECT -57.725 88.945 -57.555 89.115 ;
        RECT -48.745 88.945 -48.575 89.115 ;
        RECT -47.805 89.865 -47.635 90.035 ;
        RECT -38.825 89.865 -38.655 90.035 ;
        RECT -38.355 89.940 -38.185 90.110 ;
        RECT -47.805 89.405 -47.635 89.575 ;
        RECT -38.825 89.405 -38.655 89.575 ;
        RECT -47.805 88.945 -47.635 89.115 ;
        RECT -38.825 88.945 -38.655 89.115 ;
        RECT -37.885 89.865 -37.715 90.035 ;
        RECT -28.905 89.865 -28.735 90.035 ;
        RECT -28.435 89.940 -28.265 90.110 ;
        RECT -37.885 89.405 -37.715 89.575 ;
        RECT -28.905 89.405 -28.735 89.575 ;
        RECT -37.885 88.945 -37.715 89.115 ;
        RECT -28.905 88.945 -28.735 89.115 ;
        RECT -27.965 89.865 -27.795 90.035 ;
        RECT -18.985 89.865 -18.815 90.035 ;
        RECT -18.515 89.940 -18.345 90.110 ;
        RECT -27.965 89.405 -27.795 89.575 ;
        RECT -18.985 89.405 -18.815 89.575 ;
        RECT -27.965 88.945 -27.795 89.115 ;
        RECT -18.985 88.945 -18.815 89.115 ;
        RECT -18.045 89.865 -17.875 90.035 ;
        RECT -9.065 89.865 -8.895 90.035 ;
        RECT -8.595 89.940 -8.425 90.110 ;
        RECT -18.045 89.405 -17.875 89.575 ;
        RECT -9.065 89.405 -8.895 89.575 ;
        RECT -18.045 88.945 -17.875 89.115 ;
        RECT -9.065 88.945 -8.895 89.115 ;
        RECT -8.125 89.865 -7.955 90.035 ;
        RECT 0.855 89.865 1.025 90.035 ;
        RECT 1.325 89.940 1.495 90.110 ;
        RECT -8.125 89.405 -7.955 89.575 ;
        RECT 0.855 89.405 1.025 89.575 ;
        RECT -8.125 88.945 -7.955 89.115 ;
        RECT 0.855 88.945 1.025 89.115 ;
        RECT 1.795 89.865 1.965 90.035 ;
        RECT 10.775 89.865 10.945 90.035 ;
        RECT 11.245 89.940 11.415 90.110 ;
        RECT 1.795 89.405 1.965 89.575 ;
        RECT 10.775 89.405 10.945 89.575 ;
        RECT 1.795 88.945 1.965 89.115 ;
        RECT 10.775 88.945 10.945 89.115 ;
        RECT 11.715 89.865 11.885 90.035 ;
        RECT 20.695 89.865 20.865 90.035 ;
        RECT 21.165 89.940 21.335 90.110 ;
        RECT 11.715 89.405 11.885 89.575 ;
        RECT 20.695 89.405 20.865 89.575 ;
        RECT 11.715 88.945 11.885 89.115 ;
        RECT 20.695 88.945 20.865 89.115 ;
        RECT 21.635 89.865 21.805 90.035 ;
        RECT 21.635 89.405 21.805 89.575 ;
        RECT 21.635 88.945 21.805 89.115 ;
      LAYER met1 ;
        RECT -281.540 95.140 -281.080 95.145 ;
        RECT -271.620 95.140 -271.160 95.145 ;
        RECT -261.700 95.140 -261.240 95.145 ;
        RECT -251.780 95.140 -251.320 95.145 ;
        RECT -241.860 95.140 -241.400 95.145 ;
        RECT -231.940 95.140 -231.480 95.145 ;
        RECT -222.020 95.140 -221.560 95.145 ;
        RECT -212.100 95.140 -211.640 95.145 ;
        RECT -202.180 95.140 -201.720 95.145 ;
        RECT -192.260 95.140 -191.800 95.145 ;
        RECT -182.340 95.140 -181.880 95.145 ;
        RECT -172.420 95.140 -171.960 95.145 ;
        RECT -162.500 95.140 -162.040 95.145 ;
        RECT -152.580 95.140 -152.120 95.145 ;
        RECT -142.660 95.140 -142.200 95.145 ;
        RECT -132.740 95.140 -132.280 95.145 ;
        RECT -122.820 95.140 -122.360 95.145 ;
        RECT -112.900 95.140 -112.440 95.145 ;
        RECT -102.980 95.140 -102.520 95.145 ;
        RECT -93.060 95.140 -92.600 95.145 ;
        RECT -83.140 95.140 -82.680 95.145 ;
        RECT -73.220 95.140 -72.760 95.145 ;
        RECT -63.300 95.140 -62.840 95.145 ;
        RECT -53.380 95.140 -52.920 95.145 ;
        RECT -43.460 95.140 -43.000 95.145 ;
        RECT -33.540 95.140 -33.080 95.145 ;
        RECT -23.620 95.140 -23.160 95.145 ;
        RECT -13.700 95.140 -13.240 95.145 ;
        RECT -3.780 95.140 -3.320 95.145 ;
        RECT 6.140 95.140 6.600 95.145 ;
        RECT 16.060 95.140 16.520 95.145 ;
        RECT 25.980 95.140 26.440 95.145 ;
        RECT -282.020 93.760 -280.600 95.140 ;
        RECT -272.100 93.760 -270.680 95.140 ;
        RECT -262.180 93.760 -260.760 95.140 ;
        RECT -252.260 93.760 -250.840 95.140 ;
        RECT -242.340 93.760 -240.920 95.140 ;
        RECT -232.420 93.760 -231.000 95.140 ;
        RECT -222.500 93.760 -221.080 95.140 ;
        RECT -212.580 93.760 -211.160 95.140 ;
        RECT -202.660 93.760 -201.240 95.140 ;
        RECT -192.740 93.760 -191.320 95.140 ;
        RECT -182.820 93.760 -181.400 95.140 ;
        RECT -172.900 93.760 -171.480 95.140 ;
        RECT -162.980 93.760 -161.560 95.140 ;
        RECT -153.060 93.760 -151.640 95.140 ;
        RECT -143.140 93.760 -141.720 95.140 ;
        RECT -133.220 93.760 -131.800 95.140 ;
        RECT -123.300 93.760 -121.880 95.140 ;
        RECT -113.380 93.760 -111.960 95.140 ;
        RECT -103.460 93.760 -102.040 95.140 ;
        RECT -93.540 93.760 -92.120 95.140 ;
        RECT -83.620 93.760 -82.200 95.140 ;
        RECT -73.700 93.760 -72.280 95.140 ;
        RECT -63.780 93.760 -62.360 95.140 ;
        RECT -53.860 93.760 -52.440 95.140 ;
        RECT -43.940 93.760 -42.520 95.140 ;
        RECT -34.020 93.760 -32.600 95.140 ;
        RECT -24.100 93.760 -22.680 95.140 ;
        RECT -14.180 93.760 -12.760 95.140 ;
        RECT -4.260 93.760 -2.840 95.140 ;
        RECT 5.660 93.760 7.080 95.140 ;
        RECT 15.580 93.760 17.000 95.140 ;
        RECT 25.500 93.760 26.440 95.140 ;
        RECT -287.880 93.090 -284.660 93.570 ;
        RECT -277.960 93.090 -274.740 93.570 ;
        RECT -268.040 93.090 -264.820 93.570 ;
        RECT -258.120 93.090 -254.900 93.570 ;
        RECT -248.200 93.090 -244.980 93.570 ;
        RECT -238.280 93.090 -235.060 93.570 ;
        RECT -228.360 93.090 -225.140 93.570 ;
        RECT -218.440 93.090 -215.220 93.570 ;
        RECT -208.520 93.090 -205.300 93.570 ;
        RECT -198.600 93.090 -195.380 93.570 ;
        RECT -188.680 93.090 -185.460 93.570 ;
        RECT -178.760 93.090 -175.540 93.570 ;
        RECT -168.840 93.090 -165.620 93.570 ;
        RECT -158.920 93.090 -155.700 93.570 ;
        RECT -149.000 93.090 -145.780 93.570 ;
        RECT -139.080 93.090 -135.860 93.570 ;
        RECT -129.160 93.090 -125.940 93.570 ;
        RECT -119.240 93.090 -116.020 93.570 ;
        RECT -109.320 93.090 -106.100 93.570 ;
        RECT -99.400 93.090 -96.180 93.570 ;
        RECT -89.480 93.090 -86.260 93.570 ;
        RECT -79.560 93.090 -76.340 93.570 ;
        RECT -69.640 93.090 -66.420 93.570 ;
        RECT -59.720 93.090 -56.500 93.570 ;
        RECT -49.800 93.090 -46.580 93.570 ;
        RECT -39.880 93.090 -36.660 93.570 ;
        RECT -29.960 93.090 -26.740 93.570 ;
        RECT -20.040 93.090 -16.820 93.570 ;
        RECT -10.120 93.090 -6.900 93.570 ;
        RECT -0.200 93.090 3.020 93.570 ;
        RECT 9.720 93.090 12.940 93.570 ;
        RECT 19.640 93.090 22.860 93.570 ;
        RECT -282.920 90.370 -279.700 90.850 ;
        RECT -273.000 90.370 -269.780 90.850 ;
        RECT -263.080 90.370 -259.860 90.850 ;
        RECT -253.160 90.370 -249.940 90.850 ;
        RECT -243.240 90.370 -240.020 90.850 ;
        RECT -233.320 90.370 -230.100 90.850 ;
        RECT -223.400 90.370 -220.180 90.850 ;
        RECT -213.480 90.370 -210.260 90.850 ;
        RECT -203.560 90.370 -200.340 90.850 ;
        RECT -193.640 90.370 -190.420 90.850 ;
        RECT -183.720 90.370 -180.500 90.850 ;
        RECT -173.800 90.370 -170.580 90.850 ;
        RECT -163.880 90.370 -160.660 90.850 ;
        RECT -153.960 90.370 -150.740 90.850 ;
        RECT -144.040 90.370 -140.820 90.850 ;
        RECT -134.120 90.370 -130.900 90.850 ;
        RECT -124.200 90.370 -120.980 90.850 ;
        RECT -114.280 90.370 -111.060 90.850 ;
        RECT -104.360 90.370 -101.140 90.850 ;
        RECT -94.440 90.370 -91.220 90.850 ;
        RECT -84.520 90.370 -81.300 90.850 ;
        RECT -74.600 90.370 -71.380 90.850 ;
        RECT -64.680 90.370 -61.460 90.850 ;
        RECT -54.760 90.370 -51.540 90.850 ;
        RECT -44.840 90.370 -41.620 90.850 ;
        RECT -34.920 90.370 -31.700 90.850 ;
        RECT -25.000 90.370 -21.780 90.850 ;
        RECT -15.080 90.370 -11.860 90.850 ;
        RECT -5.160 90.370 -1.940 90.850 ;
        RECT 4.760 90.370 7.980 90.850 ;
        RECT 14.680 90.370 17.900 90.850 ;
        RECT 24.600 90.370 26.440 90.850 ;
        RECT -286.980 88.800 -285.560 90.180 ;
        RECT -277.060 88.800 -275.640 90.180 ;
        RECT -267.140 88.800 -265.720 90.180 ;
        RECT -257.220 88.800 -255.800 90.180 ;
        RECT -247.300 88.800 -245.880 90.180 ;
        RECT -237.380 88.800 -235.960 90.180 ;
        RECT -227.460 88.800 -226.040 90.180 ;
        RECT -217.540 88.800 -216.120 90.180 ;
        RECT -207.620 88.800 -206.200 90.180 ;
        RECT -197.700 88.800 -196.280 90.180 ;
        RECT -187.780 88.800 -186.360 90.180 ;
        RECT -177.860 88.800 -176.440 90.180 ;
        RECT -167.940 88.800 -166.520 90.180 ;
        RECT -158.020 88.800 -156.600 90.180 ;
        RECT -148.100 88.800 -146.680 90.180 ;
        RECT -138.180 88.800 -136.760 90.180 ;
        RECT -128.260 88.800 -126.840 90.180 ;
        RECT -118.340 88.800 -116.920 90.180 ;
        RECT -108.420 88.800 -107.000 90.180 ;
        RECT -98.500 88.800 -97.080 90.180 ;
        RECT -88.580 88.800 -87.160 90.180 ;
        RECT -78.660 88.800 -77.240 90.180 ;
        RECT -68.740 88.800 -67.320 90.180 ;
        RECT -58.820 88.800 -57.400 90.180 ;
        RECT -48.900 88.800 -47.480 90.180 ;
        RECT -38.980 88.800 -37.560 90.180 ;
        RECT -29.060 88.800 -27.640 90.180 ;
        RECT -19.140 88.800 -17.720 90.180 ;
        RECT -9.220 88.800 -7.800 90.180 ;
        RECT 0.700 88.800 2.120 90.180 ;
        RECT 10.620 88.800 12.040 90.180 ;
        RECT 20.540 88.800 21.960 90.180 ;
      LAYER via ;
        RECT -281.920 94.780 -281.645 95.045 ;
        RECT -280.980 94.770 -280.705 95.035 ;
        RECT -272.000 95.040 -271.725 95.045 ;
        RECT -272.000 94.780 -271.490 95.040 ;
        RECT -271.760 94.770 -271.490 94.780 ;
        RECT -271.290 95.035 -271.020 95.040 ;
        RECT -271.290 94.770 -270.785 95.035 ;
        RECT -262.080 94.780 -261.805 95.045 ;
        RECT -261.140 94.770 -260.865 95.035 ;
        RECT -252.160 94.780 -251.885 95.045 ;
        RECT -251.220 94.770 -250.945 95.035 ;
        RECT -242.240 94.780 -241.965 95.045 ;
        RECT -241.300 94.770 -241.025 95.035 ;
        RECT -232.320 94.780 -232.045 95.045 ;
        RECT -231.380 94.770 -231.105 95.035 ;
        RECT -222.400 94.780 -222.125 95.045 ;
        RECT -221.460 94.770 -221.185 95.035 ;
        RECT -212.480 94.780 -212.205 95.045 ;
        RECT -211.540 94.770 -211.265 95.035 ;
        RECT -202.560 94.780 -202.285 95.045 ;
        RECT -201.620 94.770 -201.345 95.035 ;
        RECT -192.640 94.780 -192.365 95.045 ;
        RECT -191.700 94.770 -191.425 95.035 ;
        RECT -182.720 94.780 -182.445 95.045 ;
        RECT -181.780 94.770 -181.505 95.035 ;
        RECT -172.800 94.780 -172.525 95.045 ;
        RECT -171.860 94.770 -171.585 95.035 ;
        RECT -162.880 94.780 -162.605 95.045 ;
        RECT -161.940 94.770 -161.665 95.035 ;
        RECT -152.960 94.780 -152.685 95.045 ;
        RECT -152.020 94.770 -151.745 95.035 ;
        RECT -143.040 94.780 -142.765 95.045 ;
        RECT -142.100 94.770 -141.825 95.035 ;
        RECT -133.120 94.780 -132.845 95.045 ;
        RECT -132.180 94.770 -131.905 95.035 ;
        RECT -123.200 94.780 -122.925 95.045 ;
        RECT -122.260 94.770 -121.985 95.035 ;
        RECT -113.280 94.780 -113.005 95.045 ;
        RECT -112.340 94.770 -112.065 95.035 ;
        RECT -103.360 94.780 -103.085 95.045 ;
        RECT -102.420 94.770 -102.145 95.035 ;
        RECT -93.440 94.780 -93.165 95.045 ;
        RECT -92.500 94.770 -92.225 95.035 ;
        RECT -83.520 94.780 -83.245 95.045 ;
        RECT -82.580 94.770 -82.305 95.035 ;
        RECT -73.600 94.780 -73.325 95.045 ;
        RECT -72.660 94.770 -72.385 95.035 ;
        RECT -63.680 94.780 -63.405 95.045 ;
        RECT -62.740 94.770 -62.465 95.035 ;
        RECT -53.760 94.780 -53.485 95.045 ;
        RECT -52.820 94.770 -52.545 95.035 ;
        RECT -43.840 94.780 -43.565 95.045 ;
        RECT -42.900 94.770 -42.625 95.035 ;
        RECT -33.920 94.780 -33.645 95.045 ;
        RECT -32.980 94.770 -32.705 95.035 ;
        RECT -24.000 94.780 -23.725 95.045 ;
        RECT -23.060 94.770 -22.785 95.035 ;
        RECT -14.080 94.780 -13.805 95.045 ;
        RECT -13.140 94.770 -12.865 95.035 ;
        RECT -4.160 94.780 -3.885 95.045 ;
        RECT -3.220 94.770 -2.945 95.035 ;
        RECT 5.760 94.780 6.035 95.045 ;
        RECT 6.700 94.770 6.975 95.035 ;
        RECT 15.680 94.780 15.955 95.045 ;
        RECT 16.620 94.770 16.895 95.035 ;
        RECT 25.600 94.780 25.875 95.045 ;
        RECT -286.640 93.190 -286.365 93.455 ;
        RECT -286.180 93.190 -285.905 93.455 ;
        RECT -276.720 93.190 -276.445 93.455 ;
        RECT -276.260 93.190 -275.985 93.455 ;
        RECT -266.800 93.190 -266.525 93.455 ;
        RECT -266.340 93.190 -266.065 93.455 ;
        RECT -256.880 93.190 -256.605 93.455 ;
        RECT -256.420 93.190 -256.145 93.455 ;
        RECT -246.960 93.190 -246.685 93.455 ;
        RECT -246.500 93.190 -246.225 93.455 ;
        RECT -237.040 93.190 -236.765 93.455 ;
        RECT -236.580 93.190 -236.305 93.455 ;
        RECT -227.120 93.190 -226.845 93.455 ;
        RECT -226.660 93.190 -226.385 93.455 ;
        RECT -217.200 93.190 -216.925 93.455 ;
        RECT -216.740 93.190 -216.465 93.455 ;
        RECT -207.280 93.190 -207.005 93.455 ;
        RECT -206.820 93.190 -206.545 93.455 ;
        RECT -197.360 93.190 -197.085 93.455 ;
        RECT -196.900 93.190 -196.625 93.455 ;
        RECT -187.440 93.190 -187.165 93.455 ;
        RECT -186.980 93.190 -186.705 93.455 ;
        RECT -177.520 93.190 -177.245 93.455 ;
        RECT -177.060 93.190 -176.785 93.455 ;
        RECT -167.600 93.190 -167.325 93.455 ;
        RECT -167.140 93.190 -166.865 93.455 ;
        RECT -157.680 93.190 -157.405 93.455 ;
        RECT -157.220 93.190 -156.945 93.455 ;
        RECT -147.760 93.190 -147.485 93.455 ;
        RECT -147.300 93.190 -147.025 93.455 ;
        RECT -137.840 93.190 -137.565 93.455 ;
        RECT -137.380 93.190 -137.105 93.455 ;
        RECT -127.920 93.190 -127.645 93.455 ;
        RECT -127.460 93.190 -127.185 93.455 ;
        RECT -118.000 93.190 -117.725 93.455 ;
        RECT -117.540 93.190 -117.265 93.455 ;
        RECT -108.080 93.190 -107.805 93.455 ;
        RECT -107.620 93.190 -107.345 93.455 ;
        RECT -98.160 93.190 -97.885 93.455 ;
        RECT -97.700 93.190 -97.425 93.455 ;
        RECT -88.240 93.190 -87.965 93.455 ;
        RECT -87.780 93.190 -87.505 93.455 ;
        RECT -78.320 93.190 -78.045 93.455 ;
        RECT -77.860 93.190 -77.585 93.455 ;
        RECT -68.400 93.190 -68.125 93.455 ;
        RECT -67.940 93.190 -67.665 93.455 ;
        RECT -58.480 93.190 -58.205 93.455 ;
        RECT -58.020 93.190 -57.745 93.455 ;
        RECT -48.560 93.190 -48.285 93.455 ;
        RECT -48.100 93.190 -47.825 93.455 ;
        RECT -38.640 93.190 -38.365 93.455 ;
        RECT -38.180 93.190 -37.905 93.455 ;
        RECT -28.720 93.190 -28.445 93.455 ;
        RECT -28.260 93.190 -27.985 93.455 ;
        RECT -18.800 93.190 -18.525 93.455 ;
        RECT -18.340 93.190 -18.065 93.455 ;
        RECT -8.880 93.190 -8.605 93.455 ;
        RECT -8.420 93.190 -8.145 93.455 ;
        RECT 1.040 93.190 1.315 93.455 ;
        RECT 1.500 93.190 1.775 93.455 ;
        RECT 10.960 93.190 11.235 93.455 ;
        RECT 11.420 93.190 11.695 93.455 ;
        RECT 20.880 93.190 21.155 93.455 ;
        RECT 21.340 93.190 21.615 93.455 ;
        RECT -281.680 90.480 -281.405 90.745 ;
        RECT -281.220 90.480 -280.945 90.745 ;
        RECT -271.760 90.480 -271.485 90.745 ;
        RECT -271.300 90.480 -271.025 90.745 ;
        RECT -261.840 90.480 -261.565 90.745 ;
        RECT -261.380 90.480 -261.105 90.745 ;
        RECT -251.920 90.480 -251.645 90.745 ;
        RECT -251.460 90.480 -251.185 90.745 ;
        RECT -242.000 90.480 -241.725 90.745 ;
        RECT -241.540 90.480 -241.265 90.745 ;
        RECT -232.080 90.480 -231.805 90.745 ;
        RECT -231.620 90.480 -231.345 90.745 ;
        RECT -222.160 90.480 -221.885 90.745 ;
        RECT -221.700 90.480 -221.425 90.745 ;
        RECT -212.240 90.480 -211.965 90.745 ;
        RECT -211.780 90.480 -211.505 90.745 ;
        RECT -202.320 90.480 -202.045 90.745 ;
        RECT -201.860 90.480 -201.585 90.745 ;
        RECT -192.400 90.480 -192.125 90.745 ;
        RECT -191.940 90.480 -191.665 90.745 ;
        RECT -182.480 90.480 -182.205 90.745 ;
        RECT -182.020 90.480 -181.745 90.745 ;
        RECT -172.560 90.480 -172.285 90.745 ;
        RECT -172.100 90.480 -171.825 90.745 ;
        RECT -162.640 90.480 -162.365 90.745 ;
        RECT -162.180 90.480 -161.905 90.745 ;
        RECT -152.720 90.480 -152.445 90.745 ;
        RECT -152.260 90.480 -151.985 90.745 ;
        RECT -142.800 90.480 -142.525 90.745 ;
        RECT -142.340 90.480 -142.065 90.745 ;
        RECT -132.880 90.480 -132.605 90.745 ;
        RECT -132.420 90.480 -132.145 90.745 ;
        RECT -122.960 90.480 -122.685 90.745 ;
        RECT -122.500 90.480 -122.225 90.745 ;
        RECT -113.040 90.480 -112.765 90.745 ;
        RECT -112.580 90.480 -112.305 90.745 ;
        RECT -103.120 90.480 -102.845 90.745 ;
        RECT -102.660 90.480 -102.385 90.745 ;
        RECT -93.200 90.480 -92.925 90.745 ;
        RECT -92.740 90.480 -92.465 90.745 ;
        RECT -83.280 90.480 -83.005 90.745 ;
        RECT -82.820 90.480 -82.545 90.745 ;
        RECT -73.360 90.480 -73.085 90.745 ;
        RECT -72.900 90.480 -72.625 90.745 ;
        RECT -63.440 90.480 -63.165 90.745 ;
        RECT -62.980 90.480 -62.705 90.745 ;
        RECT -53.520 90.480 -53.245 90.745 ;
        RECT -53.060 90.480 -52.785 90.745 ;
        RECT -43.600 90.480 -43.325 90.745 ;
        RECT -43.140 90.480 -42.865 90.745 ;
        RECT -33.680 90.480 -33.405 90.745 ;
        RECT -33.220 90.480 -32.945 90.745 ;
        RECT -23.760 90.480 -23.485 90.745 ;
        RECT -23.300 90.480 -23.025 90.745 ;
        RECT -13.840 90.480 -13.565 90.745 ;
        RECT -13.380 90.480 -13.105 90.745 ;
        RECT -3.920 90.480 -3.645 90.745 ;
        RECT -3.460 90.480 -3.185 90.745 ;
        RECT 6.000 90.480 6.275 90.745 ;
        RECT 6.460 90.480 6.735 90.745 ;
        RECT 15.920 90.480 16.195 90.745 ;
        RECT 16.380 90.480 16.655 90.745 ;
        RECT 25.840 90.480 26.115 90.745 ;
        RECT -286.870 88.890 -286.595 89.155 ;
        RECT -285.940 88.890 -285.665 89.155 ;
        RECT -276.950 88.890 -276.675 89.155 ;
        RECT -276.020 88.890 -275.745 89.155 ;
        RECT -267.030 88.890 -266.755 89.155 ;
        RECT -266.100 88.890 -265.825 89.155 ;
        RECT -257.110 88.890 -256.835 89.155 ;
        RECT -256.180 88.890 -255.905 89.155 ;
        RECT -247.190 88.890 -246.915 89.155 ;
        RECT -246.260 88.890 -245.985 89.155 ;
        RECT -237.270 88.890 -236.995 89.155 ;
        RECT -236.340 88.890 -236.065 89.155 ;
        RECT -227.350 88.890 -227.075 89.155 ;
        RECT -226.420 88.890 -226.145 89.155 ;
        RECT -217.430 88.890 -217.155 89.155 ;
        RECT -216.500 88.890 -216.225 89.155 ;
        RECT -207.510 88.890 -207.235 89.155 ;
        RECT -206.580 88.890 -206.305 89.155 ;
        RECT -197.590 88.890 -197.315 89.155 ;
        RECT -196.660 88.890 -196.385 89.155 ;
        RECT -187.670 88.890 -187.395 89.155 ;
        RECT -186.740 88.890 -186.465 89.155 ;
        RECT -177.750 88.890 -177.475 89.155 ;
        RECT -176.820 88.890 -176.545 89.155 ;
        RECT -167.830 88.890 -167.555 89.155 ;
        RECT -166.900 88.890 -166.625 89.155 ;
        RECT -157.910 88.890 -157.635 89.155 ;
        RECT -156.980 88.890 -156.705 89.155 ;
        RECT -147.990 88.890 -147.715 89.155 ;
        RECT -147.060 88.890 -146.785 89.155 ;
        RECT -138.070 88.890 -137.795 89.155 ;
        RECT -137.140 88.890 -136.865 89.155 ;
        RECT -128.150 88.890 -127.875 89.155 ;
        RECT -127.220 88.890 -126.945 89.155 ;
        RECT -118.230 88.890 -117.955 89.155 ;
        RECT -117.300 88.890 -117.025 89.155 ;
        RECT -108.310 88.890 -108.035 89.155 ;
        RECT -107.380 88.890 -107.105 89.155 ;
        RECT -98.390 88.890 -98.115 89.155 ;
        RECT -97.460 88.890 -97.185 89.155 ;
        RECT -88.470 88.890 -88.195 89.155 ;
        RECT -87.540 88.890 -87.265 89.155 ;
        RECT -78.550 88.890 -78.275 89.155 ;
        RECT -77.620 88.890 -77.345 89.155 ;
        RECT -68.630 88.890 -68.355 89.155 ;
        RECT -67.700 88.890 -67.425 89.155 ;
        RECT -58.710 88.890 -58.435 89.155 ;
        RECT -57.780 88.890 -57.505 89.155 ;
        RECT -48.790 88.890 -48.515 89.155 ;
        RECT -47.860 88.890 -47.585 89.155 ;
        RECT -38.870 88.890 -38.595 89.155 ;
        RECT -37.940 88.890 -37.665 89.155 ;
        RECT -28.950 88.890 -28.675 89.155 ;
        RECT -28.020 88.890 -27.745 89.155 ;
        RECT -19.030 88.890 -18.755 89.155 ;
        RECT -18.100 88.890 -17.825 89.155 ;
        RECT -9.110 88.890 -8.835 89.155 ;
        RECT -8.180 88.890 -7.905 89.155 ;
        RECT 0.810 88.890 1.085 89.155 ;
        RECT 1.740 88.890 2.015 89.155 ;
        RECT 10.730 88.890 11.005 89.155 ;
        RECT 11.660 88.890 11.935 89.155 ;
        RECT 20.650 88.890 20.925 89.155 ;
        RECT 21.580 88.890 21.855 89.155 ;
      LAYER met2 ;
        RECT -282.020 94.730 -280.600 95.140 ;
        RECT -272.100 94.730 -270.680 95.140 ;
        RECT -262.180 94.730 -260.760 95.140 ;
        RECT -252.260 94.730 -250.840 95.140 ;
        RECT -242.340 94.730 -240.920 95.140 ;
        RECT -232.420 94.730 -231.000 95.140 ;
        RECT -222.500 94.730 -221.080 95.140 ;
        RECT -212.580 94.730 -211.160 95.140 ;
        RECT -202.660 94.730 -201.240 95.140 ;
        RECT -192.740 94.730 -191.320 95.140 ;
        RECT -182.820 94.730 -181.400 95.140 ;
        RECT -172.900 94.730 -171.480 95.140 ;
        RECT -162.980 94.730 -161.560 95.140 ;
        RECT -153.060 94.730 -151.640 95.140 ;
        RECT -143.140 94.730 -141.720 95.140 ;
        RECT -133.220 94.730 -131.800 95.140 ;
        RECT -123.300 94.730 -121.880 95.140 ;
        RECT -113.380 94.730 -111.960 95.140 ;
        RECT -103.460 94.730 -102.040 95.140 ;
        RECT -93.540 94.730 -92.120 95.140 ;
        RECT -83.620 94.730 -82.200 95.140 ;
        RECT -73.700 94.730 -72.280 95.140 ;
        RECT -63.780 94.730 -62.360 95.140 ;
        RECT -53.860 94.730 -52.440 95.140 ;
        RECT -43.940 94.730 -42.520 95.140 ;
        RECT -34.020 94.730 -32.600 95.140 ;
        RECT -24.100 94.730 -22.680 95.140 ;
        RECT -14.180 94.730 -12.760 95.140 ;
        RECT -4.260 94.730 -2.840 95.140 ;
        RECT 5.660 94.730 7.080 95.140 ;
        RECT 15.580 94.730 17.000 95.140 ;
        RECT 25.500 94.730 26.440 95.140 ;
        RECT -272.100 94.360 -270.690 94.730 ;
        RECT -286.870 93.090 -285.670 93.570 ;
        RECT -276.950 93.090 -275.750 93.570 ;
        RECT -267.030 93.090 -265.830 93.570 ;
        RECT -257.110 93.090 -255.910 93.570 ;
        RECT -247.190 93.090 -245.990 93.570 ;
        RECT -237.270 93.090 -236.070 93.570 ;
        RECT -227.350 93.090 -226.150 93.570 ;
        RECT -217.430 93.090 -216.230 93.570 ;
        RECT -207.510 93.090 -206.310 93.570 ;
        RECT -197.590 93.090 -196.390 93.570 ;
        RECT -187.670 93.090 -186.470 93.570 ;
        RECT -177.750 93.090 -176.550 93.570 ;
        RECT -167.830 93.090 -166.630 93.570 ;
        RECT -157.910 93.090 -156.710 93.570 ;
        RECT -147.990 93.090 -146.790 93.570 ;
        RECT -138.070 93.090 -136.870 93.570 ;
        RECT -128.150 93.090 -126.950 93.570 ;
        RECT -118.230 93.090 -117.030 93.570 ;
        RECT -108.310 93.090 -107.110 93.570 ;
        RECT -98.390 93.090 -97.190 93.570 ;
        RECT -88.470 93.090 -87.270 93.570 ;
        RECT -78.550 93.090 -77.350 93.570 ;
        RECT -68.630 93.090 -67.430 93.570 ;
        RECT -58.710 93.090 -57.510 93.570 ;
        RECT -48.790 93.090 -47.590 93.570 ;
        RECT -38.870 93.090 -37.670 93.570 ;
        RECT -28.950 93.090 -27.750 93.570 ;
        RECT -19.030 93.090 -17.830 93.570 ;
        RECT -9.110 93.090 -7.910 93.570 ;
        RECT 0.810 93.090 2.010 93.570 ;
        RECT 10.730 93.090 11.930 93.570 ;
        RECT 20.650 93.090 21.850 93.570 ;
        RECT -281.910 90.370 -280.710 90.850 ;
        RECT -271.990 90.370 -270.790 90.850 ;
        RECT -262.070 90.370 -260.870 90.850 ;
        RECT -252.150 90.370 -250.950 90.850 ;
        RECT -242.230 90.370 -241.030 90.850 ;
        RECT -232.310 90.370 -231.110 90.850 ;
        RECT -222.390 90.370 -221.190 90.850 ;
        RECT -212.470 90.370 -211.270 90.850 ;
        RECT -202.550 90.370 -201.350 90.850 ;
        RECT -192.630 90.370 -191.430 90.850 ;
        RECT -182.710 90.370 -181.510 90.850 ;
        RECT -172.790 90.370 -171.590 90.850 ;
        RECT -162.870 90.370 -161.670 90.850 ;
        RECT -152.950 90.370 -151.750 90.850 ;
        RECT -143.030 90.370 -141.830 90.850 ;
        RECT -133.110 90.370 -131.910 90.850 ;
        RECT -123.190 90.370 -121.990 90.850 ;
        RECT -113.270 90.370 -112.070 90.850 ;
        RECT -103.350 90.370 -102.150 90.850 ;
        RECT -93.430 90.370 -92.230 90.850 ;
        RECT -83.510 90.370 -82.310 90.850 ;
        RECT -73.590 90.370 -72.390 90.850 ;
        RECT -63.670 90.370 -62.470 90.850 ;
        RECT -53.750 90.370 -52.550 90.850 ;
        RECT -43.830 90.370 -42.630 90.850 ;
        RECT -33.910 90.370 -32.710 90.850 ;
        RECT -23.990 90.370 -22.790 90.850 ;
        RECT -14.070 90.370 -12.870 90.850 ;
        RECT -4.150 90.370 -2.950 90.850 ;
        RECT 5.770 90.370 6.970 90.850 ;
        RECT 15.690 90.370 16.890 90.850 ;
        RECT 25.610 90.370 26.440 90.850 ;
        RECT -286.980 88.800 -285.560 89.210 ;
        RECT -277.060 88.800 -275.640 89.210 ;
        RECT -267.140 88.800 -265.720 89.210 ;
        RECT -257.220 88.800 -255.800 89.210 ;
        RECT -247.300 88.800 -245.880 89.210 ;
        RECT -237.380 88.800 -235.960 89.210 ;
        RECT -227.460 88.800 -226.040 89.210 ;
        RECT -217.540 88.800 -216.120 89.210 ;
        RECT -207.620 88.800 -206.200 89.210 ;
        RECT -197.700 88.800 -196.280 89.210 ;
        RECT -187.780 88.800 -186.360 89.210 ;
        RECT -177.860 88.800 -176.440 89.210 ;
        RECT -167.940 88.800 -166.520 89.210 ;
        RECT -158.020 88.800 -156.600 89.210 ;
        RECT -148.100 88.800 -146.680 89.210 ;
        RECT -138.180 88.800 -136.760 89.210 ;
        RECT -128.260 88.800 -126.840 89.210 ;
        RECT -118.340 88.800 -116.920 89.210 ;
        RECT -108.420 88.800 -107.000 89.210 ;
        RECT -98.500 88.800 -97.080 89.210 ;
        RECT -88.580 88.800 -87.160 89.210 ;
        RECT -78.660 88.800 -77.240 89.210 ;
        RECT -68.740 88.800 -67.320 89.210 ;
        RECT -58.820 88.800 -57.400 89.210 ;
        RECT -48.900 88.800 -47.480 89.210 ;
        RECT -38.980 88.800 -37.560 89.210 ;
        RECT -29.060 88.800 -27.640 89.210 ;
        RECT -19.140 88.800 -17.720 89.210 ;
        RECT -9.220 88.800 -7.800 89.210 ;
        RECT 0.700 88.800 2.120 89.210 ;
        RECT 10.620 88.800 12.040 89.210 ;
        RECT 20.540 88.800 21.960 89.210 ;
      LAYER via2 ;
        RECT -281.920 94.770 -281.630 95.050 ;
        RECT -280.990 94.760 -280.700 95.040 ;
        RECT -272.000 94.770 -271.710 95.050 ;
        RECT -271.070 94.760 -270.780 95.040 ;
        RECT -262.080 94.770 -261.790 95.050 ;
        RECT -261.150 94.760 -260.860 95.040 ;
        RECT -252.160 94.770 -251.870 95.050 ;
        RECT -251.230 94.760 -250.940 95.040 ;
        RECT -242.240 94.770 -241.950 95.050 ;
        RECT -241.310 94.760 -241.020 95.040 ;
        RECT -232.320 94.770 -232.030 95.050 ;
        RECT -231.390 94.760 -231.100 95.040 ;
        RECT -222.400 94.770 -222.110 95.050 ;
        RECT -221.470 94.760 -221.180 95.040 ;
        RECT -212.480 94.770 -212.190 95.050 ;
        RECT -211.550 94.760 -211.260 95.040 ;
        RECT -202.560 94.770 -202.270 95.050 ;
        RECT -201.630 94.760 -201.340 95.040 ;
        RECT -192.640 94.770 -192.350 95.050 ;
        RECT -191.710 94.760 -191.420 95.040 ;
        RECT -182.720 94.770 -182.430 95.050 ;
        RECT -181.790 94.760 -181.500 95.040 ;
        RECT -172.800 94.770 -172.510 95.050 ;
        RECT -171.870 94.760 -171.580 95.040 ;
        RECT -162.880 94.770 -162.590 95.050 ;
        RECT -161.950 94.760 -161.660 95.040 ;
        RECT -152.960 94.770 -152.670 95.050 ;
        RECT -152.030 94.760 -151.740 95.040 ;
        RECT -143.040 94.770 -142.750 95.050 ;
        RECT -142.110 94.760 -141.820 95.040 ;
        RECT -133.120 94.770 -132.830 95.050 ;
        RECT -132.190 94.760 -131.900 95.040 ;
        RECT -123.200 94.770 -122.910 95.050 ;
        RECT -122.270 94.760 -121.980 95.040 ;
        RECT -113.280 94.770 -112.990 95.050 ;
        RECT -112.350 94.760 -112.060 95.040 ;
        RECT -103.360 94.770 -103.070 95.050 ;
        RECT -102.430 94.760 -102.140 95.040 ;
        RECT -93.440 94.770 -93.150 95.050 ;
        RECT -92.510 94.760 -92.220 95.040 ;
        RECT -83.520 94.770 -83.230 95.050 ;
        RECT -82.590 94.760 -82.300 95.040 ;
        RECT -73.600 94.770 -73.310 95.050 ;
        RECT -72.670 94.760 -72.380 95.040 ;
        RECT -63.680 94.770 -63.390 95.050 ;
        RECT -62.750 94.760 -62.460 95.040 ;
        RECT -53.760 94.770 -53.470 95.050 ;
        RECT -52.830 94.760 -52.540 95.040 ;
        RECT -43.840 94.770 -43.550 95.050 ;
        RECT -42.910 94.760 -42.620 95.040 ;
        RECT -33.920 94.770 -33.630 95.050 ;
        RECT -32.990 94.760 -32.700 95.040 ;
        RECT -24.000 94.770 -23.710 95.050 ;
        RECT -23.070 94.760 -22.780 95.040 ;
        RECT -14.080 94.770 -13.790 95.050 ;
        RECT -13.150 94.760 -12.860 95.040 ;
        RECT -4.160 94.770 -3.870 95.050 ;
        RECT -3.230 94.760 -2.940 95.040 ;
        RECT 5.760 94.770 6.050 95.050 ;
        RECT 6.690 94.760 6.980 95.040 ;
        RECT 15.680 94.770 15.970 95.050 ;
        RECT 16.610 94.760 16.900 95.040 ;
        RECT 25.600 94.770 25.890 95.050 ;
        RECT -286.580 93.280 -286.290 93.560 ;
        RECT -276.660 93.280 -276.370 93.560 ;
        RECT -266.740 93.280 -266.450 93.560 ;
        RECT -256.820 93.280 -256.530 93.560 ;
        RECT -246.900 93.280 -246.610 93.560 ;
        RECT -236.980 93.280 -236.690 93.560 ;
        RECT -227.060 93.280 -226.770 93.560 ;
        RECT -217.140 93.280 -216.850 93.560 ;
        RECT -207.220 93.280 -206.930 93.560 ;
        RECT -197.300 93.280 -197.010 93.560 ;
        RECT -187.380 93.280 -187.090 93.560 ;
        RECT -177.460 93.280 -177.170 93.560 ;
        RECT -167.540 93.280 -167.250 93.560 ;
        RECT -157.620 93.280 -157.330 93.560 ;
        RECT -147.700 93.280 -147.410 93.560 ;
        RECT -137.780 93.280 -137.490 93.560 ;
        RECT -127.860 93.280 -127.570 93.560 ;
        RECT -117.940 93.280 -117.650 93.560 ;
        RECT -108.020 93.280 -107.730 93.560 ;
        RECT -98.100 93.280 -97.810 93.560 ;
        RECT -88.180 93.280 -87.890 93.560 ;
        RECT -78.260 93.280 -77.970 93.560 ;
        RECT -68.340 93.280 -68.050 93.560 ;
        RECT -58.420 93.280 -58.130 93.560 ;
        RECT -48.500 93.280 -48.210 93.560 ;
        RECT -38.580 93.280 -38.290 93.560 ;
        RECT -28.660 93.280 -28.370 93.560 ;
        RECT -18.740 93.280 -18.450 93.560 ;
        RECT -8.820 93.280 -8.530 93.560 ;
        RECT 1.100 93.280 1.390 93.560 ;
        RECT 11.020 93.280 11.310 93.560 ;
        RECT 20.940 93.280 21.230 93.560 ;
        RECT -281.540 90.420 -281.250 90.700 ;
        RECT -271.620 90.420 -271.330 90.700 ;
        RECT -261.700 90.420 -261.410 90.700 ;
        RECT -251.780 90.420 -251.490 90.700 ;
        RECT -241.860 90.420 -241.570 90.700 ;
        RECT -231.940 90.420 -231.650 90.700 ;
        RECT -222.020 90.420 -221.730 90.700 ;
        RECT -212.100 90.420 -211.810 90.700 ;
        RECT -202.180 90.420 -201.890 90.700 ;
        RECT -192.260 90.420 -191.970 90.700 ;
        RECT -182.340 90.420 -182.050 90.700 ;
        RECT -172.420 90.420 -172.130 90.700 ;
        RECT -162.500 90.420 -162.210 90.700 ;
        RECT -152.580 90.420 -152.290 90.700 ;
        RECT -142.660 90.420 -142.370 90.700 ;
        RECT -132.740 90.420 -132.450 90.700 ;
        RECT -122.820 90.420 -122.530 90.700 ;
        RECT -112.900 90.420 -112.610 90.700 ;
        RECT -102.980 90.420 -102.690 90.700 ;
        RECT -93.060 90.420 -92.770 90.700 ;
        RECT -83.140 90.420 -82.850 90.700 ;
        RECT -73.220 90.420 -72.930 90.700 ;
        RECT -63.300 90.420 -63.010 90.700 ;
        RECT -53.380 90.420 -53.090 90.700 ;
        RECT -43.460 90.420 -43.170 90.700 ;
        RECT -33.540 90.420 -33.250 90.700 ;
        RECT -23.620 90.420 -23.330 90.700 ;
        RECT -13.700 90.420 -13.410 90.700 ;
        RECT -3.780 90.420 -3.490 90.700 ;
        RECT 6.140 90.420 6.430 90.700 ;
        RECT 16.060 90.420 16.350 90.700 ;
        RECT 25.980 90.420 26.270 90.700 ;
        RECT -286.880 88.880 -286.590 89.160 ;
        RECT -285.950 88.880 -285.660 89.160 ;
        RECT -276.960 88.880 -276.670 89.160 ;
        RECT -276.030 88.880 -275.740 89.160 ;
        RECT -267.040 88.880 -266.750 89.160 ;
        RECT -266.110 88.880 -265.820 89.160 ;
        RECT -257.120 88.880 -256.830 89.160 ;
        RECT -256.190 88.880 -255.900 89.160 ;
        RECT -247.200 88.880 -246.910 89.160 ;
        RECT -246.270 88.880 -245.980 89.160 ;
        RECT -237.280 88.880 -236.990 89.160 ;
        RECT -236.350 88.880 -236.060 89.160 ;
        RECT -227.360 88.880 -227.070 89.160 ;
        RECT -226.430 88.880 -226.140 89.160 ;
        RECT -217.440 88.880 -217.150 89.160 ;
        RECT -216.510 88.880 -216.220 89.160 ;
        RECT -207.520 88.880 -207.230 89.160 ;
        RECT -206.590 88.880 -206.300 89.160 ;
        RECT -197.600 88.880 -197.310 89.160 ;
        RECT -196.670 88.880 -196.380 89.160 ;
        RECT -187.680 88.880 -187.390 89.160 ;
        RECT -186.750 88.880 -186.460 89.160 ;
        RECT -177.760 88.880 -177.470 89.160 ;
        RECT -176.830 88.880 -176.540 89.160 ;
        RECT -167.840 88.880 -167.550 89.160 ;
        RECT -166.910 88.880 -166.620 89.160 ;
        RECT -157.920 88.880 -157.630 89.160 ;
        RECT -156.990 88.880 -156.700 89.160 ;
        RECT -148.000 88.880 -147.710 89.160 ;
        RECT -147.070 88.880 -146.780 89.160 ;
        RECT -138.080 88.880 -137.790 89.160 ;
        RECT -137.150 88.880 -136.860 89.160 ;
        RECT -128.160 88.880 -127.870 89.160 ;
        RECT -127.230 88.880 -126.940 89.160 ;
        RECT -118.240 88.880 -117.950 89.160 ;
        RECT -117.310 88.880 -117.020 89.160 ;
        RECT -108.320 88.880 -108.030 89.160 ;
        RECT -107.390 88.880 -107.100 89.160 ;
        RECT -98.400 88.880 -98.110 89.160 ;
        RECT -97.470 88.880 -97.180 89.160 ;
        RECT -88.480 88.880 -88.190 89.160 ;
        RECT -87.550 88.880 -87.260 89.160 ;
        RECT -78.560 88.880 -78.270 89.160 ;
        RECT -77.630 88.880 -77.340 89.160 ;
        RECT -68.640 88.880 -68.350 89.160 ;
        RECT -67.710 88.880 -67.420 89.160 ;
        RECT -58.720 88.880 -58.430 89.160 ;
        RECT -57.790 88.880 -57.500 89.160 ;
        RECT -48.800 88.880 -48.510 89.160 ;
        RECT -47.870 88.880 -47.580 89.160 ;
        RECT -38.880 88.880 -38.590 89.160 ;
        RECT -37.950 88.880 -37.660 89.160 ;
        RECT -28.960 88.880 -28.670 89.160 ;
        RECT -28.030 88.880 -27.740 89.160 ;
        RECT -19.040 88.880 -18.750 89.160 ;
        RECT -18.110 88.880 -17.820 89.160 ;
        RECT -9.120 88.880 -8.830 89.160 ;
        RECT -8.190 88.880 -7.900 89.160 ;
        RECT 0.800 88.880 1.090 89.160 ;
        RECT 1.730 88.880 2.020 89.160 ;
        RECT 10.720 88.880 11.010 89.160 ;
        RECT 11.650 88.880 11.940 89.160 ;
        RECT 20.640 88.880 20.930 89.160 ;
        RECT 21.570 88.880 21.860 89.160 ;
      LAYER met3 ;
        RECT -298.750 109.690 -293.660 109.870 ;
        RECT 29.330 109.690 34.420 109.750 ;
        RECT -298.750 100.060 34.420 109.690 ;
        RECT -298.750 82.780 -293.660 100.060 ;
        RECT -291.620 82.780 -290.850 100.060 ;
        RECT -286.660 89.210 -285.890 100.060 ;
        RECT -281.700 95.140 -280.930 100.060 ;
        RECT -282.020 94.730 -280.600 95.140 ;
        RECT -281.700 90.850 -280.930 94.730 ;
        RECT -281.910 90.370 -280.710 90.850 ;
        RECT -286.980 88.800 -285.560 89.210 ;
        RECT -286.660 82.780 -285.890 88.800 ;
        RECT -281.700 82.780 -280.930 90.370 ;
        RECT -276.760 89.210 -275.990 100.060 ;
        RECT -271.780 95.230 -271.010 100.060 ;
        RECT -271.780 95.140 -271.000 95.230 ;
        RECT -272.100 94.730 -270.680 95.140 ;
        RECT -271.780 92.780 -271.000 94.730 ;
        RECT -271.820 90.850 -271.000 92.780 ;
        RECT -271.990 90.370 -270.790 90.850 ;
        RECT -277.060 88.800 -275.640 89.210 ;
        RECT -271.820 88.880 -271.000 90.370 ;
        RECT -266.810 89.210 -266.040 100.060 ;
        RECT -261.820 95.140 -261.050 100.060 ;
        RECT -262.180 94.730 -260.760 95.140 ;
        RECT -261.820 90.850 -261.050 94.730 ;
        RECT -262.070 90.370 -260.870 90.850 ;
        RECT -276.760 82.780 -275.990 88.800 ;
        RECT -271.830 85.270 -271.000 88.880 ;
        RECT -267.140 88.800 -265.720 89.210 ;
        RECT -271.830 82.780 -271.010 85.270 ;
        RECT -266.810 82.780 -266.040 88.800 ;
        RECT -261.820 82.780 -261.050 90.370 ;
        RECT -256.920 89.210 -256.150 100.060 ;
        RECT -251.930 95.140 -251.160 100.060 ;
        RECT -252.260 94.730 -250.840 95.140 ;
        RECT -251.930 90.850 -251.160 94.730 ;
        RECT -252.150 90.370 -250.950 90.850 ;
        RECT -257.220 88.800 -255.800 89.210 ;
        RECT -256.920 82.780 -256.150 88.800 ;
        RECT -251.930 82.780 -251.160 90.370 ;
        RECT -246.990 89.210 -246.220 100.060 ;
        RECT -242.020 95.140 -241.250 100.060 ;
        RECT -242.340 94.730 -240.920 95.140 ;
        RECT -242.020 90.850 -241.250 94.730 ;
        RECT -242.230 90.370 -241.030 90.850 ;
        RECT -247.300 88.800 -245.880 89.210 ;
        RECT -246.990 82.780 -246.220 88.800 ;
        RECT -242.020 82.780 -241.250 90.370 ;
        RECT -237.080 89.210 -236.310 100.060 ;
        RECT -232.120 95.140 -231.350 100.060 ;
        RECT -232.420 94.730 -231.000 95.140 ;
        RECT -232.120 90.850 -231.350 94.730 ;
        RECT -232.310 90.370 -231.110 90.850 ;
        RECT -237.380 88.800 -235.960 89.210 ;
        RECT -237.080 82.780 -236.310 88.800 ;
        RECT -232.120 82.780 -231.350 90.370 ;
        RECT -227.150 89.210 -226.380 100.060 ;
        RECT -222.180 95.140 -221.410 100.060 ;
        RECT -222.500 94.730 -221.080 95.140 ;
        RECT -222.180 90.850 -221.410 94.730 ;
        RECT -222.390 90.370 -221.190 90.850 ;
        RECT -227.460 88.800 -226.040 89.210 ;
        RECT -227.150 82.780 -226.380 88.800 ;
        RECT -222.180 82.780 -221.410 90.370 ;
        RECT -217.200 89.210 -216.430 100.060 ;
        RECT -212.240 95.140 -211.470 100.060 ;
        RECT -212.580 94.730 -211.160 95.140 ;
        RECT -212.240 90.850 -211.470 94.730 ;
        RECT -212.470 90.370 -211.270 90.850 ;
        RECT -217.540 88.800 -216.120 89.210 ;
        RECT -217.200 82.780 -216.430 88.800 ;
        RECT -212.240 82.780 -211.470 90.370 ;
        RECT -207.290 89.210 -206.520 100.060 ;
        RECT -202.350 95.140 -201.580 100.060 ;
        RECT -202.660 94.730 -201.240 95.140 ;
        RECT -202.350 90.850 -201.580 94.730 ;
        RECT -202.550 90.370 -201.350 90.850 ;
        RECT -207.620 88.800 -206.200 89.210 ;
        RECT -207.290 82.780 -206.520 88.800 ;
        RECT -202.350 82.780 -201.580 90.370 ;
        RECT -197.420 89.210 -196.650 100.060 ;
        RECT -192.420 95.140 -191.650 100.060 ;
        RECT -192.740 94.730 -191.320 95.140 ;
        RECT -192.420 90.850 -191.650 94.730 ;
        RECT -192.630 90.370 -191.430 90.850 ;
        RECT -197.700 88.800 -196.280 89.210 ;
        RECT -197.420 82.780 -196.650 88.800 ;
        RECT -192.420 82.780 -191.650 90.370 ;
        RECT -187.460 89.210 -186.690 100.060 ;
        RECT -182.510 95.140 -181.740 100.060 ;
        RECT -182.820 94.730 -181.400 95.140 ;
        RECT -182.510 90.850 -181.740 94.730 ;
        RECT -182.710 90.370 -181.510 90.850 ;
        RECT -187.780 88.800 -186.360 89.210 ;
        RECT -187.460 82.780 -186.690 88.800 ;
        RECT -182.510 82.780 -181.740 90.370 ;
        RECT -177.550 89.210 -176.780 100.060 ;
        RECT -172.560 95.140 -171.790 100.060 ;
        RECT -172.900 94.730 -171.480 95.140 ;
        RECT -172.560 90.850 -171.790 94.730 ;
        RECT -172.790 90.370 -171.590 90.850 ;
        RECT -177.860 88.800 -176.440 89.210 ;
        RECT -177.550 82.780 -176.780 88.800 ;
        RECT -172.560 82.780 -171.790 90.370 ;
        RECT -167.620 89.210 -166.850 100.060 ;
        RECT -162.620 95.140 -161.850 100.060 ;
        RECT -162.980 94.730 -161.560 95.140 ;
        RECT -162.620 90.850 -161.850 94.730 ;
        RECT -162.870 90.370 -161.670 90.850 ;
        RECT -167.940 88.800 -166.520 89.210 ;
        RECT -167.620 82.780 -166.850 88.800 ;
        RECT -162.620 82.780 -161.850 90.370 ;
        RECT -157.710 89.210 -156.940 100.060 ;
        RECT -152.760 95.140 -151.990 100.060 ;
        RECT -153.060 94.730 -151.640 95.140 ;
        RECT -152.760 90.850 -151.990 94.730 ;
        RECT -152.950 90.370 -151.750 90.850 ;
        RECT -158.020 88.800 -156.600 89.210 ;
        RECT -157.710 82.780 -156.940 88.800 ;
        RECT -152.760 82.780 -151.990 90.370 ;
        RECT -147.790 89.210 -147.020 100.060 ;
        RECT -142.830 95.140 -142.060 100.060 ;
        RECT -143.140 94.730 -141.720 95.140 ;
        RECT -142.830 90.850 -142.060 94.730 ;
        RECT -143.030 90.370 -141.830 90.850 ;
        RECT -148.100 88.800 -146.680 89.210 ;
        RECT -147.790 82.780 -147.020 88.800 ;
        RECT -142.830 82.780 -142.060 90.370 ;
        RECT -137.850 89.210 -137.080 100.060 ;
        RECT -132.920 95.140 -132.150 100.060 ;
        RECT -133.220 94.730 -131.800 95.140 ;
        RECT -132.920 90.850 -132.150 94.730 ;
        RECT -133.110 90.370 -131.910 90.850 ;
        RECT -138.180 88.800 -136.760 89.210 ;
        RECT -137.850 82.780 -137.080 88.800 ;
        RECT -132.920 82.780 -132.150 90.370 ;
        RECT -127.940 89.210 -127.170 100.060 ;
        RECT -122.960 95.140 -122.190 100.060 ;
        RECT -123.300 94.730 -121.880 95.140 ;
        RECT -122.960 90.850 -122.190 94.730 ;
        RECT -123.190 90.370 -121.990 90.850 ;
        RECT -128.260 88.800 -126.840 89.210 ;
        RECT -127.940 82.780 -127.170 88.800 ;
        RECT -122.960 82.780 -122.190 90.370 ;
        RECT -118.040 89.210 -117.270 100.060 ;
        RECT -113.080 95.140 -112.310 100.060 ;
        RECT -113.380 94.730 -111.960 95.140 ;
        RECT -113.080 90.850 -112.310 94.730 ;
        RECT -113.270 90.370 -112.070 90.850 ;
        RECT -118.340 88.800 -116.920 89.210 ;
        RECT -118.040 82.780 -117.270 88.800 ;
        RECT -113.080 82.780 -112.310 90.370 ;
        RECT -108.110 89.210 -107.340 100.060 ;
        RECT -103.150 95.140 -102.380 100.060 ;
        RECT -103.460 94.730 -102.040 95.140 ;
        RECT -103.150 90.850 -102.380 94.730 ;
        RECT -103.350 90.370 -102.150 90.850 ;
        RECT -108.420 88.800 -107.000 89.210 ;
        RECT -108.110 82.780 -107.340 88.800 ;
        RECT -103.150 82.780 -102.380 90.370 ;
        RECT -98.160 89.210 -97.390 100.060 ;
        RECT -93.210 95.140 -92.440 100.060 ;
        RECT -93.540 94.730 -92.120 95.140 ;
        RECT -93.210 90.850 -92.440 94.730 ;
        RECT -93.430 90.370 -92.230 90.850 ;
        RECT -98.500 88.800 -97.080 89.210 ;
        RECT -98.160 82.780 -97.390 88.800 ;
        RECT -93.210 82.780 -92.440 90.370 ;
        RECT -88.260 89.210 -87.490 100.060 ;
        RECT -83.270 95.140 -82.500 100.060 ;
        RECT -83.620 94.730 -82.200 95.140 ;
        RECT -83.270 90.850 -82.500 94.730 ;
        RECT -83.510 90.370 -82.310 90.850 ;
        RECT -88.580 88.800 -87.160 89.210 ;
        RECT -88.260 82.780 -87.490 88.800 ;
        RECT -83.270 82.780 -82.500 90.370 ;
        RECT -78.350 89.210 -77.580 100.060 ;
        RECT -73.390 95.140 -72.620 100.060 ;
        RECT -73.700 94.730 -72.280 95.140 ;
        RECT -73.390 90.850 -72.620 94.730 ;
        RECT -73.590 90.370 -72.390 90.850 ;
        RECT -78.660 88.800 -77.240 89.210 ;
        RECT -78.350 82.780 -77.580 88.800 ;
        RECT -73.390 82.780 -72.620 90.370 ;
        RECT -68.410 89.210 -67.640 100.060 ;
        RECT -63.430 95.140 -62.660 100.060 ;
        RECT -63.780 94.730 -62.360 95.140 ;
        RECT -63.430 90.850 -62.660 94.730 ;
        RECT -63.670 90.370 -62.470 90.850 ;
        RECT -68.740 88.800 -67.320 89.210 ;
        RECT -68.410 82.780 -67.640 88.800 ;
        RECT -63.430 82.780 -62.660 90.370 ;
        RECT -58.520 89.210 -57.750 100.060 ;
        RECT -53.520 95.140 -52.750 100.060 ;
        RECT -53.860 94.730 -52.440 95.140 ;
        RECT -53.520 90.850 -52.750 94.730 ;
        RECT -53.750 90.370 -52.550 90.850 ;
        RECT -58.820 88.800 -57.400 89.210 ;
        RECT -58.520 82.780 -57.750 88.800 ;
        RECT -53.520 82.780 -52.750 90.370 ;
        RECT -48.560 89.210 -47.790 100.060 ;
        RECT -43.630 95.140 -42.860 100.060 ;
        RECT -43.940 94.730 -42.520 95.140 ;
        RECT -43.630 90.850 -42.860 94.730 ;
        RECT -43.830 90.370 -42.630 90.850 ;
        RECT -48.900 88.800 -47.480 89.210 ;
        RECT -48.560 82.780 -47.790 88.800 ;
        RECT -43.630 82.780 -42.860 90.370 ;
        RECT -38.680 89.210 -37.910 100.060 ;
        RECT -33.700 95.140 -32.930 100.060 ;
        RECT -34.020 94.730 -32.600 95.140 ;
        RECT -33.700 90.850 -32.930 94.730 ;
        RECT -33.910 90.370 -32.710 90.850 ;
        RECT -38.980 88.800 -37.560 89.210 ;
        RECT -38.680 82.780 -37.910 88.800 ;
        RECT -33.700 82.780 -32.930 90.370 ;
        RECT -28.750 89.210 -27.980 100.060 ;
        RECT -23.800 95.140 -23.030 100.060 ;
        RECT -24.100 94.730 -22.680 95.140 ;
        RECT -23.800 90.850 -23.030 94.730 ;
        RECT -23.990 90.370 -22.790 90.850 ;
        RECT -29.060 88.800 -27.640 89.210 ;
        RECT -28.750 82.780 -27.980 88.800 ;
        RECT -23.800 82.780 -23.030 90.370 ;
        RECT -18.820 89.210 -18.050 100.060 ;
        RECT -13.870 95.140 -13.100 100.060 ;
        RECT -14.180 94.730 -12.760 95.140 ;
        RECT -13.870 90.850 -13.100 94.730 ;
        RECT -14.070 90.370 -12.870 90.850 ;
        RECT -19.140 88.800 -17.720 89.210 ;
        RECT -18.820 82.780 -18.050 88.800 ;
        RECT -13.870 82.780 -13.100 90.370 ;
        RECT -8.920 89.210 -8.150 100.060 ;
        RECT -3.940 95.140 -3.170 100.060 ;
        RECT -4.260 94.730 -2.840 95.140 ;
        RECT -3.940 90.850 -3.170 94.730 ;
        RECT -4.150 90.370 -2.950 90.850 ;
        RECT -9.220 88.800 -7.800 89.210 ;
        RECT -8.920 82.780 -8.150 88.800 ;
        RECT -3.940 82.780 -3.170 90.370 ;
        RECT 1.010 89.210 1.780 100.060 ;
        RECT 5.940 95.140 6.710 100.060 ;
        RECT 5.660 94.730 7.080 95.140 ;
        RECT 5.940 90.850 6.710 94.730 ;
        RECT 5.770 90.370 6.970 90.850 ;
        RECT 0.700 88.800 2.120 89.210 ;
        RECT 1.010 82.780 1.780 88.800 ;
        RECT 5.940 82.780 6.710 90.370 ;
        RECT 10.940 89.210 11.710 100.060 ;
        RECT 15.890 95.140 16.660 100.060 ;
        RECT 15.580 94.730 17.000 95.140 ;
        RECT 15.890 90.850 16.660 94.730 ;
        RECT 15.690 90.370 16.890 90.850 ;
        RECT 10.620 88.800 12.040 89.210 ;
        RECT 10.940 82.780 11.710 88.800 ;
        RECT 15.890 82.780 16.660 90.370 ;
        RECT 20.870 89.210 21.640 100.060 ;
        RECT 25.880 95.140 26.650 100.060 ;
        RECT 25.500 94.730 26.650 95.140 ;
        RECT 25.880 90.850 26.650 94.730 ;
        RECT 25.610 90.370 26.440 90.850 ;
        RECT 20.540 88.800 21.960 89.210 ;
        RECT 20.870 82.780 21.640 88.800 ;
        RECT 25.880 82.780 26.650 90.370 ;
        RECT 29.330 83.200 34.420 100.060 ;
        RECT 27.700 82.780 164.350 83.200 ;
        RECT -298.750 73.570 164.350 82.780 ;
        RECT -298.750 73.150 34.420 73.570 ;
        RECT -298.750 73.140 -293.660 73.150 ;
        RECT 29.330 73.020 34.420 73.150 ;
    END
  END VPWR
  OBS
      LAYER pwell ;
        RECT -280.030 159.090 142.600 365.400 ;
      LAYER nwell ;
        RECT -290.950 95.095 -289.345 95.330 ;
        RECT -291.650 93.570 -289.345 95.095 ;
        RECT -291.650 93.510 -290.810 93.570 ;
      LAYER pwell ;
        RECT -290.860 93.225 -290.690 93.415 ;
        RECT 25.670 93.225 25.840 93.415 ;
        RECT -290.975 93.220 -289.625 93.225 ;
        RECT -291.440 93.140 -289.625 93.220 ;
        RECT -291.445 92.355 -289.625 93.140 ;
        RECT -291.440 92.350 -289.625 92.355 ;
        RECT -290.975 92.315 -289.625 92.350 ;
        RECT 24.605 93.220 25.955 93.225 ;
        RECT 24.605 93.140 26.420 93.220 ;
        RECT 24.605 92.355 26.425 93.140 ;
        RECT 24.605 92.320 26.420 92.355 ;
        RECT 24.605 92.315 25.955 92.320 ;
      LAYER nwell ;
        RECT -291.650 90.420 -289.430 92.025 ;
      LAYER pwell ;
        RECT -289.355 90.025 -288.575 90.175 ;
        RECT -289.545 90.020 -288.575 90.025 ;
        RECT -290.140 90.015 -288.575 90.020 ;
        RECT -290.145 89.230 -288.575 90.015 ;
        RECT -289.355 88.805 -288.575 89.230 ;
        RECT 23.555 90.025 24.335 90.175 ;
        RECT 23.555 90.020 24.525 90.025 ;
        RECT 23.555 88.810 25.130 90.020 ;
        RECT 23.555 88.805 24.335 88.810 ;
      LAYER nwell ;
        RECT -291.450 -182.150 131.180 24.160 ;
      LAYER li1 ;
        RECT -290.845 94.990 -290.675 95.140 ;
        RECT -291.460 94.820 -290.675 94.990 ;
        RECT -291.375 93.655 -291.085 94.820 ;
        RECT -290.845 94.615 -290.675 94.820 ;
        RECT -290.505 94.875 -288.295 95.055 ;
        RECT -290.505 94.785 -289.600 94.875 ;
        RECT -288.800 94.795 -288.295 94.875 ;
        RECT -280.585 94.875 -278.375 95.055 ;
        RECT -280.585 94.785 -279.680 94.875 ;
        RECT -278.880 94.795 -278.375 94.875 ;
        RECT -270.665 94.875 -268.455 95.055 ;
        RECT -270.665 94.785 -269.760 94.875 ;
        RECT -268.960 94.795 -268.455 94.875 ;
        RECT -260.745 94.875 -258.535 95.055 ;
        RECT -260.745 94.785 -259.840 94.875 ;
        RECT -259.040 94.795 -258.535 94.875 ;
        RECT -250.825 94.875 -248.615 95.055 ;
        RECT -250.825 94.785 -249.920 94.875 ;
        RECT -249.120 94.795 -248.615 94.875 ;
        RECT -240.905 94.875 -238.695 95.055 ;
        RECT -240.905 94.785 -240.000 94.875 ;
        RECT -239.200 94.795 -238.695 94.875 ;
        RECT -230.985 94.875 -228.775 95.055 ;
        RECT -230.985 94.785 -230.080 94.875 ;
        RECT -229.280 94.795 -228.775 94.875 ;
        RECT -221.065 94.875 -218.855 95.055 ;
        RECT -221.065 94.785 -220.160 94.875 ;
        RECT -219.360 94.795 -218.855 94.875 ;
        RECT -211.145 94.875 -208.935 95.055 ;
        RECT -211.145 94.785 -210.240 94.875 ;
        RECT -209.440 94.795 -208.935 94.875 ;
        RECT -201.225 94.875 -199.015 95.055 ;
        RECT -201.225 94.785 -200.320 94.875 ;
        RECT -199.520 94.795 -199.015 94.875 ;
        RECT -191.305 94.875 -189.095 95.055 ;
        RECT -191.305 94.785 -190.400 94.875 ;
        RECT -189.600 94.795 -189.095 94.875 ;
        RECT -181.385 94.875 -179.175 95.055 ;
        RECT -181.385 94.785 -180.480 94.875 ;
        RECT -179.680 94.795 -179.175 94.875 ;
        RECT -171.465 94.875 -169.255 95.055 ;
        RECT -171.465 94.785 -170.560 94.875 ;
        RECT -169.760 94.795 -169.255 94.875 ;
        RECT -161.545 94.875 -159.335 95.055 ;
        RECT -161.545 94.785 -160.640 94.875 ;
        RECT -159.840 94.795 -159.335 94.875 ;
        RECT -151.625 94.875 -149.415 95.055 ;
        RECT -151.625 94.785 -150.720 94.875 ;
        RECT -149.920 94.795 -149.415 94.875 ;
        RECT -141.705 94.875 -139.495 95.055 ;
        RECT -141.705 94.785 -140.800 94.875 ;
        RECT -140.000 94.795 -139.495 94.875 ;
        RECT -131.785 94.875 -129.575 95.055 ;
        RECT -131.785 94.785 -130.880 94.875 ;
        RECT -130.080 94.795 -129.575 94.875 ;
        RECT -121.865 94.875 -119.655 95.055 ;
        RECT -121.865 94.785 -120.960 94.875 ;
        RECT -120.160 94.795 -119.655 94.875 ;
        RECT -111.945 94.875 -109.735 95.055 ;
        RECT -111.945 94.785 -111.040 94.875 ;
        RECT -110.240 94.795 -109.735 94.875 ;
        RECT -102.025 94.875 -99.815 95.055 ;
        RECT -102.025 94.785 -101.120 94.875 ;
        RECT -100.320 94.795 -99.815 94.875 ;
        RECT -92.105 94.875 -89.895 95.055 ;
        RECT -92.105 94.785 -91.200 94.875 ;
        RECT -90.400 94.795 -89.895 94.875 ;
        RECT -82.185 94.875 -79.975 95.055 ;
        RECT -82.185 94.785 -81.280 94.875 ;
        RECT -80.480 94.795 -79.975 94.875 ;
        RECT -72.265 94.875 -70.055 95.055 ;
        RECT -72.265 94.785 -71.360 94.875 ;
        RECT -70.560 94.795 -70.055 94.875 ;
        RECT -62.345 94.875 -60.135 95.055 ;
        RECT -62.345 94.785 -61.440 94.875 ;
        RECT -60.640 94.795 -60.135 94.875 ;
        RECT -52.425 94.875 -50.215 95.055 ;
        RECT -52.425 94.785 -51.520 94.875 ;
        RECT -50.720 94.795 -50.215 94.875 ;
        RECT -42.505 94.875 -40.295 95.055 ;
        RECT -42.505 94.785 -41.600 94.875 ;
        RECT -40.800 94.795 -40.295 94.875 ;
        RECT -32.585 94.875 -30.375 95.055 ;
        RECT -32.585 94.785 -31.680 94.875 ;
        RECT -30.880 94.795 -30.375 94.875 ;
        RECT -22.665 94.875 -20.455 95.055 ;
        RECT -22.665 94.785 -21.760 94.875 ;
        RECT -20.960 94.795 -20.455 94.875 ;
        RECT -12.745 94.875 -10.535 95.055 ;
        RECT -12.745 94.785 -11.840 94.875 ;
        RECT -11.040 94.795 -10.535 94.875 ;
        RECT -2.825 94.875 -0.615 95.055 ;
        RECT -2.825 94.785 -1.920 94.875 ;
        RECT -1.120 94.795 -0.615 94.875 ;
        RECT 7.095 94.875 9.305 95.055 ;
        RECT 7.095 94.785 8.000 94.875 ;
        RECT 8.800 94.795 9.305 94.875 ;
        RECT 17.015 94.875 19.225 95.055 ;
        RECT 17.015 94.785 17.920 94.875 ;
        RECT 18.720 94.795 19.225 94.875 ;
        RECT -290.845 94.285 -289.915 94.615 ;
        RECT -289.430 94.600 -289.100 94.705 ;
        RECT -283.440 94.600 -283.110 94.705 ;
        RECT -279.510 94.600 -279.180 94.705 ;
        RECT -273.520 94.600 -273.190 94.705 ;
        RECT -269.590 94.600 -269.260 94.705 ;
        RECT -263.600 94.600 -263.270 94.705 ;
        RECT -259.670 94.600 -259.340 94.705 ;
        RECT -253.680 94.600 -253.350 94.705 ;
        RECT -249.750 94.600 -249.420 94.705 ;
        RECT -243.760 94.600 -243.430 94.705 ;
        RECT -239.830 94.600 -239.500 94.705 ;
        RECT -233.840 94.600 -233.510 94.705 ;
        RECT -229.910 94.600 -229.580 94.705 ;
        RECT -223.920 94.600 -223.590 94.705 ;
        RECT -219.990 94.600 -219.660 94.705 ;
        RECT -214.000 94.600 -213.670 94.705 ;
        RECT -210.070 94.600 -209.740 94.705 ;
        RECT -204.080 94.600 -203.750 94.705 ;
        RECT -200.150 94.600 -199.820 94.705 ;
        RECT -194.160 94.600 -193.830 94.705 ;
        RECT -190.230 94.600 -189.900 94.705 ;
        RECT -184.240 94.600 -183.910 94.705 ;
        RECT -180.310 94.600 -179.980 94.705 ;
        RECT -174.320 94.600 -173.990 94.705 ;
        RECT -170.390 94.600 -170.060 94.705 ;
        RECT -164.400 94.600 -164.070 94.705 ;
        RECT -160.470 94.600 -160.140 94.705 ;
        RECT -154.480 94.600 -154.150 94.705 ;
        RECT -150.550 94.600 -150.220 94.705 ;
        RECT -144.560 94.600 -144.230 94.705 ;
        RECT -140.630 94.600 -140.300 94.705 ;
        RECT -134.640 94.600 -134.310 94.705 ;
        RECT -130.710 94.600 -130.380 94.705 ;
        RECT -124.720 94.600 -124.390 94.705 ;
        RECT -120.790 94.600 -120.460 94.705 ;
        RECT -114.800 94.600 -114.470 94.705 ;
        RECT -110.870 94.600 -110.540 94.705 ;
        RECT -104.880 94.600 -104.550 94.705 ;
        RECT -100.950 94.600 -100.620 94.705 ;
        RECT -94.960 94.600 -94.630 94.705 ;
        RECT -91.030 94.600 -90.700 94.705 ;
        RECT -85.040 94.600 -84.710 94.705 ;
        RECT -81.110 94.600 -80.780 94.705 ;
        RECT -75.120 94.600 -74.790 94.705 ;
        RECT -71.190 94.600 -70.860 94.705 ;
        RECT -65.200 94.600 -64.870 94.705 ;
        RECT -61.270 94.600 -60.940 94.705 ;
        RECT -55.280 94.600 -54.950 94.705 ;
        RECT -51.350 94.600 -51.020 94.705 ;
        RECT -45.360 94.600 -45.030 94.705 ;
        RECT -41.430 94.600 -41.100 94.705 ;
        RECT -35.440 94.600 -35.110 94.705 ;
        RECT -31.510 94.600 -31.180 94.705 ;
        RECT -25.520 94.600 -25.190 94.705 ;
        RECT -21.590 94.600 -21.260 94.705 ;
        RECT -15.600 94.600 -15.270 94.705 ;
        RECT -11.670 94.600 -11.340 94.705 ;
        RECT -5.680 94.600 -5.350 94.705 ;
        RECT -1.750 94.600 -1.420 94.705 ;
        RECT 4.240 94.600 4.570 94.705 ;
        RECT 8.170 94.600 8.500 94.705 ;
        RECT 14.160 94.600 14.490 94.705 ;
        RECT 18.090 94.600 18.420 94.705 ;
        RECT 24.080 94.600 24.410 94.705 ;
        RECT -289.745 94.430 -288.675 94.600 ;
        RECT -290.845 93.760 -290.675 94.285 ;
        RECT -289.745 94.105 -289.575 94.430 ;
        RECT -290.505 93.925 -289.575 94.105 ;
        RECT -289.395 93.865 -289.025 94.205 ;
        RECT -288.845 94.105 -288.675 94.430 ;
        RECT -283.865 94.430 -282.795 94.600 ;
        RECT -283.865 94.105 -283.695 94.430 ;
        RECT -288.845 93.935 -288.295 94.105 ;
        RECT -284.245 93.935 -283.695 94.105 ;
        RECT -283.515 93.865 -283.145 94.205 ;
        RECT -282.965 94.105 -282.795 94.430 ;
        RECT -279.825 94.430 -278.755 94.600 ;
        RECT -279.825 94.105 -279.655 94.430 ;
        RECT -282.965 93.925 -282.035 94.105 ;
        RECT -280.585 93.925 -279.655 94.105 ;
        RECT -279.475 93.865 -279.105 94.205 ;
        RECT -278.925 94.105 -278.755 94.430 ;
        RECT -273.945 94.430 -272.875 94.600 ;
        RECT -273.945 94.105 -273.775 94.430 ;
        RECT -278.925 93.935 -278.375 94.105 ;
        RECT -274.325 93.935 -273.775 94.105 ;
        RECT -273.595 93.865 -273.225 94.205 ;
        RECT -273.045 94.105 -272.875 94.430 ;
        RECT -269.905 94.430 -268.835 94.600 ;
        RECT -269.905 94.105 -269.735 94.430 ;
        RECT -273.045 93.925 -272.115 94.105 ;
        RECT -270.665 93.925 -269.735 94.105 ;
        RECT -269.555 93.865 -269.185 94.205 ;
        RECT -269.005 94.105 -268.835 94.430 ;
        RECT -264.025 94.430 -262.955 94.600 ;
        RECT -264.025 94.105 -263.855 94.430 ;
        RECT -269.005 93.935 -268.455 94.105 ;
        RECT -264.405 93.935 -263.855 94.105 ;
        RECT -263.675 93.865 -263.305 94.205 ;
        RECT -263.125 94.105 -262.955 94.430 ;
        RECT -259.985 94.430 -258.915 94.600 ;
        RECT -259.985 94.105 -259.815 94.430 ;
        RECT -263.125 93.925 -262.195 94.105 ;
        RECT -260.745 93.925 -259.815 94.105 ;
        RECT -259.635 93.865 -259.265 94.205 ;
        RECT -259.085 94.105 -258.915 94.430 ;
        RECT -254.105 94.430 -253.035 94.600 ;
        RECT -254.105 94.105 -253.935 94.430 ;
        RECT -259.085 93.935 -258.535 94.105 ;
        RECT -254.485 93.935 -253.935 94.105 ;
        RECT -253.755 93.865 -253.385 94.205 ;
        RECT -253.205 94.105 -253.035 94.430 ;
        RECT -250.065 94.430 -248.995 94.600 ;
        RECT -250.065 94.105 -249.895 94.430 ;
        RECT -253.205 93.925 -252.275 94.105 ;
        RECT -250.825 93.925 -249.895 94.105 ;
        RECT -249.715 93.865 -249.345 94.205 ;
        RECT -249.165 94.105 -248.995 94.430 ;
        RECT -244.185 94.430 -243.115 94.600 ;
        RECT -244.185 94.105 -244.015 94.430 ;
        RECT -249.165 93.935 -248.615 94.105 ;
        RECT -244.565 93.935 -244.015 94.105 ;
        RECT -243.835 93.865 -243.465 94.205 ;
        RECT -243.285 94.105 -243.115 94.430 ;
        RECT -240.145 94.430 -239.075 94.600 ;
        RECT -240.145 94.105 -239.975 94.430 ;
        RECT -243.285 93.925 -242.355 94.105 ;
        RECT -240.905 93.925 -239.975 94.105 ;
        RECT -239.795 93.865 -239.425 94.205 ;
        RECT -239.245 94.105 -239.075 94.430 ;
        RECT -234.265 94.430 -233.195 94.600 ;
        RECT -234.265 94.105 -234.095 94.430 ;
        RECT -239.245 93.935 -238.695 94.105 ;
        RECT -234.645 93.935 -234.095 94.105 ;
        RECT -233.915 93.865 -233.545 94.205 ;
        RECT -233.365 94.105 -233.195 94.430 ;
        RECT -230.225 94.430 -229.155 94.600 ;
        RECT -230.225 94.105 -230.055 94.430 ;
        RECT -233.365 93.925 -232.435 94.105 ;
        RECT -230.985 93.925 -230.055 94.105 ;
        RECT -229.875 93.865 -229.505 94.205 ;
        RECT -229.325 94.105 -229.155 94.430 ;
        RECT -224.345 94.430 -223.275 94.600 ;
        RECT -224.345 94.105 -224.175 94.430 ;
        RECT -229.325 93.935 -228.775 94.105 ;
        RECT -224.725 93.935 -224.175 94.105 ;
        RECT -223.995 93.865 -223.625 94.205 ;
        RECT -223.445 94.105 -223.275 94.430 ;
        RECT -220.305 94.430 -219.235 94.600 ;
        RECT -220.305 94.105 -220.135 94.430 ;
        RECT -223.445 93.925 -222.515 94.105 ;
        RECT -221.065 93.925 -220.135 94.105 ;
        RECT -219.955 93.865 -219.585 94.205 ;
        RECT -219.405 94.105 -219.235 94.430 ;
        RECT -214.425 94.430 -213.355 94.600 ;
        RECT -214.425 94.105 -214.255 94.430 ;
        RECT -219.405 93.935 -218.855 94.105 ;
        RECT -214.805 93.935 -214.255 94.105 ;
        RECT -214.075 93.865 -213.705 94.205 ;
        RECT -213.525 94.105 -213.355 94.430 ;
        RECT -210.385 94.430 -209.315 94.600 ;
        RECT -210.385 94.105 -210.215 94.430 ;
        RECT -213.525 93.925 -212.595 94.105 ;
        RECT -211.145 93.925 -210.215 94.105 ;
        RECT -210.035 93.865 -209.665 94.205 ;
        RECT -209.485 94.105 -209.315 94.430 ;
        RECT -204.505 94.430 -203.435 94.600 ;
        RECT -204.505 94.105 -204.335 94.430 ;
        RECT -209.485 93.935 -208.935 94.105 ;
        RECT -204.885 93.935 -204.335 94.105 ;
        RECT -204.155 93.865 -203.785 94.205 ;
        RECT -203.605 94.105 -203.435 94.430 ;
        RECT -200.465 94.430 -199.395 94.600 ;
        RECT -200.465 94.105 -200.295 94.430 ;
        RECT -203.605 93.925 -202.675 94.105 ;
        RECT -201.225 93.925 -200.295 94.105 ;
        RECT -200.115 93.865 -199.745 94.205 ;
        RECT -199.565 94.105 -199.395 94.430 ;
        RECT -194.585 94.430 -193.515 94.600 ;
        RECT -194.585 94.105 -194.415 94.430 ;
        RECT -199.565 93.935 -199.015 94.105 ;
        RECT -194.965 93.935 -194.415 94.105 ;
        RECT -194.235 93.865 -193.865 94.205 ;
        RECT -193.685 94.105 -193.515 94.430 ;
        RECT -190.545 94.430 -189.475 94.600 ;
        RECT -190.545 94.105 -190.375 94.430 ;
        RECT -193.685 93.925 -192.755 94.105 ;
        RECT -191.305 93.925 -190.375 94.105 ;
        RECT -190.195 93.865 -189.825 94.205 ;
        RECT -189.645 94.105 -189.475 94.430 ;
        RECT -184.665 94.430 -183.595 94.600 ;
        RECT -184.665 94.105 -184.495 94.430 ;
        RECT -189.645 93.935 -189.095 94.105 ;
        RECT -185.045 93.935 -184.495 94.105 ;
        RECT -184.315 93.865 -183.945 94.205 ;
        RECT -183.765 94.105 -183.595 94.430 ;
        RECT -180.625 94.430 -179.555 94.600 ;
        RECT -180.625 94.105 -180.455 94.430 ;
        RECT -183.765 93.925 -182.835 94.105 ;
        RECT -181.385 93.925 -180.455 94.105 ;
        RECT -180.275 93.865 -179.905 94.205 ;
        RECT -179.725 94.105 -179.555 94.430 ;
        RECT -174.745 94.430 -173.675 94.600 ;
        RECT -174.745 94.105 -174.575 94.430 ;
        RECT -179.725 93.935 -179.175 94.105 ;
        RECT -175.125 93.935 -174.575 94.105 ;
        RECT -174.395 93.865 -174.025 94.205 ;
        RECT -173.845 94.105 -173.675 94.430 ;
        RECT -170.705 94.430 -169.635 94.600 ;
        RECT -170.705 94.105 -170.535 94.430 ;
        RECT -173.845 93.925 -172.915 94.105 ;
        RECT -171.465 93.925 -170.535 94.105 ;
        RECT -170.355 93.865 -169.985 94.205 ;
        RECT -169.805 94.105 -169.635 94.430 ;
        RECT -164.825 94.430 -163.755 94.600 ;
        RECT -164.825 94.105 -164.655 94.430 ;
        RECT -169.805 93.935 -169.255 94.105 ;
        RECT -165.205 93.935 -164.655 94.105 ;
        RECT -164.475 93.865 -164.105 94.205 ;
        RECT -163.925 94.105 -163.755 94.430 ;
        RECT -160.785 94.430 -159.715 94.600 ;
        RECT -160.785 94.105 -160.615 94.430 ;
        RECT -163.925 93.925 -162.995 94.105 ;
        RECT -161.545 93.925 -160.615 94.105 ;
        RECT -160.435 93.865 -160.065 94.205 ;
        RECT -159.885 94.105 -159.715 94.430 ;
        RECT -154.905 94.430 -153.835 94.600 ;
        RECT -154.905 94.105 -154.735 94.430 ;
        RECT -159.885 93.935 -159.335 94.105 ;
        RECT -155.285 93.935 -154.735 94.105 ;
        RECT -154.555 93.865 -154.185 94.205 ;
        RECT -154.005 94.105 -153.835 94.430 ;
        RECT -150.865 94.430 -149.795 94.600 ;
        RECT -150.865 94.105 -150.695 94.430 ;
        RECT -154.005 93.925 -153.075 94.105 ;
        RECT -151.625 93.925 -150.695 94.105 ;
        RECT -150.515 93.865 -150.145 94.205 ;
        RECT -149.965 94.105 -149.795 94.430 ;
        RECT -144.985 94.430 -143.915 94.600 ;
        RECT -144.985 94.105 -144.815 94.430 ;
        RECT -149.965 93.935 -149.415 94.105 ;
        RECT -145.365 93.935 -144.815 94.105 ;
        RECT -144.635 93.865 -144.265 94.205 ;
        RECT -144.085 94.105 -143.915 94.430 ;
        RECT -140.945 94.430 -139.875 94.600 ;
        RECT -140.945 94.105 -140.775 94.430 ;
        RECT -144.085 93.925 -143.155 94.105 ;
        RECT -141.705 93.925 -140.775 94.105 ;
        RECT -140.595 93.865 -140.225 94.205 ;
        RECT -140.045 94.105 -139.875 94.430 ;
        RECT -135.065 94.430 -133.995 94.600 ;
        RECT -135.065 94.105 -134.895 94.430 ;
        RECT -140.045 93.935 -139.495 94.105 ;
        RECT -135.445 93.935 -134.895 94.105 ;
        RECT -134.715 93.865 -134.345 94.205 ;
        RECT -134.165 94.105 -133.995 94.430 ;
        RECT -131.025 94.430 -129.955 94.600 ;
        RECT -131.025 94.105 -130.855 94.430 ;
        RECT -134.165 93.925 -133.235 94.105 ;
        RECT -131.785 93.925 -130.855 94.105 ;
        RECT -130.675 93.865 -130.305 94.205 ;
        RECT -130.125 94.105 -129.955 94.430 ;
        RECT -125.145 94.430 -124.075 94.600 ;
        RECT -125.145 94.105 -124.975 94.430 ;
        RECT -130.125 93.935 -129.575 94.105 ;
        RECT -125.525 93.935 -124.975 94.105 ;
        RECT -124.795 93.865 -124.425 94.205 ;
        RECT -124.245 94.105 -124.075 94.430 ;
        RECT -121.105 94.430 -120.035 94.600 ;
        RECT -121.105 94.105 -120.935 94.430 ;
        RECT -124.245 93.925 -123.315 94.105 ;
        RECT -121.865 93.925 -120.935 94.105 ;
        RECT -120.755 93.865 -120.385 94.205 ;
        RECT -120.205 94.105 -120.035 94.430 ;
        RECT -115.225 94.430 -114.155 94.600 ;
        RECT -115.225 94.105 -115.055 94.430 ;
        RECT -120.205 93.935 -119.655 94.105 ;
        RECT -115.605 93.935 -115.055 94.105 ;
        RECT -114.875 93.865 -114.505 94.205 ;
        RECT -114.325 94.105 -114.155 94.430 ;
        RECT -111.185 94.430 -110.115 94.600 ;
        RECT -111.185 94.105 -111.015 94.430 ;
        RECT -114.325 93.925 -113.395 94.105 ;
        RECT -111.945 93.925 -111.015 94.105 ;
        RECT -110.835 93.865 -110.465 94.205 ;
        RECT -110.285 94.105 -110.115 94.430 ;
        RECT -105.305 94.430 -104.235 94.600 ;
        RECT -105.305 94.105 -105.135 94.430 ;
        RECT -110.285 93.935 -109.735 94.105 ;
        RECT -105.685 93.935 -105.135 94.105 ;
        RECT -104.955 93.865 -104.585 94.205 ;
        RECT -104.405 94.105 -104.235 94.430 ;
        RECT -101.265 94.430 -100.195 94.600 ;
        RECT -101.265 94.105 -101.095 94.430 ;
        RECT -104.405 93.925 -103.475 94.105 ;
        RECT -102.025 93.925 -101.095 94.105 ;
        RECT -100.915 93.865 -100.545 94.205 ;
        RECT -100.365 94.105 -100.195 94.430 ;
        RECT -95.385 94.430 -94.315 94.600 ;
        RECT -95.385 94.105 -95.215 94.430 ;
        RECT -100.365 93.935 -99.815 94.105 ;
        RECT -95.765 93.935 -95.215 94.105 ;
        RECT -95.035 93.865 -94.665 94.205 ;
        RECT -94.485 94.105 -94.315 94.430 ;
        RECT -91.345 94.430 -90.275 94.600 ;
        RECT -91.345 94.105 -91.175 94.430 ;
        RECT -94.485 93.925 -93.555 94.105 ;
        RECT -92.105 93.925 -91.175 94.105 ;
        RECT -90.995 93.865 -90.625 94.205 ;
        RECT -90.445 94.105 -90.275 94.430 ;
        RECT -85.465 94.430 -84.395 94.600 ;
        RECT -85.465 94.105 -85.295 94.430 ;
        RECT -90.445 93.935 -89.895 94.105 ;
        RECT -85.845 93.935 -85.295 94.105 ;
        RECT -85.115 93.865 -84.745 94.205 ;
        RECT -84.565 94.105 -84.395 94.430 ;
        RECT -81.425 94.430 -80.355 94.600 ;
        RECT -81.425 94.105 -81.255 94.430 ;
        RECT -84.565 93.925 -83.635 94.105 ;
        RECT -82.185 93.925 -81.255 94.105 ;
        RECT -81.075 93.865 -80.705 94.205 ;
        RECT -80.525 94.105 -80.355 94.430 ;
        RECT -75.545 94.430 -74.475 94.600 ;
        RECT -75.545 94.105 -75.375 94.430 ;
        RECT -80.525 93.935 -79.975 94.105 ;
        RECT -75.925 93.935 -75.375 94.105 ;
        RECT -75.195 93.865 -74.825 94.205 ;
        RECT -74.645 94.105 -74.475 94.430 ;
        RECT -71.505 94.430 -70.435 94.600 ;
        RECT -71.505 94.105 -71.335 94.430 ;
        RECT -74.645 93.925 -73.715 94.105 ;
        RECT -72.265 93.925 -71.335 94.105 ;
        RECT -71.155 93.865 -70.785 94.205 ;
        RECT -70.605 94.105 -70.435 94.430 ;
        RECT -65.625 94.430 -64.555 94.600 ;
        RECT -65.625 94.105 -65.455 94.430 ;
        RECT -70.605 93.935 -70.055 94.105 ;
        RECT -66.005 93.935 -65.455 94.105 ;
        RECT -65.275 93.865 -64.905 94.205 ;
        RECT -64.725 94.105 -64.555 94.430 ;
        RECT -61.585 94.430 -60.515 94.600 ;
        RECT -61.585 94.105 -61.415 94.430 ;
        RECT -64.725 93.925 -63.795 94.105 ;
        RECT -62.345 93.925 -61.415 94.105 ;
        RECT -61.235 93.865 -60.865 94.205 ;
        RECT -60.685 94.105 -60.515 94.430 ;
        RECT -55.705 94.430 -54.635 94.600 ;
        RECT -55.705 94.105 -55.535 94.430 ;
        RECT -60.685 93.935 -60.135 94.105 ;
        RECT -56.085 93.935 -55.535 94.105 ;
        RECT -55.355 93.865 -54.985 94.205 ;
        RECT -54.805 94.105 -54.635 94.430 ;
        RECT -51.665 94.430 -50.595 94.600 ;
        RECT -51.665 94.105 -51.495 94.430 ;
        RECT -54.805 93.925 -53.875 94.105 ;
        RECT -52.425 93.925 -51.495 94.105 ;
        RECT -51.315 93.865 -50.945 94.205 ;
        RECT -50.765 94.105 -50.595 94.430 ;
        RECT -45.785 94.430 -44.715 94.600 ;
        RECT -45.785 94.105 -45.615 94.430 ;
        RECT -50.765 93.935 -50.215 94.105 ;
        RECT -46.165 93.935 -45.615 94.105 ;
        RECT -45.435 93.865 -45.065 94.205 ;
        RECT -44.885 94.105 -44.715 94.430 ;
        RECT -41.745 94.430 -40.675 94.600 ;
        RECT -41.745 94.105 -41.575 94.430 ;
        RECT -44.885 93.925 -43.955 94.105 ;
        RECT -42.505 93.925 -41.575 94.105 ;
        RECT -41.395 93.865 -41.025 94.205 ;
        RECT -40.845 94.105 -40.675 94.430 ;
        RECT -35.865 94.430 -34.795 94.600 ;
        RECT -35.865 94.105 -35.695 94.430 ;
        RECT -40.845 93.935 -40.295 94.105 ;
        RECT -36.245 93.935 -35.695 94.105 ;
        RECT -35.515 93.865 -35.145 94.205 ;
        RECT -34.965 94.105 -34.795 94.430 ;
        RECT -31.825 94.430 -30.755 94.600 ;
        RECT -31.825 94.105 -31.655 94.430 ;
        RECT -34.965 93.925 -34.035 94.105 ;
        RECT -32.585 93.925 -31.655 94.105 ;
        RECT -31.475 93.865 -31.105 94.205 ;
        RECT -30.925 94.105 -30.755 94.430 ;
        RECT -25.945 94.430 -24.875 94.600 ;
        RECT -25.945 94.105 -25.775 94.430 ;
        RECT -30.925 93.935 -30.375 94.105 ;
        RECT -26.325 93.935 -25.775 94.105 ;
        RECT -25.595 93.865 -25.225 94.205 ;
        RECT -25.045 94.105 -24.875 94.430 ;
        RECT -21.905 94.430 -20.835 94.600 ;
        RECT -21.905 94.105 -21.735 94.430 ;
        RECT -25.045 93.925 -24.115 94.105 ;
        RECT -22.665 93.925 -21.735 94.105 ;
        RECT -21.555 93.865 -21.185 94.205 ;
        RECT -21.005 94.105 -20.835 94.430 ;
        RECT -16.025 94.430 -14.955 94.600 ;
        RECT -16.025 94.105 -15.855 94.430 ;
        RECT -21.005 93.935 -20.455 94.105 ;
        RECT -16.405 93.935 -15.855 94.105 ;
        RECT -15.675 93.865 -15.305 94.205 ;
        RECT -15.125 94.105 -14.955 94.430 ;
        RECT -11.985 94.430 -10.915 94.600 ;
        RECT -11.985 94.105 -11.815 94.430 ;
        RECT -15.125 93.925 -14.195 94.105 ;
        RECT -12.745 93.925 -11.815 94.105 ;
        RECT -11.635 93.865 -11.265 94.205 ;
        RECT -11.085 94.105 -10.915 94.430 ;
        RECT -6.105 94.430 -5.035 94.600 ;
        RECT -6.105 94.105 -5.935 94.430 ;
        RECT -11.085 93.935 -10.535 94.105 ;
        RECT -6.485 93.935 -5.935 94.105 ;
        RECT -5.755 93.865 -5.385 94.205 ;
        RECT -5.205 94.105 -5.035 94.430 ;
        RECT -2.065 94.430 -0.995 94.600 ;
        RECT -2.065 94.105 -1.895 94.430 ;
        RECT -5.205 93.925 -4.275 94.105 ;
        RECT -2.825 93.925 -1.895 94.105 ;
        RECT -1.715 93.865 -1.345 94.205 ;
        RECT -1.165 94.105 -0.995 94.430 ;
        RECT 3.815 94.430 4.885 94.600 ;
        RECT 3.815 94.105 3.985 94.430 ;
        RECT -1.165 93.935 -0.615 94.105 ;
        RECT 3.435 93.935 3.985 94.105 ;
        RECT 4.165 93.865 4.535 94.205 ;
        RECT 4.715 94.105 4.885 94.430 ;
        RECT 7.855 94.430 8.925 94.600 ;
        RECT 7.855 94.105 8.025 94.430 ;
        RECT 4.715 93.925 5.645 94.105 ;
        RECT 7.095 93.925 8.025 94.105 ;
        RECT 8.205 93.865 8.575 94.205 ;
        RECT 8.755 94.105 8.925 94.430 ;
        RECT 13.735 94.430 14.805 94.600 ;
        RECT 13.735 94.105 13.905 94.430 ;
        RECT 8.755 93.935 9.305 94.105 ;
        RECT 13.355 93.935 13.905 94.105 ;
        RECT 14.085 93.865 14.455 94.205 ;
        RECT 14.635 94.105 14.805 94.430 ;
        RECT 17.775 94.430 18.845 94.600 ;
        RECT 17.775 94.105 17.945 94.430 ;
        RECT 14.635 93.925 15.565 94.105 ;
        RECT 17.015 93.925 17.945 94.105 ;
        RECT 18.125 93.865 18.495 94.205 ;
        RECT 18.675 94.105 18.845 94.430 ;
        RECT 23.655 94.430 24.725 94.600 ;
        RECT 23.655 94.105 23.825 94.430 ;
        RECT 18.675 93.935 19.225 94.105 ;
        RECT 23.275 93.935 23.825 94.105 ;
        RECT 24.005 93.865 24.375 94.205 ;
        RECT 24.555 94.105 24.725 94.430 ;
        RECT 24.555 93.925 25.485 94.105 ;
        RECT -291.460 93.245 -289.620 93.415 ;
        RECT 24.600 93.245 26.440 93.415 ;
        RECT -291.375 92.520 -291.085 93.245 ;
        RECT -290.915 92.445 -290.605 93.245 ;
        RECT -290.400 92.445 -289.705 93.075 ;
        RECT -291.375 90.695 -291.085 91.860 ;
        RECT -290.400 91.845 -290.230 92.445 ;
        RECT -290.060 92.005 -289.725 92.255 ;
        RECT -287.365 92.095 -287.035 93.075 ;
        RECT -285.505 92.095 -285.175 93.075 ;
        RECT -282.835 92.445 -282.140 93.075 ;
        RECT -290.915 90.695 -290.635 91.835 ;
        RECT -290.465 90.865 -290.135 91.845 ;
        RECT -289.965 90.695 -289.705 91.835 ;
        RECT -287.775 91.685 -287.440 91.935 ;
        RECT -287.270 91.495 -287.100 92.095 ;
        RECT -287.795 90.865 -287.100 91.495 ;
        RECT -285.440 91.495 -285.270 92.095 ;
        RECT -282.815 92.005 -282.480 92.255 ;
        RECT -285.100 91.685 -284.765 91.935 ;
        RECT -282.310 91.845 -282.140 92.445 ;
        RECT -280.480 92.445 -279.785 93.075 ;
        RECT -280.480 91.845 -280.310 92.445 ;
        RECT -280.140 92.005 -279.805 92.255 ;
        RECT -277.445 92.095 -277.115 93.075 ;
        RECT -275.585 92.095 -275.255 93.075 ;
        RECT -272.915 92.445 -272.220 93.075 ;
        RECT -285.440 90.865 -284.745 91.495 ;
        RECT -282.405 90.865 -282.075 91.845 ;
        RECT -280.545 90.865 -280.215 91.845 ;
        RECT -277.855 91.685 -277.520 91.935 ;
        RECT -277.350 91.495 -277.180 92.095 ;
        RECT -277.875 90.865 -277.180 91.495 ;
        RECT -275.520 91.495 -275.350 92.095 ;
        RECT -272.895 92.005 -272.560 92.255 ;
        RECT -275.180 91.685 -274.845 91.935 ;
        RECT -272.390 91.845 -272.220 92.445 ;
        RECT -270.560 92.445 -269.865 93.075 ;
        RECT -270.560 91.845 -270.390 92.445 ;
        RECT -270.220 92.005 -269.885 92.255 ;
        RECT -267.525 92.095 -267.195 93.075 ;
        RECT -265.665 92.095 -265.335 93.075 ;
        RECT -262.995 92.445 -262.300 93.075 ;
        RECT -275.520 90.865 -274.825 91.495 ;
        RECT -272.485 90.865 -272.155 91.845 ;
        RECT -270.625 90.865 -270.295 91.845 ;
        RECT -267.935 91.685 -267.600 91.935 ;
        RECT -267.430 91.495 -267.260 92.095 ;
        RECT -267.955 90.865 -267.260 91.495 ;
        RECT -265.600 91.495 -265.430 92.095 ;
        RECT -262.975 92.005 -262.640 92.255 ;
        RECT -265.260 91.685 -264.925 91.935 ;
        RECT -262.470 91.845 -262.300 92.445 ;
        RECT -260.640 92.445 -259.945 93.075 ;
        RECT -260.640 91.845 -260.470 92.445 ;
        RECT -260.300 92.005 -259.965 92.255 ;
        RECT -257.605 92.095 -257.275 93.075 ;
        RECT -255.745 92.095 -255.415 93.075 ;
        RECT -253.075 92.445 -252.380 93.075 ;
        RECT -265.600 90.865 -264.905 91.495 ;
        RECT -262.565 90.865 -262.235 91.845 ;
        RECT -260.705 90.865 -260.375 91.845 ;
        RECT -258.015 91.685 -257.680 91.935 ;
        RECT -257.510 91.495 -257.340 92.095 ;
        RECT -258.035 90.865 -257.340 91.495 ;
        RECT -255.680 91.495 -255.510 92.095 ;
        RECT -253.055 92.005 -252.720 92.255 ;
        RECT -255.340 91.685 -255.005 91.935 ;
        RECT -252.550 91.845 -252.380 92.445 ;
        RECT -250.720 92.445 -250.025 93.075 ;
        RECT -250.720 91.845 -250.550 92.445 ;
        RECT -250.380 92.005 -250.045 92.255 ;
        RECT -247.685 92.095 -247.355 93.075 ;
        RECT -245.825 92.095 -245.495 93.075 ;
        RECT -243.155 92.445 -242.460 93.075 ;
        RECT -255.680 90.865 -254.985 91.495 ;
        RECT -252.645 90.865 -252.315 91.845 ;
        RECT -250.785 90.865 -250.455 91.845 ;
        RECT -248.095 91.685 -247.760 91.935 ;
        RECT -247.590 91.495 -247.420 92.095 ;
        RECT -248.115 90.865 -247.420 91.495 ;
        RECT -245.760 91.495 -245.590 92.095 ;
        RECT -243.135 92.005 -242.800 92.255 ;
        RECT -245.420 91.685 -245.085 91.935 ;
        RECT -242.630 91.845 -242.460 92.445 ;
        RECT -240.800 92.445 -240.105 93.075 ;
        RECT -240.800 91.845 -240.630 92.445 ;
        RECT -240.460 92.005 -240.125 92.255 ;
        RECT -237.765 92.095 -237.435 93.075 ;
        RECT -235.905 92.095 -235.575 93.075 ;
        RECT -233.235 92.445 -232.540 93.075 ;
        RECT -245.760 90.865 -245.065 91.495 ;
        RECT -242.725 90.865 -242.395 91.845 ;
        RECT -240.865 90.865 -240.535 91.845 ;
        RECT -238.175 91.685 -237.840 91.935 ;
        RECT -237.670 91.495 -237.500 92.095 ;
        RECT -238.195 90.865 -237.500 91.495 ;
        RECT -235.840 91.495 -235.670 92.095 ;
        RECT -233.215 92.005 -232.880 92.255 ;
        RECT -235.500 91.685 -235.165 91.935 ;
        RECT -232.710 91.845 -232.540 92.445 ;
        RECT -230.880 92.445 -230.185 93.075 ;
        RECT -230.880 91.845 -230.710 92.445 ;
        RECT -230.540 92.005 -230.205 92.255 ;
        RECT -227.845 92.095 -227.515 93.075 ;
        RECT -225.985 92.095 -225.655 93.075 ;
        RECT -223.315 92.445 -222.620 93.075 ;
        RECT -235.840 90.865 -235.145 91.495 ;
        RECT -232.805 90.865 -232.475 91.845 ;
        RECT -230.945 90.865 -230.615 91.845 ;
        RECT -228.255 91.685 -227.920 91.935 ;
        RECT -227.750 91.495 -227.580 92.095 ;
        RECT -228.275 90.865 -227.580 91.495 ;
        RECT -225.920 91.495 -225.750 92.095 ;
        RECT -223.295 92.005 -222.960 92.255 ;
        RECT -225.580 91.685 -225.245 91.935 ;
        RECT -222.790 91.845 -222.620 92.445 ;
        RECT -220.960 92.445 -220.265 93.075 ;
        RECT -220.960 91.845 -220.790 92.445 ;
        RECT -220.620 92.005 -220.285 92.255 ;
        RECT -217.925 92.095 -217.595 93.075 ;
        RECT -216.065 92.095 -215.735 93.075 ;
        RECT -213.395 92.445 -212.700 93.075 ;
        RECT -225.920 90.865 -225.225 91.495 ;
        RECT -222.885 90.865 -222.555 91.845 ;
        RECT -221.025 90.865 -220.695 91.845 ;
        RECT -218.335 91.685 -218.000 91.935 ;
        RECT -217.830 91.495 -217.660 92.095 ;
        RECT -218.355 90.865 -217.660 91.495 ;
        RECT -216.000 91.495 -215.830 92.095 ;
        RECT -213.375 92.005 -213.040 92.255 ;
        RECT -215.660 91.685 -215.325 91.935 ;
        RECT -212.870 91.845 -212.700 92.445 ;
        RECT -211.040 92.445 -210.345 93.075 ;
        RECT -211.040 91.845 -210.870 92.445 ;
        RECT -210.700 92.005 -210.365 92.255 ;
        RECT -208.005 92.095 -207.675 93.075 ;
        RECT -206.145 92.095 -205.815 93.075 ;
        RECT -203.475 92.445 -202.780 93.075 ;
        RECT -216.000 90.865 -215.305 91.495 ;
        RECT -212.965 90.865 -212.635 91.845 ;
        RECT -211.105 90.865 -210.775 91.845 ;
        RECT -208.415 91.685 -208.080 91.935 ;
        RECT -207.910 91.495 -207.740 92.095 ;
        RECT -208.435 90.865 -207.740 91.495 ;
        RECT -206.080 91.495 -205.910 92.095 ;
        RECT -203.455 92.005 -203.120 92.255 ;
        RECT -205.740 91.685 -205.405 91.935 ;
        RECT -202.950 91.845 -202.780 92.445 ;
        RECT -201.120 92.445 -200.425 93.075 ;
        RECT -201.120 91.845 -200.950 92.445 ;
        RECT -200.780 92.005 -200.445 92.255 ;
        RECT -198.085 92.095 -197.755 93.075 ;
        RECT -196.225 92.095 -195.895 93.075 ;
        RECT -193.555 92.445 -192.860 93.075 ;
        RECT -206.080 90.865 -205.385 91.495 ;
        RECT -203.045 90.865 -202.715 91.845 ;
        RECT -201.185 90.865 -200.855 91.845 ;
        RECT -198.495 91.685 -198.160 91.935 ;
        RECT -197.990 91.495 -197.820 92.095 ;
        RECT -198.515 90.865 -197.820 91.495 ;
        RECT -196.160 91.495 -195.990 92.095 ;
        RECT -193.535 92.005 -193.200 92.255 ;
        RECT -195.820 91.685 -195.485 91.935 ;
        RECT -193.030 91.845 -192.860 92.445 ;
        RECT -191.200 92.445 -190.505 93.075 ;
        RECT -191.200 91.845 -191.030 92.445 ;
        RECT -190.860 92.005 -190.525 92.255 ;
        RECT -188.165 92.095 -187.835 93.075 ;
        RECT -186.305 92.095 -185.975 93.075 ;
        RECT -183.635 92.445 -182.940 93.075 ;
        RECT -196.160 90.865 -195.465 91.495 ;
        RECT -193.125 90.865 -192.795 91.845 ;
        RECT -191.265 90.865 -190.935 91.845 ;
        RECT -188.575 91.685 -188.240 91.935 ;
        RECT -188.070 91.495 -187.900 92.095 ;
        RECT -188.595 90.865 -187.900 91.495 ;
        RECT -186.240 91.495 -186.070 92.095 ;
        RECT -183.615 92.005 -183.280 92.255 ;
        RECT -185.900 91.685 -185.565 91.935 ;
        RECT -183.110 91.845 -182.940 92.445 ;
        RECT -181.280 92.445 -180.585 93.075 ;
        RECT -181.280 91.845 -181.110 92.445 ;
        RECT -180.940 92.005 -180.605 92.255 ;
        RECT -178.245 92.095 -177.915 93.075 ;
        RECT -176.385 92.095 -176.055 93.075 ;
        RECT -173.715 92.445 -173.020 93.075 ;
        RECT -186.240 90.865 -185.545 91.495 ;
        RECT -183.205 90.865 -182.875 91.845 ;
        RECT -181.345 90.865 -181.015 91.845 ;
        RECT -178.655 91.685 -178.320 91.935 ;
        RECT -178.150 91.495 -177.980 92.095 ;
        RECT -178.675 90.865 -177.980 91.495 ;
        RECT -176.320 91.495 -176.150 92.095 ;
        RECT -173.695 92.005 -173.360 92.255 ;
        RECT -175.980 91.685 -175.645 91.935 ;
        RECT -173.190 91.845 -173.020 92.445 ;
        RECT -171.360 92.445 -170.665 93.075 ;
        RECT -171.360 91.845 -171.190 92.445 ;
        RECT -171.020 92.005 -170.685 92.255 ;
        RECT -168.325 92.095 -167.995 93.075 ;
        RECT -166.465 92.095 -166.135 93.075 ;
        RECT -163.795 92.445 -163.100 93.075 ;
        RECT -176.320 90.865 -175.625 91.495 ;
        RECT -173.285 90.865 -172.955 91.845 ;
        RECT -171.425 90.865 -171.095 91.845 ;
        RECT -168.735 91.685 -168.400 91.935 ;
        RECT -168.230 91.495 -168.060 92.095 ;
        RECT -168.755 90.865 -168.060 91.495 ;
        RECT -166.400 91.495 -166.230 92.095 ;
        RECT -163.775 92.005 -163.440 92.255 ;
        RECT -166.060 91.685 -165.725 91.935 ;
        RECT -163.270 91.845 -163.100 92.445 ;
        RECT -161.440 92.445 -160.745 93.075 ;
        RECT -161.440 91.845 -161.270 92.445 ;
        RECT -161.100 92.005 -160.765 92.255 ;
        RECT -158.405 92.095 -158.075 93.075 ;
        RECT -156.545 92.095 -156.215 93.075 ;
        RECT -153.875 92.445 -153.180 93.075 ;
        RECT -166.400 90.865 -165.705 91.495 ;
        RECT -163.365 90.865 -163.035 91.845 ;
        RECT -161.505 90.865 -161.175 91.845 ;
        RECT -158.815 91.685 -158.480 91.935 ;
        RECT -158.310 91.495 -158.140 92.095 ;
        RECT -158.835 90.865 -158.140 91.495 ;
        RECT -156.480 91.495 -156.310 92.095 ;
        RECT -153.855 92.005 -153.520 92.255 ;
        RECT -156.140 91.685 -155.805 91.935 ;
        RECT -153.350 91.845 -153.180 92.445 ;
        RECT -151.520 92.445 -150.825 93.075 ;
        RECT -151.520 91.845 -151.350 92.445 ;
        RECT -151.180 92.005 -150.845 92.255 ;
        RECT -148.485 92.095 -148.155 93.075 ;
        RECT -146.625 92.095 -146.295 93.075 ;
        RECT -143.955 92.445 -143.260 93.075 ;
        RECT -156.480 90.865 -155.785 91.495 ;
        RECT -153.445 90.865 -153.115 91.845 ;
        RECT -151.585 90.865 -151.255 91.845 ;
        RECT -148.895 91.685 -148.560 91.935 ;
        RECT -148.390 91.495 -148.220 92.095 ;
        RECT -148.915 90.865 -148.220 91.495 ;
        RECT -146.560 91.495 -146.390 92.095 ;
        RECT -143.935 92.005 -143.600 92.255 ;
        RECT -146.220 91.685 -145.885 91.935 ;
        RECT -143.430 91.845 -143.260 92.445 ;
        RECT -141.600 92.445 -140.905 93.075 ;
        RECT -141.600 91.845 -141.430 92.445 ;
        RECT -141.260 92.005 -140.925 92.255 ;
        RECT -138.565 92.095 -138.235 93.075 ;
        RECT -136.705 92.095 -136.375 93.075 ;
        RECT -134.035 92.445 -133.340 93.075 ;
        RECT -146.560 90.865 -145.865 91.495 ;
        RECT -143.525 90.865 -143.195 91.845 ;
        RECT -141.665 90.865 -141.335 91.845 ;
        RECT -138.975 91.685 -138.640 91.935 ;
        RECT -138.470 91.495 -138.300 92.095 ;
        RECT -138.995 90.865 -138.300 91.495 ;
        RECT -136.640 91.495 -136.470 92.095 ;
        RECT -134.015 92.005 -133.680 92.255 ;
        RECT -136.300 91.685 -135.965 91.935 ;
        RECT -133.510 91.845 -133.340 92.445 ;
        RECT -131.680 92.445 -130.985 93.075 ;
        RECT -131.680 91.845 -131.510 92.445 ;
        RECT -131.340 92.005 -131.005 92.255 ;
        RECT -128.645 92.095 -128.315 93.075 ;
        RECT -126.785 92.095 -126.455 93.075 ;
        RECT -124.115 92.445 -123.420 93.075 ;
        RECT -136.640 90.865 -135.945 91.495 ;
        RECT -133.605 90.865 -133.275 91.845 ;
        RECT -131.745 90.865 -131.415 91.845 ;
        RECT -129.055 91.685 -128.720 91.935 ;
        RECT -128.550 91.495 -128.380 92.095 ;
        RECT -129.075 90.865 -128.380 91.495 ;
        RECT -126.720 91.495 -126.550 92.095 ;
        RECT -124.095 92.005 -123.760 92.255 ;
        RECT -126.380 91.685 -126.045 91.935 ;
        RECT -123.590 91.845 -123.420 92.445 ;
        RECT -121.760 92.445 -121.065 93.075 ;
        RECT -121.760 91.845 -121.590 92.445 ;
        RECT -121.420 92.005 -121.085 92.255 ;
        RECT -118.725 92.095 -118.395 93.075 ;
        RECT -116.865 92.095 -116.535 93.075 ;
        RECT -114.195 92.445 -113.500 93.075 ;
        RECT -126.720 90.865 -126.025 91.495 ;
        RECT -123.685 90.865 -123.355 91.845 ;
        RECT -121.825 90.865 -121.495 91.845 ;
        RECT -119.135 91.685 -118.800 91.935 ;
        RECT -118.630 91.495 -118.460 92.095 ;
        RECT -119.155 90.865 -118.460 91.495 ;
        RECT -116.800 91.495 -116.630 92.095 ;
        RECT -114.175 92.005 -113.840 92.255 ;
        RECT -116.460 91.685 -116.125 91.935 ;
        RECT -113.670 91.845 -113.500 92.445 ;
        RECT -111.840 92.445 -111.145 93.075 ;
        RECT -111.840 91.845 -111.670 92.445 ;
        RECT -111.500 92.005 -111.165 92.255 ;
        RECT -108.805 92.095 -108.475 93.075 ;
        RECT -106.945 92.095 -106.615 93.075 ;
        RECT -104.275 92.445 -103.580 93.075 ;
        RECT -116.800 90.865 -116.105 91.495 ;
        RECT -113.765 90.865 -113.435 91.845 ;
        RECT -111.905 90.865 -111.575 91.845 ;
        RECT -109.215 91.685 -108.880 91.935 ;
        RECT -108.710 91.495 -108.540 92.095 ;
        RECT -109.235 90.865 -108.540 91.495 ;
        RECT -106.880 91.495 -106.710 92.095 ;
        RECT -104.255 92.005 -103.920 92.255 ;
        RECT -106.540 91.685 -106.205 91.935 ;
        RECT -103.750 91.845 -103.580 92.445 ;
        RECT -101.920 92.445 -101.225 93.075 ;
        RECT -101.920 91.845 -101.750 92.445 ;
        RECT -101.580 92.005 -101.245 92.255 ;
        RECT -98.885 92.095 -98.555 93.075 ;
        RECT -97.025 92.095 -96.695 93.075 ;
        RECT -94.355 92.445 -93.660 93.075 ;
        RECT -106.880 90.865 -106.185 91.495 ;
        RECT -103.845 90.865 -103.515 91.845 ;
        RECT -101.985 90.865 -101.655 91.845 ;
        RECT -99.295 91.685 -98.960 91.935 ;
        RECT -98.790 91.495 -98.620 92.095 ;
        RECT -99.315 90.865 -98.620 91.495 ;
        RECT -96.960 91.495 -96.790 92.095 ;
        RECT -94.335 92.005 -94.000 92.255 ;
        RECT -96.620 91.685 -96.285 91.935 ;
        RECT -93.830 91.845 -93.660 92.445 ;
        RECT -92.000 92.445 -91.305 93.075 ;
        RECT -92.000 91.845 -91.830 92.445 ;
        RECT -91.660 92.005 -91.325 92.255 ;
        RECT -88.965 92.095 -88.635 93.075 ;
        RECT -87.105 92.095 -86.775 93.075 ;
        RECT -84.435 92.445 -83.740 93.075 ;
        RECT -96.960 90.865 -96.265 91.495 ;
        RECT -93.925 90.865 -93.595 91.845 ;
        RECT -92.065 90.865 -91.735 91.845 ;
        RECT -89.375 91.685 -89.040 91.935 ;
        RECT -88.870 91.495 -88.700 92.095 ;
        RECT -89.395 90.865 -88.700 91.495 ;
        RECT -87.040 91.495 -86.870 92.095 ;
        RECT -84.415 92.005 -84.080 92.255 ;
        RECT -86.700 91.685 -86.365 91.935 ;
        RECT -83.910 91.845 -83.740 92.445 ;
        RECT -82.080 92.445 -81.385 93.075 ;
        RECT -82.080 91.845 -81.910 92.445 ;
        RECT -81.740 92.005 -81.405 92.255 ;
        RECT -79.045 92.095 -78.715 93.075 ;
        RECT -77.185 92.095 -76.855 93.075 ;
        RECT -74.515 92.445 -73.820 93.075 ;
        RECT -87.040 90.865 -86.345 91.495 ;
        RECT -84.005 90.865 -83.675 91.845 ;
        RECT -82.145 90.865 -81.815 91.845 ;
        RECT -79.455 91.685 -79.120 91.935 ;
        RECT -78.950 91.495 -78.780 92.095 ;
        RECT -79.475 90.865 -78.780 91.495 ;
        RECT -77.120 91.495 -76.950 92.095 ;
        RECT -74.495 92.005 -74.160 92.255 ;
        RECT -76.780 91.685 -76.445 91.935 ;
        RECT -73.990 91.845 -73.820 92.445 ;
        RECT -72.160 92.445 -71.465 93.075 ;
        RECT -72.160 91.845 -71.990 92.445 ;
        RECT -71.820 92.005 -71.485 92.255 ;
        RECT -69.125 92.095 -68.795 93.075 ;
        RECT -67.265 92.095 -66.935 93.075 ;
        RECT -64.595 92.445 -63.900 93.075 ;
        RECT -77.120 90.865 -76.425 91.495 ;
        RECT -74.085 90.865 -73.755 91.845 ;
        RECT -72.225 90.865 -71.895 91.845 ;
        RECT -69.535 91.685 -69.200 91.935 ;
        RECT -69.030 91.495 -68.860 92.095 ;
        RECT -69.555 90.865 -68.860 91.495 ;
        RECT -67.200 91.495 -67.030 92.095 ;
        RECT -64.575 92.005 -64.240 92.255 ;
        RECT -66.860 91.685 -66.525 91.935 ;
        RECT -64.070 91.845 -63.900 92.445 ;
        RECT -62.240 92.445 -61.545 93.075 ;
        RECT -62.240 91.845 -62.070 92.445 ;
        RECT -61.900 92.005 -61.565 92.255 ;
        RECT -59.205 92.095 -58.875 93.075 ;
        RECT -57.345 92.095 -57.015 93.075 ;
        RECT -54.675 92.445 -53.980 93.075 ;
        RECT -67.200 90.865 -66.505 91.495 ;
        RECT -64.165 90.865 -63.835 91.845 ;
        RECT -62.305 90.865 -61.975 91.845 ;
        RECT -59.615 91.685 -59.280 91.935 ;
        RECT -59.110 91.495 -58.940 92.095 ;
        RECT -59.635 90.865 -58.940 91.495 ;
        RECT -57.280 91.495 -57.110 92.095 ;
        RECT -54.655 92.005 -54.320 92.255 ;
        RECT -56.940 91.685 -56.605 91.935 ;
        RECT -54.150 91.845 -53.980 92.445 ;
        RECT -52.320 92.445 -51.625 93.075 ;
        RECT -52.320 91.845 -52.150 92.445 ;
        RECT -51.980 92.005 -51.645 92.255 ;
        RECT -49.285 92.095 -48.955 93.075 ;
        RECT -47.425 92.095 -47.095 93.075 ;
        RECT -44.755 92.445 -44.060 93.075 ;
        RECT -57.280 90.865 -56.585 91.495 ;
        RECT -54.245 90.865 -53.915 91.845 ;
        RECT -52.385 90.865 -52.055 91.845 ;
        RECT -49.695 91.685 -49.360 91.935 ;
        RECT -49.190 91.495 -49.020 92.095 ;
        RECT -49.715 90.865 -49.020 91.495 ;
        RECT -47.360 91.495 -47.190 92.095 ;
        RECT -44.735 92.005 -44.400 92.255 ;
        RECT -47.020 91.685 -46.685 91.935 ;
        RECT -44.230 91.845 -44.060 92.445 ;
        RECT -42.400 92.445 -41.705 93.075 ;
        RECT -42.400 91.845 -42.230 92.445 ;
        RECT -42.060 92.005 -41.725 92.255 ;
        RECT -39.365 92.095 -39.035 93.075 ;
        RECT -37.505 92.095 -37.175 93.075 ;
        RECT -34.835 92.445 -34.140 93.075 ;
        RECT -47.360 90.865 -46.665 91.495 ;
        RECT -44.325 90.865 -43.995 91.845 ;
        RECT -42.465 90.865 -42.135 91.845 ;
        RECT -39.775 91.685 -39.440 91.935 ;
        RECT -39.270 91.495 -39.100 92.095 ;
        RECT -39.795 90.865 -39.100 91.495 ;
        RECT -37.440 91.495 -37.270 92.095 ;
        RECT -34.815 92.005 -34.480 92.255 ;
        RECT -37.100 91.685 -36.765 91.935 ;
        RECT -34.310 91.845 -34.140 92.445 ;
        RECT -32.480 92.445 -31.785 93.075 ;
        RECT -32.480 91.845 -32.310 92.445 ;
        RECT -32.140 92.005 -31.805 92.255 ;
        RECT -29.445 92.095 -29.115 93.075 ;
        RECT -27.585 92.095 -27.255 93.075 ;
        RECT -24.915 92.445 -24.220 93.075 ;
        RECT -37.440 90.865 -36.745 91.495 ;
        RECT -34.405 90.865 -34.075 91.845 ;
        RECT -32.545 90.865 -32.215 91.845 ;
        RECT -29.855 91.685 -29.520 91.935 ;
        RECT -29.350 91.495 -29.180 92.095 ;
        RECT -29.875 90.865 -29.180 91.495 ;
        RECT -27.520 91.495 -27.350 92.095 ;
        RECT -24.895 92.005 -24.560 92.255 ;
        RECT -27.180 91.685 -26.845 91.935 ;
        RECT -24.390 91.845 -24.220 92.445 ;
        RECT -22.560 92.445 -21.865 93.075 ;
        RECT -22.560 91.845 -22.390 92.445 ;
        RECT -22.220 92.005 -21.885 92.255 ;
        RECT -19.525 92.095 -19.195 93.075 ;
        RECT -17.665 92.095 -17.335 93.075 ;
        RECT -14.995 92.445 -14.300 93.075 ;
        RECT -27.520 90.865 -26.825 91.495 ;
        RECT -24.485 90.865 -24.155 91.845 ;
        RECT -22.625 90.865 -22.295 91.845 ;
        RECT -19.935 91.685 -19.600 91.935 ;
        RECT -19.430 91.495 -19.260 92.095 ;
        RECT -19.955 90.865 -19.260 91.495 ;
        RECT -17.600 91.495 -17.430 92.095 ;
        RECT -14.975 92.005 -14.640 92.255 ;
        RECT -17.260 91.685 -16.925 91.935 ;
        RECT -14.470 91.845 -14.300 92.445 ;
        RECT -12.640 92.445 -11.945 93.075 ;
        RECT -12.640 91.845 -12.470 92.445 ;
        RECT -12.300 92.005 -11.965 92.255 ;
        RECT -9.605 92.095 -9.275 93.075 ;
        RECT -7.745 92.095 -7.415 93.075 ;
        RECT -5.075 92.445 -4.380 93.075 ;
        RECT -17.600 90.865 -16.905 91.495 ;
        RECT -14.565 90.865 -14.235 91.845 ;
        RECT -12.705 90.865 -12.375 91.845 ;
        RECT -10.015 91.685 -9.680 91.935 ;
        RECT -9.510 91.495 -9.340 92.095 ;
        RECT -10.035 90.865 -9.340 91.495 ;
        RECT -7.680 91.495 -7.510 92.095 ;
        RECT -5.055 92.005 -4.720 92.255 ;
        RECT -7.340 91.685 -7.005 91.935 ;
        RECT -4.550 91.845 -4.380 92.445 ;
        RECT -2.720 92.445 -2.025 93.075 ;
        RECT -2.720 91.845 -2.550 92.445 ;
        RECT -2.380 92.005 -2.045 92.255 ;
        RECT 0.315 92.095 0.645 93.075 ;
        RECT 2.175 92.095 2.505 93.075 ;
        RECT 4.845 92.445 5.540 93.075 ;
        RECT -7.680 90.865 -6.985 91.495 ;
        RECT -4.645 90.865 -4.315 91.845 ;
        RECT -2.785 90.865 -2.455 91.845 ;
        RECT -0.095 91.685 0.240 91.935 ;
        RECT 0.410 91.495 0.580 92.095 ;
        RECT -0.115 90.865 0.580 91.495 ;
        RECT 2.240 91.495 2.410 92.095 ;
        RECT 4.865 92.005 5.200 92.255 ;
        RECT 2.580 91.685 2.915 91.935 ;
        RECT 5.370 91.845 5.540 92.445 ;
        RECT 7.200 92.445 7.895 93.075 ;
        RECT 7.200 91.845 7.370 92.445 ;
        RECT 7.540 92.005 7.875 92.255 ;
        RECT 10.235 92.095 10.565 93.075 ;
        RECT 12.095 92.095 12.425 93.075 ;
        RECT 14.765 92.445 15.460 93.075 ;
        RECT 2.240 90.865 2.935 91.495 ;
        RECT 5.275 90.865 5.605 91.845 ;
        RECT 7.135 90.865 7.465 91.845 ;
        RECT 9.825 91.685 10.160 91.935 ;
        RECT 10.330 91.495 10.500 92.095 ;
        RECT 9.805 90.865 10.500 91.495 ;
        RECT 12.160 91.495 12.330 92.095 ;
        RECT 14.785 92.005 15.120 92.255 ;
        RECT 12.500 91.685 12.835 91.935 ;
        RECT 15.290 91.845 15.460 92.445 ;
        RECT 17.120 92.445 17.815 93.075 ;
        RECT 17.120 91.845 17.290 92.445 ;
        RECT 17.460 92.005 17.795 92.255 ;
        RECT 20.155 92.095 20.485 93.075 ;
        RECT 22.015 92.095 22.345 93.075 ;
        RECT 24.685 92.445 25.380 93.075 ;
        RECT 25.585 92.445 25.895 93.245 ;
        RECT 26.065 92.520 26.355 93.245 ;
        RECT 12.160 90.865 12.855 91.495 ;
        RECT 15.195 90.865 15.525 91.845 ;
        RECT 17.055 90.865 17.385 91.845 ;
        RECT 19.745 91.685 20.080 91.935 ;
        RECT 20.250 91.495 20.420 92.095 ;
        RECT 19.725 90.865 20.420 91.495 ;
        RECT 22.080 91.495 22.250 92.095 ;
        RECT 24.705 92.005 25.040 92.255 ;
        RECT 22.420 91.685 22.755 91.935 ;
        RECT 25.210 91.845 25.380 92.445 ;
        RECT 22.080 90.865 22.775 91.495 ;
        RECT 25.115 90.865 25.445 91.845 ;
        RECT -291.460 90.525 -289.620 90.695 ;
        RECT -290.075 89.140 -289.785 89.850 ;
        RECT -289.545 89.655 -289.375 90.180 ;
        RECT -289.205 89.835 -288.655 90.005 ;
        RECT -289.545 89.325 -288.995 89.655 ;
        RECT -288.825 89.510 -288.655 89.835 ;
        RECT -288.475 89.735 -288.105 90.075 ;
        RECT -287.925 89.835 -286.995 90.015 ;
        RECT -285.545 89.835 -284.615 90.015 ;
        RECT -287.925 89.510 -287.755 89.835 ;
        RECT -288.825 89.340 -287.755 89.510 ;
        RECT -284.785 89.510 -284.615 89.835 ;
        RECT -284.435 89.735 -284.065 90.075 ;
        RECT -283.885 89.835 -283.335 90.005 ;
        RECT -279.285 89.835 -278.735 90.005 ;
        RECT -283.885 89.510 -283.715 89.835 ;
        RECT -284.785 89.340 -283.715 89.510 ;
        RECT -278.905 89.510 -278.735 89.835 ;
        RECT -278.555 89.735 -278.185 90.075 ;
        RECT -278.005 89.835 -277.075 90.015 ;
        RECT -275.625 89.835 -274.695 90.015 ;
        RECT -278.005 89.510 -277.835 89.835 ;
        RECT -278.905 89.340 -277.835 89.510 ;
        RECT -274.865 89.510 -274.695 89.835 ;
        RECT -274.515 89.735 -274.145 90.075 ;
        RECT -273.965 89.835 -273.415 90.005 ;
        RECT -269.365 89.835 -268.815 90.005 ;
        RECT -273.965 89.510 -273.795 89.835 ;
        RECT -274.865 89.340 -273.795 89.510 ;
        RECT -268.985 89.510 -268.815 89.835 ;
        RECT -268.635 89.735 -268.265 90.075 ;
        RECT -268.085 89.835 -267.155 90.015 ;
        RECT -265.705 89.835 -264.775 90.015 ;
        RECT -268.085 89.510 -267.915 89.835 ;
        RECT -268.985 89.340 -267.915 89.510 ;
        RECT -264.945 89.510 -264.775 89.835 ;
        RECT -264.595 89.735 -264.225 90.075 ;
        RECT -264.045 89.835 -263.495 90.005 ;
        RECT -259.445 89.835 -258.895 90.005 ;
        RECT -264.045 89.510 -263.875 89.835 ;
        RECT -264.945 89.340 -263.875 89.510 ;
        RECT -259.065 89.510 -258.895 89.835 ;
        RECT -258.715 89.735 -258.345 90.075 ;
        RECT -258.165 89.835 -257.235 90.015 ;
        RECT -255.785 89.835 -254.855 90.015 ;
        RECT -258.165 89.510 -257.995 89.835 ;
        RECT -259.065 89.340 -257.995 89.510 ;
        RECT -255.025 89.510 -254.855 89.835 ;
        RECT -254.675 89.735 -254.305 90.075 ;
        RECT -254.125 89.835 -253.575 90.005 ;
        RECT -249.525 89.835 -248.975 90.005 ;
        RECT -254.125 89.510 -253.955 89.835 ;
        RECT -255.025 89.340 -253.955 89.510 ;
        RECT -249.145 89.510 -248.975 89.835 ;
        RECT -248.795 89.735 -248.425 90.075 ;
        RECT -248.245 89.835 -247.315 90.015 ;
        RECT -245.865 89.835 -244.935 90.015 ;
        RECT -248.245 89.510 -248.075 89.835 ;
        RECT -249.145 89.340 -248.075 89.510 ;
        RECT -245.105 89.510 -244.935 89.835 ;
        RECT -244.755 89.735 -244.385 90.075 ;
        RECT -244.205 89.835 -243.655 90.005 ;
        RECT -239.605 89.835 -239.055 90.005 ;
        RECT -244.205 89.510 -244.035 89.835 ;
        RECT -245.105 89.340 -244.035 89.510 ;
        RECT -239.225 89.510 -239.055 89.835 ;
        RECT -238.875 89.735 -238.505 90.075 ;
        RECT -238.325 89.835 -237.395 90.015 ;
        RECT -235.945 89.835 -235.015 90.015 ;
        RECT -238.325 89.510 -238.155 89.835 ;
        RECT -239.225 89.340 -238.155 89.510 ;
        RECT -235.185 89.510 -235.015 89.835 ;
        RECT -234.835 89.735 -234.465 90.075 ;
        RECT -234.285 89.835 -233.735 90.005 ;
        RECT -229.685 89.835 -229.135 90.005 ;
        RECT -234.285 89.510 -234.115 89.835 ;
        RECT -235.185 89.340 -234.115 89.510 ;
        RECT -229.305 89.510 -229.135 89.835 ;
        RECT -228.955 89.735 -228.585 90.075 ;
        RECT -228.405 89.835 -227.475 90.015 ;
        RECT -226.025 89.835 -225.095 90.015 ;
        RECT -228.405 89.510 -228.235 89.835 ;
        RECT -229.305 89.340 -228.235 89.510 ;
        RECT -225.265 89.510 -225.095 89.835 ;
        RECT -224.915 89.735 -224.545 90.075 ;
        RECT -224.365 89.835 -223.815 90.005 ;
        RECT -219.765 89.835 -219.215 90.005 ;
        RECT -224.365 89.510 -224.195 89.835 ;
        RECT -225.265 89.340 -224.195 89.510 ;
        RECT -219.385 89.510 -219.215 89.835 ;
        RECT -219.035 89.735 -218.665 90.075 ;
        RECT -218.485 89.835 -217.555 90.015 ;
        RECT -216.105 89.835 -215.175 90.015 ;
        RECT -218.485 89.510 -218.315 89.835 ;
        RECT -219.385 89.340 -218.315 89.510 ;
        RECT -215.345 89.510 -215.175 89.835 ;
        RECT -214.995 89.735 -214.625 90.075 ;
        RECT -214.445 89.835 -213.895 90.005 ;
        RECT -209.845 89.835 -209.295 90.005 ;
        RECT -214.445 89.510 -214.275 89.835 ;
        RECT -215.345 89.340 -214.275 89.510 ;
        RECT -209.465 89.510 -209.295 89.835 ;
        RECT -209.115 89.735 -208.745 90.075 ;
        RECT -208.565 89.835 -207.635 90.015 ;
        RECT -206.185 89.835 -205.255 90.015 ;
        RECT -208.565 89.510 -208.395 89.835 ;
        RECT -209.465 89.340 -208.395 89.510 ;
        RECT -205.425 89.510 -205.255 89.835 ;
        RECT -205.075 89.735 -204.705 90.075 ;
        RECT -204.525 89.835 -203.975 90.005 ;
        RECT -199.925 89.835 -199.375 90.005 ;
        RECT -204.525 89.510 -204.355 89.835 ;
        RECT -205.425 89.340 -204.355 89.510 ;
        RECT -199.545 89.510 -199.375 89.835 ;
        RECT -199.195 89.735 -198.825 90.075 ;
        RECT -198.645 89.835 -197.715 90.015 ;
        RECT -196.265 89.835 -195.335 90.015 ;
        RECT -198.645 89.510 -198.475 89.835 ;
        RECT -199.545 89.340 -198.475 89.510 ;
        RECT -195.505 89.510 -195.335 89.835 ;
        RECT -195.155 89.735 -194.785 90.075 ;
        RECT -194.605 89.835 -194.055 90.005 ;
        RECT -190.005 89.835 -189.455 90.005 ;
        RECT -194.605 89.510 -194.435 89.835 ;
        RECT -195.505 89.340 -194.435 89.510 ;
        RECT -189.625 89.510 -189.455 89.835 ;
        RECT -189.275 89.735 -188.905 90.075 ;
        RECT -188.725 89.835 -187.795 90.015 ;
        RECT -186.345 89.835 -185.415 90.015 ;
        RECT -188.725 89.510 -188.555 89.835 ;
        RECT -189.625 89.340 -188.555 89.510 ;
        RECT -185.585 89.510 -185.415 89.835 ;
        RECT -185.235 89.735 -184.865 90.075 ;
        RECT -184.685 89.835 -184.135 90.005 ;
        RECT -180.085 89.835 -179.535 90.005 ;
        RECT -184.685 89.510 -184.515 89.835 ;
        RECT -185.585 89.340 -184.515 89.510 ;
        RECT -179.705 89.510 -179.535 89.835 ;
        RECT -179.355 89.735 -178.985 90.075 ;
        RECT -178.805 89.835 -177.875 90.015 ;
        RECT -176.425 89.835 -175.495 90.015 ;
        RECT -178.805 89.510 -178.635 89.835 ;
        RECT -179.705 89.340 -178.635 89.510 ;
        RECT -175.665 89.510 -175.495 89.835 ;
        RECT -175.315 89.735 -174.945 90.075 ;
        RECT -174.765 89.835 -174.215 90.005 ;
        RECT -170.165 89.835 -169.615 90.005 ;
        RECT -174.765 89.510 -174.595 89.835 ;
        RECT -175.665 89.340 -174.595 89.510 ;
        RECT -169.785 89.510 -169.615 89.835 ;
        RECT -169.435 89.735 -169.065 90.075 ;
        RECT -168.885 89.835 -167.955 90.015 ;
        RECT -166.505 89.835 -165.575 90.015 ;
        RECT -168.885 89.510 -168.715 89.835 ;
        RECT -169.785 89.340 -168.715 89.510 ;
        RECT -165.745 89.510 -165.575 89.835 ;
        RECT -165.395 89.735 -165.025 90.075 ;
        RECT -164.845 89.835 -164.295 90.005 ;
        RECT -160.245 89.835 -159.695 90.005 ;
        RECT -164.845 89.510 -164.675 89.835 ;
        RECT -165.745 89.340 -164.675 89.510 ;
        RECT -159.865 89.510 -159.695 89.835 ;
        RECT -159.515 89.735 -159.145 90.075 ;
        RECT -158.965 89.835 -158.035 90.015 ;
        RECT -156.585 89.835 -155.655 90.015 ;
        RECT -158.965 89.510 -158.795 89.835 ;
        RECT -159.865 89.340 -158.795 89.510 ;
        RECT -155.825 89.510 -155.655 89.835 ;
        RECT -155.475 89.735 -155.105 90.075 ;
        RECT -154.925 89.835 -154.375 90.005 ;
        RECT -150.325 89.835 -149.775 90.005 ;
        RECT -154.925 89.510 -154.755 89.835 ;
        RECT -155.825 89.340 -154.755 89.510 ;
        RECT -149.945 89.510 -149.775 89.835 ;
        RECT -149.595 89.735 -149.225 90.075 ;
        RECT -149.045 89.835 -148.115 90.015 ;
        RECT -146.665 89.835 -145.735 90.015 ;
        RECT -149.045 89.510 -148.875 89.835 ;
        RECT -149.945 89.340 -148.875 89.510 ;
        RECT -145.905 89.510 -145.735 89.835 ;
        RECT -145.555 89.735 -145.185 90.075 ;
        RECT -145.005 89.835 -144.455 90.005 ;
        RECT -140.405 89.835 -139.855 90.005 ;
        RECT -145.005 89.510 -144.835 89.835 ;
        RECT -145.905 89.340 -144.835 89.510 ;
        RECT -140.025 89.510 -139.855 89.835 ;
        RECT -139.675 89.735 -139.305 90.075 ;
        RECT -139.125 89.835 -138.195 90.015 ;
        RECT -136.745 89.835 -135.815 90.015 ;
        RECT -139.125 89.510 -138.955 89.835 ;
        RECT -140.025 89.340 -138.955 89.510 ;
        RECT -135.985 89.510 -135.815 89.835 ;
        RECT -135.635 89.735 -135.265 90.075 ;
        RECT -135.085 89.835 -134.535 90.005 ;
        RECT -130.485 89.835 -129.935 90.005 ;
        RECT -135.085 89.510 -134.915 89.835 ;
        RECT -135.985 89.340 -134.915 89.510 ;
        RECT -130.105 89.510 -129.935 89.835 ;
        RECT -129.755 89.735 -129.385 90.075 ;
        RECT -129.205 89.835 -128.275 90.015 ;
        RECT -126.825 89.835 -125.895 90.015 ;
        RECT -129.205 89.510 -129.035 89.835 ;
        RECT -130.105 89.340 -129.035 89.510 ;
        RECT -126.065 89.510 -125.895 89.835 ;
        RECT -125.715 89.735 -125.345 90.075 ;
        RECT -125.165 89.835 -124.615 90.005 ;
        RECT -120.565 89.835 -120.015 90.005 ;
        RECT -125.165 89.510 -124.995 89.835 ;
        RECT -126.065 89.340 -124.995 89.510 ;
        RECT -120.185 89.510 -120.015 89.835 ;
        RECT -119.835 89.735 -119.465 90.075 ;
        RECT -119.285 89.835 -118.355 90.015 ;
        RECT -116.905 89.835 -115.975 90.015 ;
        RECT -119.285 89.510 -119.115 89.835 ;
        RECT -120.185 89.340 -119.115 89.510 ;
        RECT -116.145 89.510 -115.975 89.835 ;
        RECT -115.795 89.735 -115.425 90.075 ;
        RECT -115.245 89.835 -114.695 90.005 ;
        RECT -110.645 89.835 -110.095 90.005 ;
        RECT -115.245 89.510 -115.075 89.835 ;
        RECT -116.145 89.340 -115.075 89.510 ;
        RECT -110.265 89.510 -110.095 89.835 ;
        RECT -109.915 89.735 -109.545 90.075 ;
        RECT -109.365 89.835 -108.435 90.015 ;
        RECT -106.985 89.835 -106.055 90.015 ;
        RECT -109.365 89.510 -109.195 89.835 ;
        RECT -110.265 89.340 -109.195 89.510 ;
        RECT -106.225 89.510 -106.055 89.835 ;
        RECT -105.875 89.735 -105.505 90.075 ;
        RECT -105.325 89.835 -104.775 90.005 ;
        RECT -100.725 89.835 -100.175 90.005 ;
        RECT -105.325 89.510 -105.155 89.835 ;
        RECT -106.225 89.340 -105.155 89.510 ;
        RECT -100.345 89.510 -100.175 89.835 ;
        RECT -99.995 89.735 -99.625 90.075 ;
        RECT -99.445 89.835 -98.515 90.015 ;
        RECT -97.065 89.835 -96.135 90.015 ;
        RECT -99.445 89.510 -99.275 89.835 ;
        RECT -100.345 89.340 -99.275 89.510 ;
        RECT -96.305 89.510 -96.135 89.835 ;
        RECT -95.955 89.735 -95.585 90.075 ;
        RECT -95.405 89.835 -94.855 90.005 ;
        RECT -90.805 89.835 -90.255 90.005 ;
        RECT -95.405 89.510 -95.235 89.835 ;
        RECT -96.305 89.340 -95.235 89.510 ;
        RECT -90.425 89.510 -90.255 89.835 ;
        RECT -90.075 89.735 -89.705 90.075 ;
        RECT -89.525 89.835 -88.595 90.015 ;
        RECT -87.145 89.835 -86.215 90.015 ;
        RECT -89.525 89.510 -89.355 89.835 ;
        RECT -90.425 89.340 -89.355 89.510 ;
        RECT -86.385 89.510 -86.215 89.835 ;
        RECT -86.035 89.735 -85.665 90.075 ;
        RECT -85.485 89.835 -84.935 90.005 ;
        RECT -80.885 89.835 -80.335 90.005 ;
        RECT -85.485 89.510 -85.315 89.835 ;
        RECT -86.385 89.340 -85.315 89.510 ;
        RECT -80.505 89.510 -80.335 89.835 ;
        RECT -80.155 89.735 -79.785 90.075 ;
        RECT -79.605 89.835 -78.675 90.015 ;
        RECT -77.225 89.835 -76.295 90.015 ;
        RECT -79.605 89.510 -79.435 89.835 ;
        RECT -80.505 89.340 -79.435 89.510 ;
        RECT -76.465 89.510 -76.295 89.835 ;
        RECT -76.115 89.735 -75.745 90.075 ;
        RECT -75.565 89.835 -75.015 90.005 ;
        RECT -70.965 89.835 -70.415 90.005 ;
        RECT -75.565 89.510 -75.395 89.835 ;
        RECT -76.465 89.340 -75.395 89.510 ;
        RECT -70.585 89.510 -70.415 89.835 ;
        RECT -70.235 89.735 -69.865 90.075 ;
        RECT -69.685 89.835 -68.755 90.015 ;
        RECT -67.305 89.835 -66.375 90.015 ;
        RECT -69.685 89.510 -69.515 89.835 ;
        RECT -70.585 89.340 -69.515 89.510 ;
        RECT -66.545 89.510 -66.375 89.835 ;
        RECT -66.195 89.735 -65.825 90.075 ;
        RECT -65.645 89.835 -65.095 90.005 ;
        RECT -61.045 89.835 -60.495 90.005 ;
        RECT -65.645 89.510 -65.475 89.835 ;
        RECT -66.545 89.340 -65.475 89.510 ;
        RECT -60.665 89.510 -60.495 89.835 ;
        RECT -60.315 89.735 -59.945 90.075 ;
        RECT -59.765 89.835 -58.835 90.015 ;
        RECT -57.385 89.835 -56.455 90.015 ;
        RECT -59.765 89.510 -59.595 89.835 ;
        RECT -60.665 89.340 -59.595 89.510 ;
        RECT -56.625 89.510 -56.455 89.835 ;
        RECT -56.275 89.735 -55.905 90.075 ;
        RECT -55.725 89.835 -55.175 90.005 ;
        RECT -51.125 89.835 -50.575 90.005 ;
        RECT -55.725 89.510 -55.555 89.835 ;
        RECT -56.625 89.340 -55.555 89.510 ;
        RECT -50.745 89.510 -50.575 89.835 ;
        RECT -50.395 89.735 -50.025 90.075 ;
        RECT -49.845 89.835 -48.915 90.015 ;
        RECT -47.465 89.835 -46.535 90.015 ;
        RECT -49.845 89.510 -49.675 89.835 ;
        RECT -50.745 89.340 -49.675 89.510 ;
        RECT -46.705 89.510 -46.535 89.835 ;
        RECT -46.355 89.735 -45.985 90.075 ;
        RECT -45.805 89.835 -45.255 90.005 ;
        RECT -41.205 89.835 -40.655 90.005 ;
        RECT -45.805 89.510 -45.635 89.835 ;
        RECT -46.705 89.340 -45.635 89.510 ;
        RECT -40.825 89.510 -40.655 89.835 ;
        RECT -40.475 89.735 -40.105 90.075 ;
        RECT -39.925 89.835 -38.995 90.015 ;
        RECT -37.545 89.835 -36.615 90.015 ;
        RECT -39.925 89.510 -39.755 89.835 ;
        RECT -40.825 89.340 -39.755 89.510 ;
        RECT -36.785 89.510 -36.615 89.835 ;
        RECT -36.435 89.735 -36.065 90.075 ;
        RECT -35.885 89.835 -35.335 90.005 ;
        RECT -31.285 89.835 -30.735 90.005 ;
        RECT -35.885 89.510 -35.715 89.835 ;
        RECT -36.785 89.340 -35.715 89.510 ;
        RECT -30.905 89.510 -30.735 89.835 ;
        RECT -30.555 89.735 -30.185 90.075 ;
        RECT -30.005 89.835 -29.075 90.015 ;
        RECT -27.625 89.835 -26.695 90.015 ;
        RECT -30.005 89.510 -29.835 89.835 ;
        RECT -30.905 89.340 -29.835 89.510 ;
        RECT -26.865 89.510 -26.695 89.835 ;
        RECT -26.515 89.735 -26.145 90.075 ;
        RECT -25.965 89.835 -25.415 90.005 ;
        RECT -21.365 89.835 -20.815 90.005 ;
        RECT -25.965 89.510 -25.795 89.835 ;
        RECT -26.865 89.340 -25.795 89.510 ;
        RECT -20.985 89.510 -20.815 89.835 ;
        RECT -20.635 89.735 -20.265 90.075 ;
        RECT -20.085 89.835 -19.155 90.015 ;
        RECT -17.705 89.835 -16.775 90.015 ;
        RECT -20.085 89.510 -19.915 89.835 ;
        RECT -20.985 89.340 -19.915 89.510 ;
        RECT -16.945 89.510 -16.775 89.835 ;
        RECT -16.595 89.735 -16.225 90.075 ;
        RECT -16.045 89.835 -15.495 90.005 ;
        RECT -11.445 89.835 -10.895 90.005 ;
        RECT -16.045 89.510 -15.875 89.835 ;
        RECT -16.945 89.340 -15.875 89.510 ;
        RECT -11.065 89.510 -10.895 89.835 ;
        RECT -10.715 89.735 -10.345 90.075 ;
        RECT -10.165 89.835 -9.235 90.015 ;
        RECT -7.785 89.835 -6.855 90.015 ;
        RECT -10.165 89.510 -9.995 89.835 ;
        RECT -11.065 89.340 -9.995 89.510 ;
        RECT -7.025 89.510 -6.855 89.835 ;
        RECT -6.675 89.735 -6.305 90.075 ;
        RECT -6.125 89.835 -5.575 90.005 ;
        RECT -1.525 89.835 -0.975 90.005 ;
        RECT -6.125 89.510 -5.955 89.835 ;
        RECT -7.025 89.340 -5.955 89.510 ;
        RECT -1.145 89.510 -0.975 89.835 ;
        RECT -0.795 89.735 -0.425 90.075 ;
        RECT -0.245 89.835 0.685 90.015 ;
        RECT 2.135 89.835 3.065 90.015 ;
        RECT -0.245 89.510 -0.075 89.835 ;
        RECT -1.145 89.340 -0.075 89.510 ;
        RECT 2.895 89.510 3.065 89.835 ;
        RECT 3.245 89.735 3.615 90.075 ;
        RECT 3.795 89.835 4.345 90.005 ;
        RECT 8.395 89.835 8.945 90.005 ;
        RECT 3.795 89.510 3.965 89.835 ;
        RECT 2.895 89.340 3.965 89.510 ;
        RECT 8.775 89.510 8.945 89.835 ;
        RECT 9.125 89.735 9.495 90.075 ;
        RECT 9.675 89.835 10.605 90.015 ;
        RECT 12.055 89.835 12.985 90.015 ;
        RECT 9.675 89.510 9.845 89.835 ;
        RECT 8.775 89.340 9.845 89.510 ;
        RECT 12.815 89.510 12.985 89.835 ;
        RECT 13.165 89.735 13.535 90.075 ;
        RECT 13.715 89.835 14.265 90.005 ;
        RECT 18.315 89.835 18.865 90.005 ;
        RECT 13.715 89.510 13.885 89.835 ;
        RECT 12.815 89.340 13.885 89.510 ;
        RECT 18.695 89.510 18.865 89.835 ;
        RECT 19.045 89.735 19.415 90.075 ;
        RECT 19.595 89.835 20.525 90.015 ;
        RECT 21.975 89.835 22.905 90.015 ;
        RECT 19.595 89.510 19.765 89.835 ;
        RECT 18.695 89.340 19.765 89.510 ;
        RECT 22.735 89.510 22.905 89.835 ;
        RECT 23.085 89.735 23.455 90.075 ;
        RECT 23.635 89.835 24.185 90.005 ;
        RECT 23.635 89.510 23.805 89.835 ;
        RECT 24.355 89.655 24.525 90.180 ;
        RECT 22.735 89.340 23.805 89.510 ;
        RECT -289.545 89.140 -289.375 89.325 ;
        RECT -288.400 89.235 -288.070 89.340 ;
        RECT -284.470 89.235 -284.140 89.340 ;
        RECT -278.480 89.235 -278.150 89.340 ;
        RECT -274.550 89.235 -274.220 89.340 ;
        RECT -268.560 89.235 -268.230 89.340 ;
        RECT -264.630 89.235 -264.300 89.340 ;
        RECT -258.640 89.235 -258.310 89.340 ;
        RECT -254.710 89.235 -254.380 89.340 ;
        RECT -248.720 89.235 -248.390 89.340 ;
        RECT -244.790 89.235 -244.460 89.340 ;
        RECT -238.800 89.235 -238.470 89.340 ;
        RECT -234.870 89.235 -234.540 89.340 ;
        RECT -228.880 89.235 -228.550 89.340 ;
        RECT -224.950 89.235 -224.620 89.340 ;
        RECT -218.960 89.235 -218.630 89.340 ;
        RECT -215.030 89.235 -214.700 89.340 ;
        RECT -209.040 89.235 -208.710 89.340 ;
        RECT -205.110 89.235 -204.780 89.340 ;
        RECT -199.120 89.235 -198.790 89.340 ;
        RECT -195.190 89.235 -194.860 89.340 ;
        RECT -189.200 89.235 -188.870 89.340 ;
        RECT -185.270 89.235 -184.940 89.340 ;
        RECT -179.280 89.235 -178.950 89.340 ;
        RECT -175.350 89.235 -175.020 89.340 ;
        RECT -169.360 89.235 -169.030 89.340 ;
        RECT -165.430 89.235 -165.100 89.340 ;
        RECT -159.440 89.235 -159.110 89.340 ;
        RECT -155.510 89.235 -155.180 89.340 ;
        RECT -149.520 89.235 -149.190 89.340 ;
        RECT -145.590 89.235 -145.260 89.340 ;
        RECT -139.600 89.235 -139.270 89.340 ;
        RECT -135.670 89.235 -135.340 89.340 ;
        RECT -129.680 89.235 -129.350 89.340 ;
        RECT -125.750 89.235 -125.420 89.340 ;
        RECT -119.760 89.235 -119.430 89.340 ;
        RECT -115.830 89.235 -115.500 89.340 ;
        RECT -109.840 89.235 -109.510 89.340 ;
        RECT -105.910 89.235 -105.580 89.340 ;
        RECT -99.920 89.235 -99.590 89.340 ;
        RECT -95.990 89.235 -95.660 89.340 ;
        RECT -90.000 89.235 -89.670 89.340 ;
        RECT -86.070 89.235 -85.740 89.340 ;
        RECT -80.080 89.235 -79.750 89.340 ;
        RECT -76.150 89.235 -75.820 89.340 ;
        RECT -70.160 89.235 -69.830 89.340 ;
        RECT -66.230 89.235 -65.900 89.340 ;
        RECT -60.240 89.235 -59.910 89.340 ;
        RECT -56.310 89.235 -55.980 89.340 ;
        RECT -50.320 89.235 -49.990 89.340 ;
        RECT -46.390 89.235 -46.060 89.340 ;
        RECT -40.400 89.235 -40.070 89.340 ;
        RECT -36.470 89.235 -36.140 89.340 ;
        RECT -30.480 89.235 -30.150 89.340 ;
        RECT -26.550 89.235 -26.220 89.340 ;
        RECT -20.560 89.235 -20.230 89.340 ;
        RECT -16.630 89.235 -16.300 89.340 ;
        RECT -10.640 89.235 -10.310 89.340 ;
        RECT -6.710 89.235 -6.380 89.340 ;
        RECT -0.720 89.235 -0.390 89.340 ;
        RECT 3.210 89.235 3.540 89.340 ;
        RECT 9.200 89.235 9.530 89.340 ;
        RECT 13.130 89.235 13.460 89.340 ;
        RECT 19.120 89.235 19.450 89.340 ;
        RECT 23.050 89.235 23.380 89.340 ;
        RECT 23.975 89.325 24.525 89.655 ;
        RECT -290.075 89.125 -289.375 89.140 ;
        RECT -290.160 88.955 -289.375 89.125 ;
        RECT -289.840 88.950 -289.375 88.955 ;
        RECT -289.545 88.800 -289.375 88.950 ;
        RECT -285.545 89.065 -284.640 89.155 ;
        RECT -283.840 89.065 -283.335 89.145 ;
        RECT -285.545 88.885 -283.335 89.065 ;
        RECT -275.625 89.065 -274.720 89.155 ;
        RECT -273.920 89.065 -273.415 89.145 ;
        RECT -275.625 88.885 -273.415 89.065 ;
        RECT -265.705 89.065 -264.800 89.155 ;
        RECT -264.000 89.065 -263.495 89.145 ;
        RECT -265.705 88.885 -263.495 89.065 ;
        RECT -255.785 89.065 -254.880 89.155 ;
        RECT -254.080 89.065 -253.575 89.145 ;
        RECT -255.785 88.885 -253.575 89.065 ;
        RECT -245.865 89.065 -244.960 89.155 ;
        RECT -244.160 89.065 -243.655 89.145 ;
        RECT -245.865 88.885 -243.655 89.065 ;
        RECT -235.945 89.065 -235.040 89.155 ;
        RECT -234.240 89.065 -233.735 89.145 ;
        RECT -235.945 88.885 -233.735 89.065 ;
        RECT -226.025 89.065 -225.120 89.155 ;
        RECT -224.320 89.065 -223.815 89.145 ;
        RECT -226.025 88.885 -223.815 89.065 ;
        RECT -216.105 89.065 -215.200 89.155 ;
        RECT -214.400 89.065 -213.895 89.145 ;
        RECT -216.105 88.885 -213.895 89.065 ;
        RECT -206.185 89.065 -205.280 89.155 ;
        RECT -204.480 89.065 -203.975 89.145 ;
        RECT -206.185 88.885 -203.975 89.065 ;
        RECT -196.265 89.065 -195.360 89.155 ;
        RECT -194.560 89.065 -194.055 89.145 ;
        RECT -196.265 88.885 -194.055 89.065 ;
        RECT -186.345 89.065 -185.440 89.155 ;
        RECT -184.640 89.065 -184.135 89.145 ;
        RECT -186.345 88.885 -184.135 89.065 ;
        RECT -176.425 89.065 -175.520 89.155 ;
        RECT -174.720 89.065 -174.215 89.145 ;
        RECT -176.425 88.885 -174.215 89.065 ;
        RECT -166.505 89.065 -165.600 89.155 ;
        RECT -164.800 89.065 -164.295 89.145 ;
        RECT -166.505 88.885 -164.295 89.065 ;
        RECT -156.585 89.065 -155.680 89.155 ;
        RECT -154.880 89.065 -154.375 89.145 ;
        RECT -156.585 88.885 -154.375 89.065 ;
        RECT -146.665 89.065 -145.760 89.155 ;
        RECT -144.960 89.065 -144.455 89.145 ;
        RECT -146.665 88.885 -144.455 89.065 ;
        RECT -136.745 89.065 -135.840 89.155 ;
        RECT -135.040 89.065 -134.535 89.145 ;
        RECT -136.745 88.885 -134.535 89.065 ;
        RECT -126.825 89.065 -125.920 89.155 ;
        RECT -125.120 89.065 -124.615 89.145 ;
        RECT -126.825 88.885 -124.615 89.065 ;
        RECT -116.905 89.065 -116.000 89.155 ;
        RECT -115.200 89.065 -114.695 89.145 ;
        RECT -116.905 88.885 -114.695 89.065 ;
        RECT -106.985 89.065 -106.080 89.155 ;
        RECT -105.280 89.065 -104.775 89.145 ;
        RECT -106.985 88.885 -104.775 89.065 ;
        RECT -97.065 89.065 -96.160 89.155 ;
        RECT -95.360 89.065 -94.855 89.145 ;
        RECT -97.065 88.885 -94.855 89.065 ;
        RECT -87.145 89.065 -86.240 89.155 ;
        RECT -85.440 89.065 -84.935 89.145 ;
        RECT -87.145 88.885 -84.935 89.065 ;
        RECT -77.225 89.065 -76.320 89.155 ;
        RECT -75.520 89.065 -75.015 89.145 ;
        RECT -77.225 88.885 -75.015 89.065 ;
        RECT -67.305 89.065 -66.400 89.155 ;
        RECT -65.600 89.065 -65.095 89.145 ;
        RECT -67.305 88.885 -65.095 89.065 ;
        RECT -57.385 89.065 -56.480 89.155 ;
        RECT -55.680 89.065 -55.175 89.145 ;
        RECT -57.385 88.885 -55.175 89.065 ;
        RECT -47.465 89.065 -46.560 89.155 ;
        RECT -45.760 89.065 -45.255 89.145 ;
        RECT -47.465 88.885 -45.255 89.065 ;
        RECT -37.545 89.065 -36.640 89.155 ;
        RECT -35.840 89.065 -35.335 89.145 ;
        RECT -37.545 88.885 -35.335 89.065 ;
        RECT -27.625 89.065 -26.720 89.155 ;
        RECT -25.920 89.065 -25.415 89.145 ;
        RECT -27.625 88.885 -25.415 89.065 ;
        RECT -17.705 89.065 -16.800 89.155 ;
        RECT -16.000 89.065 -15.495 89.145 ;
        RECT -17.705 88.885 -15.495 89.065 ;
        RECT -7.785 89.065 -6.880 89.155 ;
        RECT -6.080 89.065 -5.575 89.145 ;
        RECT -7.785 88.885 -5.575 89.065 ;
        RECT 2.135 89.065 3.040 89.155 ;
        RECT 3.840 89.065 4.345 89.145 ;
        RECT 2.135 88.885 4.345 89.065 ;
        RECT 12.055 89.065 12.960 89.155 ;
        RECT 13.760 89.065 14.265 89.145 ;
        RECT 12.055 88.885 14.265 89.065 ;
        RECT 21.975 89.065 22.880 89.155 ;
        RECT 23.680 89.065 24.185 89.145 ;
        RECT 21.975 88.885 24.185 89.065 ;
        RECT 24.355 89.130 24.525 89.325 ;
        RECT 24.765 89.130 25.055 89.850 ;
        RECT 24.355 89.125 25.055 89.130 ;
        RECT 24.355 88.955 25.140 89.125 ;
        RECT 24.355 88.950 24.820 88.955 ;
        RECT 24.355 88.800 24.525 88.950 ;
      LAYER mcon ;
        RECT -291.315 94.820 -291.145 94.990 ;
        RECT -290.845 94.825 -290.675 94.995 ;
        RECT -290.020 94.795 -289.850 94.965 ;
        RECT -288.655 94.795 -288.485 94.965 ;
        RECT -280.100 94.795 -279.930 94.965 ;
        RECT -278.735 94.795 -278.565 94.965 ;
        RECT -270.180 94.795 -270.010 94.965 ;
        RECT -268.815 94.795 -268.645 94.965 ;
        RECT -260.260 94.795 -260.090 94.965 ;
        RECT -258.895 94.795 -258.725 94.965 ;
        RECT -250.340 94.795 -250.170 94.965 ;
        RECT -248.975 94.795 -248.805 94.965 ;
        RECT -240.420 94.795 -240.250 94.965 ;
        RECT -239.055 94.795 -238.885 94.965 ;
        RECT -230.500 94.795 -230.330 94.965 ;
        RECT -229.135 94.795 -228.965 94.965 ;
        RECT -220.580 94.795 -220.410 94.965 ;
        RECT -219.215 94.795 -219.045 94.965 ;
        RECT -210.660 94.795 -210.490 94.965 ;
        RECT -209.295 94.795 -209.125 94.965 ;
        RECT -200.740 94.795 -200.570 94.965 ;
        RECT -199.375 94.795 -199.205 94.965 ;
        RECT -190.820 94.795 -190.650 94.965 ;
        RECT -189.455 94.795 -189.285 94.965 ;
        RECT -180.900 94.795 -180.730 94.965 ;
        RECT -179.535 94.795 -179.365 94.965 ;
        RECT -170.980 94.795 -170.810 94.965 ;
        RECT -169.615 94.795 -169.445 94.965 ;
        RECT -161.060 94.795 -160.890 94.965 ;
        RECT -159.695 94.795 -159.525 94.965 ;
        RECT -151.140 94.795 -150.970 94.965 ;
        RECT -149.775 94.795 -149.605 94.965 ;
        RECT -141.220 94.795 -141.050 94.965 ;
        RECT -139.855 94.795 -139.685 94.965 ;
        RECT -131.300 94.795 -131.130 94.965 ;
        RECT -129.935 94.795 -129.765 94.965 ;
        RECT -121.380 94.795 -121.210 94.965 ;
        RECT -120.015 94.795 -119.845 94.965 ;
        RECT -111.460 94.795 -111.290 94.965 ;
        RECT -110.095 94.795 -109.925 94.965 ;
        RECT -101.540 94.795 -101.370 94.965 ;
        RECT -100.175 94.795 -100.005 94.965 ;
        RECT -91.620 94.795 -91.450 94.965 ;
        RECT -90.255 94.795 -90.085 94.965 ;
        RECT -81.700 94.795 -81.530 94.965 ;
        RECT -80.335 94.795 -80.165 94.965 ;
        RECT -71.780 94.795 -71.610 94.965 ;
        RECT -70.415 94.795 -70.245 94.965 ;
        RECT -61.860 94.795 -61.690 94.965 ;
        RECT -60.495 94.795 -60.325 94.965 ;
        RECT -51.940 94.795 -51.770 94.965 ;
        RECT -50.575 94.795 -50.405 94.965 ;
        RECT -42.020 94.795 -41.850 94.965 ;
        RECT -40.655 94.795 -40.485 94.965 ;
        RECT -32.100 94.795 -31.930 94.965 ;
        RECT -30.735 94.795 -30.565 94.965 ;
        RECT -22.180 94.795 -22.010 94.965 ;
        RECT -20.815 94.795 -20.645 94.965 ;
        RECT -12.260 94.795 -12.090 94.965 ;
        RECT -10.895 94.795 -10.725 94.965 ;
        RECT -2.340 94.795 -2.170 94.965 ;
        RECT -0.975 94.795 -0.805 94.965 ;
        RECT 7.580 94.795 7.750 94.965 ;
        RECT 8.945 94.795 9.115 94.965 ;
        RECT 17.500 94.795 17.670 94.965 ;
        RECT 18.865 94.795 19.035 94.965 ;
        RECT -290.845 94.365 -290.675 94.535 ;
        RECT -290.845 93.905 -290.675 94.075 ;
        RECT -289.285 93.945 -289.115 94.115 ;
        RECT -283.425 93.945 -283.255 94.115 ;
        RECT -279.365 93.945 -279.195 94.115 ;
        RECT -273.505 93.945 -273.335 94.115 ;
        RECT -269.445 93.945 -269.275 94.115 ;
        RECT -263.585 93.945 -263.415 94.115 ;
        RECT -259.525 93.945 -259.355 94.115 ;
        RECT -253.665 93.945 -253.495 94.115 ;
        RECT -249.605 93.945 -249.435 94.115 ;
        RECT -243.745 93.945 -243.575 94.115 ;
        RECT -239.685 93.945 -239.515 94.115 ;
        RECT -233.825 93.945 -233.655 94.115 ;
        RECT -229.765 93.945 -229.595 94.115 ;
        RECT -223.905 93.945 -223.735 94.115 ;
        RECT -219.845 93.945 -219.675 94.115 ;
        RECT -213.985 93.945 -213.815 94.115 ;
        RECT -209.925 93.945 -209.755 94.115 ;
        RECT -204.065 93.945 -203.895 94.115 ;
        RECT -200.005 93.945 -199.835 94.115 ;
        RECT -194.145 93.945 -193.975 94.115 ;
        RECT -190.085 93.945 -189.915 94.115 ;
        RECT -184.225 93.945 -184.055 94.115 ;
        RECT -180.165 93.945 -179.995 94.115 ;
        RECT -174.305 93.945 -174.135 94.115 ;
        RECT -170.245 93.945 -170.075 94.115 ;
        RECT -164.385 93.945 -164.215 94.115 ;
        RECT -160.325 93.945 -160.155 94.115 ;
        RECT -154.465 93.945 -154.295 94.115 ;
        RECT -150.405 93.945 -150.235 94.115 ;
        RECT -144.545 93.945 -144.375 94.115 ;
        RECT -140.485 93.945 -140.315 94.115 ;
        RECT -134.625 93.945 -134.455 94.115 ;
        RECT -130.565 93.945 -130.395 94.115 ;
        RECT -124.705 93.945 -124.535 94.115 ;
        RECT -120.645 93.945 -120.475 94.115 ;
        RECT -114.785 93.945 -114.615 94.115 ;
        RECT -110.725 93.945 -110.555 94.115 ;
        RECT -104.865 93.945 -104.695 94.115 ;
        RECT -100.805 93.945 -100.635 94.115 ;
        RECT -94.945 93.945 -94.775 94.115 ;
        RECT -90.885 93.945 -90.715 94.115 ;
        RECT -85.025 93.945 -84.855 94.115 ;
        RECT -80.965 93.945 -80.795 94.115 ;
        RECT -75.105 93.945 -74.935 94.115 ;
        RECT -71.045 93.945 -70.875 94.115 ;
        RECT -65.185 93.945 -65.015 94.115 ;
        RECT -61.125 93.945 -60.955 94.115 ;
        RECT -55.265 93.945 -55.095 94.115 ;
        RECT -51.205 93.945 -51.035 94.115 ;
        RECT -45.345 93.945 -45.175 94.115 ;
        RECT -41.285 93.945 -41.115 94.115 ;
        RECT -35.425 93.945 -35.255 94.115 ;
        RECT -31.365 93.945 -31.195 94.115 ;
        RECT -25.505 93.945 -25.335 94.115 ;
        RECT -21.445 93.945 -21.275 94.115 ;
        RECT -15.585 93.945 -15.415 94.115 ;
        RECT -11.525 93.945 -11.355 94.115 ;
        RECT -5.665 93.945 -5.495 94.115 ;
        RECT -1.605 93.945 -1.435 94.115 ;
        RECT 4.255 93.945 4.425 94.115 ;
        RECT 8.315 93.945 8.485 94.115 ;
        RECT 14.175 93.945 14.345 94.115 ;
        RECT 18.235 93.945 18.405 94.115 ;
        RECT 24.095 93.945 24.265 94.115 ;
        RECT -291.315 93.245 -291.145 93.415 ;
        RECT -290.855 93.245 -290.685 93.415 ;
        RECT -290.395 93.245 -290.225 93.415 ;
        RECT -289.935 93.245 -289.765 93.415 ;
        RECT 24.745 93.245 24.915 93.415 ;
        RECT 25.205 93.245 25.375 93.415 ;
        RECT 25.665 93.245 25.835 93.415 ;
        RECT 26.125 93.245 26.295 93.415 ;
        RECT -289.965 92.525 -289.795 92.695 ;
        RECT -289.980 92.085 -289.810 92.255 ;
        RECT -282.745 92.525 -282.575 92.695 ;
        RECT -287.690 91.685 -287.520 91.855 ;
        RECT -287.705 91.245 -287.535 91.415 ;
        RECT -282.730 92.085 -282.560 92.255 ;
        RECT -285.020 91.685 -284.850 91.855 ;
        RECT -280.045 92.525 -279.875 92.695 ;
        RECT -280.060 92.085 -279.890 92.255 ;
        RECT -272.825 92.525 -272.655 92.695 ;
        RECT -285.005 91.245 -284.835 91.415 ;
        RECT -277.770 91.685 -277.600 91.855 ;
        RECT -277.785 91.245 -277.615 91.415 ;
        RECT -272.810 92.085 -272.640 92.255 ;
        RECT -275.100 91.685 -274.930 91.855 ;
        RECT -270.125 92.525 -269.955 92.695 ;
        RECT -270.140 92.085 -269.970 92.255 ;
        RECT -262.905 92.525 -262.735 92.695 ;
        RECT -275.085 91.245 -274.915 91.415 ;
        RECT -267.850 91.685 -267.680 91.855 ;
        RECT -267.865 91.245 -267.695 91.415 ;
        RECT -262.890 92.085 -262.720 92.255 ;
        RECT -265.180 91.685 -265.010 91.855 ;
        RECT -260.205 92.525 -260.035 92.695 ;
        RECT -260.220 92.085 -260.050 92.255 ;
        RECT -252.985 92.525 -252.815 92.695 ;
        RECT -265.165 91.245 -264.995 91.415 ;
        RECT -257.930 91.685 -257.760 91.855 ;
        RECT -257.945 91.245 -257.775 91.415 ;
        RECT -252.970 92.085 -252.800 92.255 ;
        RECT -255.260 91.685 -255.090 91.855 ;
        RECT -250.285 92.525 -250.115 92.695 ;
        RECT -250.300 92.085 -250.130 92.255 ;
        RECT -243.065 92.525 -242.895 92.695 ;
        RECT -255.245 91.245 -255.075 91.415 ;
        RECT -248.010 91.685 -247.840 91.855 ;
        RECT -248.025 91.245 -247.855 91.415 ;
        RECT -243.050 92.085 -242.880 92.255 ;
        RECT -245.340 91.685 -245.170 91.855 ;
        RECT -240.365 92.525 -240.195 92.695 ;
        RECT -240.380 92.085 -240.210 92.255 ;
        RECT -233.145 92.525 -232.975 92.695 ;
        RECT -245.325 91.245 -245.155 91.415 ;
        RECT -238.090 91.685 -237.920 91.855 ;
        RECT -238.105 91.245 -237.935 91.415 ;
        RECT -233.130 92.085 -232.960 92.255 ;
        RECT -235.420 91.685 -235.250 91.855 ;
        RECT -230.445 92.525 -230.275 92.695 ;
        RECT -230.460 92.085 -230.290 92.255 ;
        RECT -223.225 92.525 -223.055 92.695 ;
        RECT -235.405 91.245 -235.235 91.415 ;
        RECT -228.170 91.685 -228.000 91.855 ;
        RECT -228.185 91.245 -228.015 91.415 ;
        RECT -223.210 92.085 -223.040 92.255 ;
        RECT -225.500 91.685 -225.330 91.855 ;
        RECT -220.525 92.525 -220.355 92.695 ;
        RECT -220.540 92.085 -220.370 92.255 ;
        RECT -213.305 92.525 -213.135 92.695 ;
        RECT -225.485 91.245 -225.315 91.415 ;
        RECT -218.250 91.685 -218.080 91.855 ;
        RECT -218.265 91.245 -218.095 91.415 ;
        RECT -213.290 92.085 -213.120 92.255 ;
        RECT -215.580 91.685 -215.410 91.855 ;
        RECT -210.605 92.525 -210.435 92.695 ;
        RECT -210.620 92.085 -210.450 92.255 ;
        RECT -203.385 92.525 -203.215 92.695 ;
        RECT -215.565 91.245 -215.395 91.415 ;
        RECT -208.330 91.685 -208.160 91.855 ;
        RECT -208.345 91.245 -208.175 91.415 ;
        RECT -203.370 92.085 -203.200 92.255 ;
        RECT -205.660 91.685 -205.490 91.855 ;
        RECT -200.685 92.525 -200.515 92.695 ;
        RECT -200.700 92.085 -200.530 92.255 ;
        RECT -193.465 92.525 -193.295 92.695 ;
        RECT -205.645 91.245 -205.475 91.415 ;
        RECT -198.410 91.685 -198.240 91.855 ;
        RECT -198.425 91.245 -198.255 91.415 ;
        RECT -193.450 92.085 -193.280 92.255 ;
        RECT -195.740 91.685 -195.570 91.855 ;
        RECT -190.765 92.525 -190.595 92.695 ;
        RECT -190.780 92.085 -190.610 92.255 ;
        RECT -183.545 92.525 -183.375 92.695 ;
        RECT -195.725 91.245 -195.555 91.415 ;
        RECT -188.490 91.685 -188.320 91.855 ;
        RECT -188.505 91.245 -188.335 91.415 ;
        RECT -183.530 92.085 -183.360 92.255 ;
        RECT -185.820 91.685 -185.650 91.855 ;
        RECT -180.845 92.525 -180.675 92.695 ;
        RECT -180.860 92.085 -180.690 92.255 ;
        RECT -173.625 92.525 -173.455 92.695 ;
        RECT -185.805 91.245 -185.635 91.415 ;
        RECT -178.570 91.685 -178.400 91.855 ;
        RECT -178.585 91.245 -178.415 91.415 ;
        RECT -173.610 92.085 -173.440 92.255 ;
        RECT -175.900 91.685 -175.730 91.855 ;
        RECT -170.925 92.525 -170.755 92.695 ;
        RECT -170.940 92.085 -170.770 92.255 ;
        RECT -163.705 92.525 -163.535 92.695 ;
        RECT -175.885 91.245 -175.715 91.415 ;
        RECT -168.650 91.685 -168.480 91.855 ;
        RECT -168.665 91.245 -168.495 91.415 ;
        RECT -163.690 92.085 -163.520 92.255 ;
        RECT -165.980 91.685 -165.810 91.855 ;
        RECT -161.005 92.525 -160.835 92.695 ;
        RECT -161.020 92.085 -160.850 92.255 ;
        RECT -153.785 92.525 -153.615 92.695 ;
        RECT -165.965 91.245 -165.795 91.415 ;
        RECT -158.730 91.685 -158.560 91.855 ;
        RECT -158.745 91.245 -158.575 91.415 ;
        RECT -153.770 92.085 -153.600 92.255 ;
        RECT -156.060 91.685 -155.890 91.855 ;
        RECT -151.085 92.525 -150.915 92.695 ;
        RECT -151.100 92.085 -150.930 92.255 ;
        RECT -143.865 92.525 -143.695 92.695 ;
        RECT -156.045 91.245 -155.875 91.415 ;
        RECT -148.810 91.685 -148.640 91.855 ;
        RECT -148.825 91.245 -148.655 91.415 ;
        RECT -143.850 92.085 -143.680 92.255 ;
        RECT -146.140 91.685 -145.970 91.855 ;
        RECT -141.165 92.525 -140.995 92.695 ;
        RECT -141.180 92.085 -141.010 92.255 ;
        RECT -133.945 92.525 -133.775 92.695 ;
        RECT -146.125 91.245 -145.955 91.415 ;
        RECT -138.890 91.685 -138.720 91.855 ;
        RECT -138.905 91.245 -138.735 91.415 ;
        RECT -133.930 92.085 -133.760 92.255 ;
        RECT -136.220 91.685 -136.050 91.855 ;
        RECT -131.245 92.525 -131.075 92.695 ;
        RECT -131.260 92.085 -131.090 92.255 ;
        RECT -124.025 92.525 -123.855 92.695 ;
        RECT -136.205 91.245 -136.035 91.415 ;
        RECT -128.970 91.685 -128.800 91.855 ;
        RECT -128.985 91.245 -128.815 91.415 ;
        RECT -124.010 92.085 -123.840 92.255 ;
        RECT -126.300 91.685 -126.130 91.855 ;
        RECT -121.325 92.525 -121.155 92.695 ;
        RECT -121.340 92.085 -121.170 92.255 ;
        RECT -114.105 92.525 -113.935 92.695 ;
        RECT -126.285 91.245 -126.115 91.415 ;
        RECT -119.050 91.685 -118.880 91.855 ;
        RECT -119.065 91.245 -118.895 91.415 ;
        RECT -114.090 92.085 -113.920 92.255 ;
        RECT -116.380 91.685 -116.210 91.855 ;
        RECT -111.405 92.525 -111.235 92.695 ;
        RECT -111.420 92.085 -111.250 92.255 ;
        RECT -104.185 92.525 -104.015 92.695 ;
        RECT -116.365 91.245 -116.195 91.415 ;
        RECT -109.130 91.685 -108.960 91.855 ;
        RECT -109.145 91.245 -108.975 91.415 ;
        RECT -104.170 92.085 -104.000 92.255 ;
        RECT -106.460 91.685 -106.290 91.855 ;
        RECT -101.485 92.525 -101.315 92.695 ;
        RECT -101.500 92.085 -101.330 92.255 ;
        RECT -94.265 92.525 -94.095 92.695 ;
        RECT -106.445 91.245 -106.275 91.415 ;
        RECT -99.210 91.685 -99.040 91.855 ;
        RECT -99.225 91.245 -99.055 91.415 ;
        RECT -94.250 92.085 -94.080 92.255 ;
        RECT -96.540 91.685 -96.370 91.855 ;
        RECT -91.565 92.525 -91.395 92.695 ;
        RECT -91.580 92.085 -91.410 92.255 ;
        RECT -84.345 92.525 -84.175 92.695 ;
        RECT -96.525 91.245 -96.355 91.415 ;
        RECT -89.290 91.685 -89.120 91.855 ;
        RECT -89.305 91.245 -89.135 91.415 ;
        RECT -84.330 92.085 -84.160 92.255 ;
        RECT -86.620 91.685 -86.450 91.855 ;
        RECT -81.645 92.525 -81.475 92.695 ;
        RECT -81.660 92.085 -81.490 92.255 ;
        RECT -74.425 92.525 -74.255 92.695 ;
        RECT -86.605 91.245 -86.435 91.415 ;
        RECT -79.370 91.685 -79.200 91.855 ;
        RECT -79.385 91.245 -79.215 91.415 ;
        RECT -74.410 92.085 -74.240 92.255 ;
        RECT -76.700 91.685 -76.530 91.855 ;
        RECT -71.725 92.525 -71.555 92.695 ;
        RECT -71.740 92.085 -71.570 92.255 ;
        RECT -64.505 92.525 -64.335 92.695 ;
        RECT -76.685 91.245 -76.515 91.415 ;
        RECT -69.450 91.685 -69.280 91.855 ;
        RECT -69.465 91.245 -69.295 91.415 ;
        RECT -64.490 92.085 -64.320 92.255 ;
        RECT -66.780 91.685 -66.610 91.855 ;
        RECT -61.805 92.525 -61.635 92.695 ;
        RECT -61.820 92.085 -61.650 92.255 ;
        RECT -54.585 92.525 -54.415 92.695 ;
        RECT -66.765 91.245 -66.595 91.415 ;
        RECT -59.530 91.685 -59.360 91.855 ;
        RECT -59.545 91.245 -59.375 91.415 ;
        RECT -54.570 92.085 -54.400 92.255 ;
        RECT -56.860 91.685 -56.690 91.855 ;
        RECT -51.885 92.525 -51.715 92.695 ;
        RECT -51.900 92.085 -51.730 92.255 ;
        RECT -44.665 92.525 -44.495 92.695 ;
        RECT -56.845 91.245 -56.675 91.415 ;
        RECT -49.610 91.685 -49.440 91.855 ;
        RECT -49.625 91.245 -49.455 91.415 ;
        RECT -44.650 92.085 -44.480 92.255 ;
        RECT -46.940 91.685 -46.770 91.855 ;
        RECT -41.965 92.525 -41.795 92.695 ;
        RECT -41.980 92.085 -41.810 92.255 ;
        RECT -34.745 92.525 -34.575 92.695 ;
        RECT -46.925 91.245 -46.755 91.415 ;
        RECT -39.690 91.685 -39.520 91.855 ;
        RECT -39.705 91.245 -39.535 91.415 ;
        RECT -34.730 92.085 -34.560 92.255 ;
        RECT -37.020 91.685 -36.850 91.855 ;
        RECT -32.045 92.525 -31.875 92.695 ;
        RECT -32.060 92.085 -31.890 92.255 ;
        RECT -24.825 92.525 -24.655 92.695 ;
        RECT -37.005 91.245 -36.835 91.415 ;
        RECT -29.770 91.685 -29.600 91.855 ;
        RECT -29.785 91.245 -29.615 91.415 ;
        RECT -24.810 92.085 -24.640 92.255 ;
        RECT -27.100 91.685 -26.930 91.855 ;
        RECT -22.125 92.525 -21.955 92.695 ;
        RECT -22.140 92.085 -21.970 92.255 ;
        RECT -14.905 92.525 -14.735 92.695 ;
        RECT -27.085 91.245 -26.915 91.415 ;
        RECT -19.850 91.685 -19.680 91.855 ;
        RECT -19.865 91.245 -19.695 91.415 ;
        RECT -14.890 92.085 -14.720 92.255 ;
        RECT -17.180 91.685 -17.010 91.855 ;
        RECT -12.205 92.525 -12.035 92.695 ;
        RECT -12.220 92.085 -12.050 92.255 ;
        RECT -4.985 92.525 -4.815 92.695 ;
        RECT -17.165 91.245 -16.995 91.415 ;
        RECT -9.930 91.685 -9.760 91.855 ;
        RECT -9.945 91.245 -9.775 91.415 ;
        RECT -4.970 92.085 -4.800 92.255 ;
        RECT -7.260 91.685 -7.090 91.855 ;
        RECT -2.285 92.525 -2.115 92.695 ;
        RECT -2.300 92.085 -2.130 92.255 ;
        RECT 4.935 92.525 5.105 92.695 ;
        RECT -7.245 91.245 -7.075 91.415 ;
        RECT -0.010 91.685 0.160 91.855 ;
        RECT -0.025 91.245 0.145 91.415 ;
        RECT 4.950 92.085 5.120 92.255 ;
        RECT 2.660 91.685 2.830 91.855 ;
        RECT 7.635 92.525 7.805 92.695 ;
        RECT 7.620 92.085 7.790 92.255 ;
        RECT 14.855 92.525 15.025 92.695 ;
        RECT 2.675 91.245 2.845 91.415 ;
        RECT 9.910 91.685 10.080 91.855 ;
        RECT 9.895 91.245 10.065 91.415 ;
        RECT 14.870 92.085 15.040 92.255 ;
        RECT 12.580 91.685 12.750 91.855 ;
        RECT 17.555 92.525 17.725 92.695 ;
        RECT 17.540 92.085 17.710 92.255 ;
        RECT 24.775 92.525 24.945 92.695 ;
        RECT 12.595 91.245 12.765 91.415 ;
        RECT 19.830 91.685 20.000 91.855 ;
        RECT 19.815 91.245 19.985 91.415 ;
        RECT 24.790 92.085 24.960 92.255 ;
        RECT 22.500 91.685 22.670 91.855 ;
        RECT 22.515 91.245 22.685 91.415 ;
        RECT -291.315 90.525 -291.145 90.695 ;
        RECT -290.855 90.525 -290.685 90.695 ;
        RECT -290.395 90.525 -290.225 90.695 ;
        RECT -289.935 90.525 -289.765 90.695 ;
        RECT -289.545 89.865 -289.375 90.035 ;
        RECT -289.545 89.405 -289.375 89.575 ;
        RECT -288.385 89.825 -288.215 89.995 ;
        RECT -284.325 89.825 -284.155 89.995 ;
        RECT -278.465 89.825 -278.295 89.995 ;
        RECT -274.405 89.825 -274.235 89.995 ;
        RECT -268.545 89.825 -268.375 89.995 ;
        RECT -264.485 89.825 -264.315 89.995 ;
        RECT -258.625 89.825 -258.455 89.995 ;
        RECT -254.565 89.825 -254.395 89.995 ;
        RECT -248.705 89.825 -248.535 89.995 ;
        RECT -244.645 89.825 -244.475 89.995 ;
        RECT -238.785 89.825 -238.615 89.995 ;
        RECT -234.725 89.825 -234.555 89.995 ;
        RECT -228.865 89.825 -228.695 89.995 ;
        RECT -224.805 89.825 -224.635 89.995 ;
        RECT -218.945 89.825 -218.775 89.995 ;
        RECT -214.885 89.825 -214.715 89.995 ;
        RECT -209.025 89.825 -208.855 89.995 ;
        RECT -204.965 89.825 -204.795 89.995 ;
        RECT -199.105 89.825 -198.935 89.995 ;
        RECT -195.045 89.825 -194.875 89.995 ;
        RECT -189.185 89.825 -189.015 89.995 ;
        RECT -185.125 89.825 -184.955 89.995 ;
        RECT -179.265 89.825 -179.095 89.995 ;
        RECT -175.205 89.825 -175.035 89.995 ;
        RECT -169.345 89.825 -169.175 89.995 ;
        RECT -165.285 89.825 -165.115 89.995 ;
        RECT -159.425 89.825 -159.255 89.995 ;
        RECT -155.365 89.825 -155.195 89.995 ;
        RECT -149.505 89.825 -149.335 89.995 ;
        RECT -145.445 89.825 -145.275 89.995 ;
        RECT -139.585 89.825 -139.415 89.995 ;
        RECT -135.525 89.825 -135.355 89.995 ;
        RECT -129.665 89.825 -129.495 89.995 ;
        RECT -125.605 89.825 -125.435 89.995 ;
        RECT -119.745 89.825 -119.575 89.995 ;
        RECT -115.685 89.825 -115.515 89.995 ;
        RECT -109.825 89.825 -109.655 89.995 ;
        RECT -105.765 89.825 -105.595 89.995 ;
        RECT -99.905 89.825 -99.735 89.995 ;
        RECT -95.845 89.825 -95.675 89.995 ;
        RECT -89.985 89.825 -89.815 89.995 ;
        RECT -85.925 89.825 -85.755 89.995 ;
        RECT -80.065 89.825 -79.895 89.995 ;
        RECT -76.005 89.825 -75.835 89.995 ;
        RECT -70.145 89.825 -69.975 89.995 ;
        RECT -66.085 89.825 -65.915 89.995 ;
        RECT -60.225 89.825 -60.055 89.995 ;
        RECT -56.165 89.825 -55.995 89.995 ;
        RECT -50.305 89.825 -50.135 89.995 ;
        RECT -46.245 89.825 -46.075 89.995 ;
        RECT -40.385 89.825 -40.215 89.995 ;
        RECT -36.325 89.825 -36.155 89.995 ;
        RECT -30.465 89.825 -30.295 89.995 ;
        RECT -26.405 89.825 -26.235 89.995 ;
        RECT -20.545 89.825 -20.375 89.995 ;
        RECT -16.485 89.825 -16.315 89.995 ;
        RECT -10.625 89.825 -10.455 89.995 ;
        RECT -6.565 89.825 -6.395 89.995 ;
        RECT -0.705 89.825 -0.535 89.995 ;
        RECT 3.355 89.825 3.525 89.995 ;
        RECT 9.215 89.825 9.385 89.995 ;
        RECT 13.275 89.825 13.445 89.995 ;
        RECT 19.135 89.825 19.305 89.995 ;
        RECT 23.195 89.825 23.365 89.995 ;
        RECT 24.355 89.865 24.525 90.035 ;
        RECT 24.355 89.405 24.525 89.575 ;
        RECT -290.015 88.955 -289.845 89.125 ;
        RECT -289.545 88.945 -289.375 89.115 ;
        RECT -285.060 88.975 -284.890 89.145 ;
        RECT -283.695 88.975 -283.525 89.145 ;
        RECT -275.140 88.975 -274.970 89.145 ;
        RECT -273.775 88.975 -273.605 89.145 ;
        RECT -265.220 88.975 -265.050 89.145 ;
        RECT -263.855 88.975 -263.685 89.145 ;
        RECT -255.300 88.975 -255.130 89.145 ;
        RECT -253.935 88.975 -253.765 89.145 ;
        RECT -245.380 88.975 -245.210 89.145 ;
        RECT -244.015 88.975 -243.845 89.145 ;
        RECT -235.460 88.975 -235.290 89.145 ;
        RECT -234.095 88.975 -233.925 89.145 ;
        RECT -225.540 88.975 -225.370 89.145 ;
        RECT -224.175 88.975 -224.005 89.145 ;
        RECT -215.620 88.975 -215.450 89.145 ;
        RECT -214.255 88.975 -214.085 89.145 ;
        RECT -205.700 88.975 -205.530 89.145 ;
        RECT -204.335 88.975 -204.165 89.145 ;
        RECT -195.780 88.975 -195.610 89.145 ;
        RECT -194.415 88.975 -194.245 89.145 ;
        RECT -185.860 88.975 -185.690 89.145 ;
        RECT -184.495 88.975 -184.325 89.145 ;
        RECT -175.940 88.975 -175.770 89.145 ;
        RECT -174.575 88.975 -174.405 89.145 ;
        RECT -166.020 88.975 -165.850 89.145 ;
        RECT -164.655 88.975 -164.485 89.145 ;
        RECT -156.100 88.975 -155.930 89.145 ;
        RECT -154.735 88.975 -154.565 89.145 ;
        RECT -146.180 88.975 -146.010 89.145 ;
        RECT -144.815 88.975 -144.645 89.145 ;
        RECT -136.260 88.975 -136.090 89.145 ;
        RECT -134.895 88.975 -134.725 89.145 ;
        RECT -126.340 88.975 -126.170 89.145 ;
        RECT -124.975 88.975 -124.805 89.145 ;
        RECT -116.420 88.975 -116.250 89.145 ;
        RECT -115.055 88.975 -114.885 89.145 ;
        RECT -106.500 88.975 -106.330 89.145 ;
        RECT -105.135 88.975 -104.965 89.145 ;
        RECT -96.580 88.975 -96.410 89.145 ;
        RECT -95.215 88.975 -95.045 89.145 ;
        RECT -86.660 88.975 -86.490 89.145 ;
        RECT -85.295 88.975 -85.125 89.145 ;
        RECT -76.740 88.975 -76.570 89.145 ;
        RECT -75.375 88.975 -75.205 89.145 ;
        RECT -66.820 88.975 -66.650 89.145 ;
        RECT -65.455 88.975 -65.285 89.145 ;
        RECT -56.900 88.975 -56.730 89.145 ;
        RECT -55.535 88.975 -55.365 89.145 ;
        RECT -46.980 88.975 -46.810 89.145 ;
        RECT -45.615 88.975 -45.445 89.145 ;
        RECT -37.060 88.975 -36.890 89.145 ;
        RECT -35.695 88.975 -35.525 89.145 ;
        RECT -27.140 88.975 -26.970 89.145 ;
        RECT -25.775 88.975 -25.605 89.145 ;
        RECT -17.220 88.975 -17.050 89.145 ;
        RECT -15.855 88.975 -15.685 89.145 ;
        RECT -7.300 88.975 -7.130 89.145 ;
        RECT -5.935 88.975 -5.765 89.145 ;
        RECT 2.620 88.975 2.790 89.145 ;
        RECT 3.985 88.975 4.155 89.145 ;
        RECT 12.540 88.975 12.710 89.145 ;
        RECT 13.905 88.975 14.075 89.145 ;
        RECT 22.460 88.975 22.630 89.145 ;
        RECT 23.825 88.975 23.995 89.145 ;
        RECT 24.355 88.945 24.525 89.115 ;
        RECT 24.825 88.955 24.995 89.125 ;
      LAYER met1 ;
        RECT -291.460 95.140 -291.000 95.145 ;
        RECT -291.460 94.665 -290.520 95.140 ;
        RECT -289.600 95.060 -288.600 95.760 ;
        RECT -279.680 95.060 -278.680 95.760 ;
        RECT -269.760 95.060 -268.760 95.760 ;
        RECT -259.840 95.060 -258.840 95.760 ;
        RECT -249.920 95.060 -248.920 95.760 ;
        RECT -240.000 95.060 -239.000 95.760 ;
        RECT -230.080 95.060 -229.080 95.760 ;
        RECT -220.160 95.060 -219.160 95.760 ;
        RECT -210.240 95.060 -209.240 95.760 ;
        RECT -200.320 95.060 -199.320 95.760 ;
        RECT -190.400 95.060 -189.400 95.760 ;
        RECT -180.480 95.060 -179.480 95.760 ;
        RECT -170.560 95.060 -169.560 95.760 ;
        RECT -160.640 95.060 -159.640 95.760 ;
        RECT -150.720 95.060 -149.720 95.760 ;
        RECT -140.800 95.060 -139.800 95.760 ;
        RECT -130.880 95.060 -129.880 95.760 ;
        RECT -120.960 95.060 -119.960 95.760 ;
        RECT -111.040 95.060 -110.040 95.760 ;
        RECT -101.120 95.060 -100.120 95.760 ;
        RECT -91.200 95.060 -90.200 95.760 ;
        RECT -81.280 95.060 -80.280 95.760 ;
        RECT -71.360 95.060 -70.360 95.760 ;
        RECT -61.440 95.060 -60.440 95.760 ;
        RECT -51.520 95.060 -50.520 95.760 ;
        RECT -41.600 95.060 -40.600 95.760 ;
        RECT -31.680 95.060 -30.680 95.760 ;
        RECT -21.760 95.060 -20.760 95.760 ;
        RECT -11.840 95.060 -10.840 95.760 ;
        RECT -1.920 95.060 -0.920 95.760 ;
        RECT 8.000 95.060 9.000 95.760 ;
        RECT 17.920 95.060 18.920 95.760 ;
        RECT -290.110 94.760 -288.420 95.060 ;
        RECT -280.190 94.760 -278.500 95.060 ;
        RECT -270.270 94.760 -268.580 95.060 ;
        RECT -260.350 94.760 -258.660 95.060 ;
        RECT -250.430 94.760 -248.740 95.060 ;
        RECT -240.510 94.760 -238.820 95.060 ;
        RECT -230.590 94.760 -228.900 95.060 ;
        RECT -220.670 94.760 -218.980 95.060 ;
        RECT -210.750 94.760 -209.060 95.060 ;
        RECT -200.830 94.760 -199.140 95.060 ;
        RECT -190.910 94.760 -189.220 95.060 ;
        RECT -180.990 94.760 -179.300 95.060 ;
        RECT -171.070 94.760 -169.380 95.060 ;
        RECT -161.150 94.760 -159.460 95.060 ;
        RECT -151.230 94.760 -149.540 95.060 ;
        RECT -141.310 94.760 -139.620 95.060 ;
        RECT -131.390 94.760 -129.700 95.060 ;
        RECT -121.470 94.760 -119.780 95.060 ;
        RECT -111.550 94.760 -109.860 95.060 ;
        RECT -101.630 94.760 -99.940 95.060 ;
        RECT -91.710 94.760 -90.020 95.060 ;
        RECT -81.790 94.760 -80.100 95.060 ;
        RECT -71.870 94.760 -70.180 95.060 ;
        RECT -61.950 94.760 -60.260 95.060 ;
        RECT -52.030 94.760 -50.340 95.060 ;
        RECT -42.110 94.760 -40.420 95.060 ;
        RECT -32.190 94.760 -30.500 95.060 ;
        RECT -22.270 94.760 -20.580 95.060 ;
        RECT -12.350 94.760 -10.660 95.060 ;
        RECT -2.430 94.760 -0.740 95.060 ;
        RECT 7.490 94.760 9.180 95.060 ;
        RECT 17.410 94.760 19.100 95.060 ;
        RECT -291.000 93.760 -290.520 94.665 ;
        RECT -289.370 93.890 -289.050 94.180 ;
        RECT -283.490 93.890 -283.170 94.180 ;
        RECT -279.450 93.890 -279.130 94.180 ;
        RECT -273.570 93.890 -273.250 94.180 ;
        RECT -269.530 93.890 -269.210 94.180 ;
        RECT -263.650 93.890 -263.330 94.180 ;
        RECT -259.610 93.890 -259.290 94.180 ;
        RECT -253.730 93.890 -253.410 94.180 ;
        RECT -249.690 93.890 -249.370 94.180 ;
        RECT -243.810 93.890 -243.490 94.180 ;
        RECT -239.770 93.890 -239.450 94.180 ;
        RECT -233.890 93.890 -233.570 94.180 ;
        RECT -229.850 93.890 -229.530 94.180 ;
        RECT -223.970 93.890 -223.650 94.180 ;
        RECT -219.930 93.890 -219.610 94.180 ;
        RECT -214.050 93.890 -213.730 94.180 ;
        RECT -210.010 93.890 -209.690 94.180 ;
        RECT -204.130 93.890 -203.810 94.180 ;
        RECT -200.090 93.890 -199.770 94.180 ;
        RECT -194.210 93.890 -193.890 94.180 ;
        RECT -190.170 93.890 -189.850 94.180 ;
        RECT -184.290 93.890 -183.970 94.180 ;
        RECT -180.250 93.890 -179.930 94.180 ;
        RECT -174.370 93.890 -174.050 94.180 ;
        RECT -170.330 93.890 -170.010 94.180 ;
        RECT -164.450 93.890 -164.130 94.180 ;
        RECT -160.410 93.890 -160.090 94.180 ;
        RECT -154.530 93.890 -154.210 94.180 ;
        RECT -150.490 93.890 -150.170 94.180 ;
        RECT -144.610 93.890 -144.290 94.180 ;
        RECT -140.570 93.890 -140.250 94.180 ;
        RECT -134.690 93.890 -134.370 94.180 ;
        RECT -130.650 93.890 -130.330 94.180 ;
        RECT -124.770 93.890 -124.450 94.180 ;
        RECT -120.730 93.890 -120.410 94.180 ;
        RECT -114.850 93.890 -114.530 94.180 ;
        RECT -110.810 93.890 -110.490 94.180 ;
        RECT -104.930 93.890 -104.610 94.180 ;
        RECT -100.890 93.890 -100.570 94.180 ;
        RECT -95.010 93.890 -94.690 94.180 ;
        RECT -90.970 93.890 -90.650 94.180 ;
        RECT -85.090 93.890 -84.770 94.180 ;
        RECT -81.050 93.890 -80.730 94.180 ;
        RECT -75.170 93.890 -74.850 94.180 ;
        RECT -71.130 93.890 -70.810 94.180 ;
        RECT -65.250 93.890 -64.930 94.180 ;
        RECT -61.210 93.890 -60.890 94.180 ;
        RECT -55.330 93.890 -55.010 94.180 ;
        RECT -51.290 93.890 -50.970 94.180 ;
        RECT -45.410 93.890 -45.090 94.180 ;
        RECT -41.370 93.890 -41.050 94.180 ;
        RECT -35.490 93.890 -35.170 94.180 ;
        RECT -31.450 93.890 -31.130 94.180 ;
        RECT -25.570 93.890 -25.250 94.180 ;
        RECT -21.530 93.890 -21.210 94.180 ;
        RECT -15.650 93.890 -15.330 94.180 ;
        RECT -11.610 93.890 -11.290 94.180 ;
        RECT -5.730 93.890 -5.410 94.180 ;
        RECT -1.690 93.890 -1.370 94.180 ;
        RECT 4.190 93.890 4.510 94.180 ;
        RECT 8.230 93.890 8.550 94.180 ;
        RECT 14.110 93.890 14.430 94.180 ;
        RECT 18.150 93.890 18.470 94.180 ;
        RECT 24.030 93.890 24.350 94.180 ;
        RECT -291.460 93.090 -289.620 93.570 ;
        RECT -289.290 92.760 -289.100 93.890 ;
        RECT -283.440 92.760 -283.250 93.890 ;
        RECT -279.370 92.760 -279.180 93.890 ;
        RECT -273.520 92.760 -273.330 93.890 ;
        RECT -269.450 92.760 -269.260 93.890 ;
        RECT -263.600 92.760 -263.410 93.890 ;
        RECT -259.530 92.760 -259.340 93.890 ;
        RECT -253.680 92.760 -253.490 93.890 ;
        RECT -249.610 92.760 -249.420 93.890 ;
        RECT -243.760 92.760 -243.570 93.890 ;
        RECT -239.690 92.760 -239.500 93.890 ;
        RECT -233.840 92.760 -233.650 93.890 ;
        RECT -229.770 92.760 -229.580 93.890 ;
        RECT -223.920 92.760 -223.730 93.890 ;
        RECT -219.850 92.760 -219.660 93.890 ;
        RECT -214.000 92.760 -213.810 93.890 ;
        RECT -209.930 92.760 -209.740 93.890 ;
        RECT -204.080 92.760 -203.890 93.890 ;
        RECT -200.010 92.760 -199.820 93.890 ;
        RECT -194.160 92.760 -193.970 93.890 ;
        RECT -190.090 92.760 -189.900 93.890 ;
        RECT -184.240 92.760 -184.050 93.890 ;
        RECT -180.170 92.760 -179.980 93.890 ;
        RECT -174.320 92.760 -174.130 93.890 ;
        RECT -170.250 92.760 -170.060 93.890 ;
        RECT -164.400 92.760 -164.210 93.890 ;
        RECT -160.330 92.760 -160.140 93.890 ;
        RECT -154.480 92.760 -154.290 93.890 ;
        RECT -150.410 92.760 -150.220 93.890 ;
        RECT -144.560 92.760 -144.370 93.890 ;
        RECT -140.490 92.760 -140.300 93.890 ;
        RECT -134.640 92.760 -134.450 93.890 ;
        RECT -130.570 92.760 -130.380 93.890 ;
        RECT -124.720 92.760 -124.530 93.890 ;
        RECT -120.650 92.760 -120.460 93.890 ;
        RECT -114.800 92.760 -114.610 93.890 ;
        RECT -110.730 92.760 -110.540 93.890 ;
        RECT -104.880 92.760 -104.690 93.890 ;
        RECT -100.810 92.760 -100.620 93.890 ;
        RECT -94.960 92.760 -94.770 93.890 ;
        RECT -90.890 92.760 -90.700 93.890 ;
        RECT -85.040 92.760 -84.850 93.890 ;
        RECT -80.970 92.760 -80.780 93.890 ;
        RECT -75.120 92.760 -74.930 93.890 ;
        RECT -71.050 92.760 -70.860 93.890 ;
        RECT -65.200 92.760 -65.010 93.890 ;
        RECT -61.130 92.760 -60.940 93.890 ;
        RECT -55.280 92.760 -55.090 93.890 ;
        RECT -51.210 92.760 -51.020 93.890 ;
        RECT -45.360 92.760 -45.170 93.890 ;
        RECT -41.290 92.760 -41.100 93.890 ;
        RECT -35.440 92.760 -35.250 93.890 ;
        RECT -31.370 92.760 -31.180 93.890 ;
        RECT -25.520 92.760 -25.330 93.890 ;
        RECT -21.450 92.760 -21.260 93.890 ;
        RECT -15.600 92.760 -15.410 93.890 ;
        RECT -11.530 92.760 -11.340 93.890 ;
        RECT -5.680 92.760 -5.490 93.890 ;
        RECT -1.610 92.760 -1.420 93.890 ;
        RECT 4.240 92.760 4.430 93.890 ;
        RECT 8.310 92.760 8.500 93.890 ;
        RECT 14.160 92.760 14.350 93.890 ;
        RECT 18.230 92.760 18.420 93.890 ;
        RECT 24.080 92.760 24.270 93.890 ;
        RECT 24.600 93.090 26.440 93.570 ;
        RECT -290.050 92.610 -288.110 92.760 ;
        RECT -290.050 92.460 -289.710 92.610 ;
        RECT -290.050 92.260 -289.730 92.290 ;
        RECT -290.050 92.120 -289.230 92.260 ;
        RECT -290.050 92.010 -289.730 92.120 ;
        RECT -289.390 91.330 -289.230 92.120 ;
        RECT -288.270 91.820 -288.110 92.610 ;
        RECT -284.430 92.610 -282.490 92.760 ;
        RECT -287.770 91.820 -287.450 91.930 ;
        RECT -288.270 91.680 -287.450 91.820 ;
        RECT -287.770 91.650 -287.450 91.680 ;
        RECT -285.090 91.820 -284.770 91.930 ;
        RECT -284.430 91.820 -284.270 92.610 ;
        RECT -282.830 92.460 -282.490 92.610 ;
        RECT -280.130 92.610 -278.190 92.760 ;
        RECT -280.130 92.460 -279.790 92.610 ;
        RECT -282.810 92.260 -282.490 92.290 ;
        RECT -285.090 91.680 -284.270 91.820 ;
        RECT -283.310 92.120 -282.490 92.260 ;
        RECT -285.090 91.650 -284.770 91.680 ;
        RECT -287.790 91.330 -287.450 91.480 ;
        RECT -289.390 91.180 -287.450 91.330 ;
        RECT -285.090 91.330 -284.750 91.480 ;
        RECT -283.310 91.330 -283.150 92.120 ;
        RECT -282.810 92.010 -282.490 92.120 ;
        RECT -280.130 92.260 -279.810 92.290 ;
        RECT -280.130 92.120 -279.310 92.260 ;
        RECT -280.130 92.010 -279.810 92.120 ;
        RECT -285.090 91.180 -283.150 91.330 ;
        RECT -279.470 91.330 -279.310 92.120 ;
        RECT -278.350 91.820 -278.190 92.610 ;
        RECT -274.510 92.610 -272.570 92.760 ;
        RECT -277.850 91.820 -277.530 91.930 ;
        RECT -278.350 91.680 -277.530 91.820 ;
        RECT -277.850 91.650 -277.530 91.680 ;
        RECT -275.170 91.820 -274.850 91.930 ;
        RECT -274.510 91.820 -274.350 92.610 ;
        RECT -272.910 92.460 -272.570 92.610 ;
        RECT -270.210 92.610 -268.270 92.760 ;
        RECT -270.210 92.460 -269.870 92.610 ;
        RECT -272.890 92.260 -272.570 92.290 ;
        RECT -275.170 91.680 -274.350 91.820 ;
        RECT -273.390 92.120 -272.570 92.260 ;
        RECT -275.170 91.650 -274.850 91.680 ;
        RECT -277.870 91.330 -277.530 91.480 ;
        RECT -279.470 91.180 -277.530 91.330 ;
        RECT -275.170 91.330 -274.830 91.480 ;
        RECT -273.390 91.330 -273.230 92.120 ;
        RECT -272.890 92.010 -272.570 92.120 ;
        RECT -270.210 92.260 -269.890 92.290 ;
        RECT -270.210 92.120 -269.390 92.260 ;
        RECT -270.210 92.010 -269.890 92.120 ;
        RECT -275.170 91.180 -273.230 91.330 ;
        RECT -269.550 91.330 -269.390 92.120 ;
        RECT -268.430 91.820 -268.270 92.610 ;
        RECT -264.590 92.610 -262.650 92.760 ;
        RECT -267.930 91.820 -267.610 91.930 ;
        RECT -268.430 91.680 -267.610 91.820 ;
        RECT -267.930 91.650 -267.610 91.680 ;
        RECT -265.250 91.820 -264.930 91.930 ;
        RECT -264.590 91.820 -264.430 92.610 ;
        RECT -262.990 92.460 -262.650 92.610 ;
        RECT -260.290 92.610 -258.350 92.760 ;
        RECT -260.290 92.460 -259.950 92.610 ;
        RECT -262.970 92.260 -262.650 92.290 ;
        RECT -265.250 91.680 -264.430 91.820 ;
        RECT -263.470 92.120 -262.650 92.260 ;
        RECT -265.250 91.650 -264.930 91.680 ;
        RECT -267.950 91.330 -267.610 91.480 ;
        RECT -269.550 91.180 -267.610 91.330 ;
        RECT -265.250 91.330 -264.910 91.480 ;
        RECT -263.470 91.330 -263.310 92.120 ;
        RECT -262.970 92.010 -262.650 92.120 ;
        RECT -260.290 92.260 -259.970 92.290 ;
        RECT -260.290 92.120 -259.470 92.260 ;
        RECT -260.290 92.010 -259.970 92.120 ;
        RECT -265.250 91.180 -263.310 91.330 ;
        RECT -259.630 91.330 -259.470 92.120 ;
        RECT -258.510 91.820 -258.350 92.610 ;
        RECT -254.670 92.610 -252.730 92.760 ;
        RECT -258.010 91.820 -257.690 91.930 ;
        RECT -258.510 91.680 -257.690 91.820 ;
        RECT -258.010 91.650 -257.690 91.680 ;
        RECT -255.330 91.820 -255.010 91.930 ;
        RECT -254.670 91.820 -254.510 92.610 ;
        RECT -253.070 92.460 -252.730 92.610 ;
        RECT -250.370 92.610 -248.430 92.760 ;
        RECT -250.370 92.460 -250.030 92.610 ;
        RECT -253.050 92.260 -252.730 92.290 ;
        RECT -255.330 91.680 -254.510 91.820 ;
        RECT -253.550 92.120 -252.730 92.260 ;
        RECT -255.330 91.650 -255.010 91.680 ;
        RECT -258.030 91.330 -257.690 91.480 ;
        RECT -259.630 91.180 -257.690 91.330 ;
        RECT -255.330 91.330 -254.990 91.480 ;
        RECT -253.550 91.330 -253.390 92.120 ;
        RECT -253.050 92.010 -252.730 92.120 ;
        RECT -250.370 92.260 -250.050 92.290 ;
        RECT -250.370 92.120 -249.550 92.260 ;
        RECT -250.370 92.010 -250.050 92.120 ;
        RECT -255.330 91.180 -253.390 91.330 ;
        RECT -249.710 91.330 -249.550 92.120 ;
        RECT -248.590 91.820 -248.430 92.610 ;
        RECT -244.750 92.610 -242.810 92.760 ;
        RECT -248.090 91.820 -247.770 91.930 ;
        RECT -248.590 91.680 -247.770 91.820 ;
        RECT -248.090 91.650 -247.770 91.680 ;
        RECT -245.410 91.820 -245.090 91.930 ;
        RECT -244.750 91.820 -244.590 92.610 ;
        RECT -243.150 92.460 -242.810 92.610 ;
        RECT -240.450 92.610 -238.510 92.760 ;
        RECT -240.450 92.460 -240.110 92.610 ;
        RECT -243.130 92.260 -242.810 92.290 ;
        RECT -245.410 91.680 -244.590 91.820 ;
        RECT -243.630 92.120 -242.810 92.260 ;
        RECT -245.410 91.650 -245.090 91.680 ;
        RECT -248.110 91.330 -247.770 91.480 ;
        RECT -249.710 91.180 -247.770 91.330 ;
        RECT -245.410 91.330 -245.070 91.480 ;
        RECT -243.630 91.330 -243.470 92.120 ;
        RECT -243.130 92.010 -242.810 92.120 ;
        RECT -240.450 92.260 -240.130 92.290 ;
        RECT -240.450 92.120 -239.630 92.260 ;
        RECT -240.450 92.010 -240.130 92.120 ;
        RECT -245.410 91.180 -243.470 91.330 ;
        RECT -239.790 91.330 -239.630 92.120 ;
        RECT -238.670 91.820 -238.510 92.610 ;
        RECT -234.830 92.610 -232.890 92.760 ;
        RECT -238.170 91.820 -237.850 91.930 ;
        RECT -238.670 91.680 -237.850 91.820 ;
        RECT -238.170 91.650 -237.850 91.680 ;
        RECT -235.490 91.820 -235.170 91.930 ;
        RECT -234.830 91.820 -234.670 92.610 ;
        RECT -233.230 92.460 -232.890 92.610 ;
        RECT -230.530 92.610 -228.590 92.760 ;
        RECT -230.530 92.460 -230.190 92.610 ;
        RECT -233.210 92.260 -232.890 92.290 ;
        RECT -235.490 91.680 -234.670 91.820 ;
        RECT -233.710 92.120 -232.890 92.260 ;
        RECT -235.490 91.650 -235.170 91.680 ;
        RECT -238.190 91.330 -237.850 91.480 ;
        RECT -239.790 91.180 -237.850 91.330 ;
        RECT -235.490 91.330 -235.150 91.480 ;
        RECT -233.710 91.330 -233.550 92.120 ;
        RECT -233.210 92.010 -232.890 92.120 ;
        RECT -230.530 92.260 -230.210 92.290 ;
        RECT -230.530 92.120 -229.710 92.260 ;
        RECT -230.530 92.010 -230.210 92.120 ;
        RECT -235.490 91.180 -233.550 91.330 ;
        RECT -229.870 91.330 -229.710 92.120 ;
        RECT -228.750 91.820 -228.590 92.610 ;
        RECT -224.910 92.610 -222.970 92.760 ;
        RECT -228.250 91.820 -227.930 91.930 ;
        RECT -228.750 91.680 -227.930 91.820 ;
        RECT -228.250 91.650 -227.930 91.680 ;
        RECT -225.570 91.820 -225.250 91.930 ;
        RECT -224.910 91.820 -224.750 92.610 ;
        RECT -223.310 92.460 -222.970 92.610 ;
        RECT -220.610 92.610 -218.670 92.760 ;
        RECT -220.610 92.460 -220.270 92.610 ;
        RECT -223.290 92.260 -222.970 92.290 ;
        RECT -225.570 91.680 -224.750 91.820 ;
        RECT -223.790 92.120 -222.970 92.260 ;
        RECT -225.570 91.650 -225.250 91.680 ;
        RECT -228.270 91.330 -227.930 91.480 ;
        RECT -229.870 91.180 -227.930 91.330 ;
        RECT -225.570 91.330 -225.230 91.480 ;
        RECT -223.790 91.330 -223.630 92.120 ;
        RECT -223.290 92.010 -222.970 92.120 ;
        RECT -220.610 92.260 -220.290 92.290 ;
        RECT -220.610 92.120 -219.790 92.260 ;
        RECT -220.610 92.010 -220.290 92.120 ;
        RECT -225.570 91.180 -223.630 91.330 ;
        RECT -219.950 91.330 -219.790 92.120 ;
        RECT -218.830 91.820 -218.670 92.610 ;
        RECT -214.990 92.610 -213.050 92.760 ;
        RECT -218.330 91.820 -218.010 91.930 ;
        RECT -218.830 91.680 -218.010 91.820 ;
        RECT -218.330 91.650 -218.010 91.680 ;
        RECT -215.650 91.820 -215.330 91.930 ;
        RECT -214.990 91.820 -214.830 92.610 ;
        RECT -213.390 92.460 -213.050 92.610 ;
        RECT -210.690 92.610 -208.750 92.760 ;
        RECT -210.690 92.460 -210.350 92.610 ;
        RECT -213.370 92.260 -213.050 92.290 ;
        RECT -215.650 91.680 -214.830 91.820 ;
        RECT -213.870 92.120 -213.050 92.260 ;
        RECT -215.650 91.650 -215.330 91.680 ;
        RECT -218.350 91.330 -218.010 91.480 ;
        RECT -219.950 91.180 -218.010 91.330 ;
        RECT -215.650 91.330 -215.310 91.480 ;
        RECT -213.870 91.330 -213.710 92.120 ;
        RECT -213.370 92.010 -213.050 92.120 ;
        RECT -210.690 92.260 -210.370 92.290 ;
        RECT -210.690 92.120 -209.870 92.260 ;
        RECT -210.690 92.010 -210.370 92.120 ;
        RECT -215.650 91.180 -213.710 91.330 ;
        RECT -210.030 91.330 -209.870 92.120 ;
        RECT -208.910 91.820 -208.750 92.610 ;
        RECT -205.070 92.610 -203.130 92.760 ;
        RECT -208.410 91.820 -208.090 91.930 ;
        RECT -208.910 91.680 -208.090 91.820 ;
        RECT -208.410 91.650 -208.090 91.680 ;
        RECT -205.730 91.820 -205.410 91.930 ;
        RECT -205.070 91.820 -204.910 92.610 ;
        RECT -203.470 92.460 -203.130 92.610 ;
        RECT -200.770 92.610 -198.830 92.760 ;
        RECT -200.770 92.460 -200.430 92.610 ;
        RECT -203.450 92.260 -203.130 92.290 ;
        RECT -205.730 91.680 -204.910 91.820 ;
        RECT -203.950 92.120 -203.130 92.260 ;
        RECT -205.730 91.650 -205.410 91.680 ;
        RECT -208.430 91.330 -208.090 91.480 ;
        RECT -210.030 91.180 -208.090 91.330 ;
        RECT -205.730 91.330 -205.390 91.480 ;
        RECT -203.950 91.330 -203.790 92.120 ;
        RECT -203.450 92.010 -203.130 92.120 ;
        RECT -200.770 92.260 -200.450 92.290 ;
        RECT -200.770 92.120 -199.950 92.260 ;
        RECT -200.770 92.010 -200.450 92.120 ;
        RECT -205.730 91.180 -203.790 91.330 ;
        RECT -200.110 91.330 -199.950 92.120 ;
        RECT -198.990 91.820 -198.830 92.610 ;
        RECT -195.150 92.610 -193.210 92.760 ;
        RECT -198.490 91.820 -198.170 91.930 ;
        RECT -198.990 91.680 -198.170 91.820 ;
        RECT -198.490 91.650 -198.170 91.680 ;
        RECT -195.810 91.820 -195.490 91.930 ;
        RECT -195.150 91.820 -194.990 92.610 ;
        RECT -193.550 92.460 -193.210 92.610 ;
        RECT -190.850 92.610 -188.910 92.760 ;
        RECT -190.850 92.460 -190.510 92.610 ;
        RECT -193.530 92.260 -193.210 92.290 ;
        RECT -195.810 91.680 -194.990 91.820 ;
        RECT -194.030 92.120 -193.210 92.260 ;
        RECT -195.810 91.650 -195.490 91.680 ;
        RECT -198.510 91.330 -198.170 91.480 ;
        RECT -200.110 91.180 -198.170 91.330 ;
        RECT -195.810 91.330 -195.470 91.480 ;
        RECT -194.030 91.330 -193.870 92.120 ;
        RECT -193.530 92.010 -193.210 92.120 ;
        RECT -190.850 92.260 -190.530 92.290 ;
        RECT -190.850 92.120 -190.030 92.260 ;
        RECT -190.850 92.010 -190.530 92.120 ;
        RECT -195.810 91.180 -193.870 91.330 ;
        RECT -190.190 91.330 -190.030 92.120 ;
        RECT -189.070 91.820 -188.910 92.610 ;
        RECT -185.230 92.610 -183.290 92.760 ;
        RECT -188.570 91.820 -188.250 91.930 ;
        RECT -189.070 91.680 -188.250 91.820 ;
        RECT -188.570 91.650 -188.250 91.680 ;
        RECT -185.890 91.820 -185.570 91.930 ;
        RECT -185.230 91.820 -185.070 92.610 ;
        RECT -183.630 92.460 -183.290 92.610 ;
        RECT -180.930 92.610 -178.990 92.760 ;
        RECT -180.930 92.460 -180.590 92.610 ;
        RECT -183.610 92.260 -183.290 92.290 ;
        RECT -185.890 91.680 -185.070 91.820 ;
        RECT -184.110 92.120 -183.290 92.260 ;
        RECT -185.890 91.650 -185.570 91.680 ;
        RECT -188.590 91.330 -188.250 91.480 ;
        RECT -190.190 91.180 -188.250 91.330 ;
        RECT -185.890 91.330 -185.550 91.480 ;
        RECT -184.110 91.330 -183.950 92.120 ;
        RECT -183.610 92.010 -183.290 92.120 ;
        RECT -180.930 92.260 -180.610 92.290 ;
        RECT -180.930 92.120 -180.110 92.260 ;
        RECT -180.930 92.010 -180.610 92.120 ;
        RECT -185.890 91.180 -183.950 91.330 ;
        RECT -180.270 91.330 -180.110 92.120 ;
        RECT -179.150 91.820 -178.990 92.610 ;
        RECT -175.310 92.610 -173.370 92.760 ;
        RECT -178.650 91.820 -178.330 91.930 ;
        RECT -179.150 91.680 -178.330 91.820 ;
        RECT -178.650 91.650 -178.330 91.680 ;
        RECT -175.970 91.820 -175.650 91.930 ;
        RECT -175.310 91.820 -175.150 92.610 ;
        RECT -173.710 92.460 -173.370 92.610 ;
        RECT -171.010 92.610 -169.070 92.760 ;
        RECT -171.010 92.460 -170.670 92.610 ;
        RECT -173.690 92.260 -173.370 92.290 ;
        RECT -175.970 91.680 -175.150 91.820 ;
        RECT -174.190 92.120 -173.370 92.260 ;
        RECT -175.970 91.650 -175.650 91.680 ;
        RECT -178.670 91.330 -178.330 91.480 ;
        RECT -180.270 91.180 -178.330 91.330 ;
        RECT -175.970 91.330 -175.630 91.480 ;
        RECT -174.190 91.330 -174.030 92.120 ;
        RECT -173.690 92.010 -173.370 92.120 ;
        RECT -171.010 92.260 -170.690 92.290 ;
        RECT -171.010 92.120 -170.190 92.260 ;
        RECT -171.010 92.010 -170.690 92.120 ;
        RECT -175.970 91.180 -174.030 91.330 ;
        RECT -170.350 91.330 -170.190 92.120 ;
        RECT -169.230 91.820 -169.070 92.610 ;
        RECT -165.390 92.610 -163.450 92.760 ;
        RECT -168.730 91.820 -168.410 91.930 ;
        RECT -169.230 91.680 -168.410 91.820 ;
        RECT -168.730 91.650 -168.410 91.680 ;
        RECT -166.050 91.820 -165.730 91.930 ;
        RECT -165.390 91.820 -165.230 92.610 ;
        RECT -163.790 92.460 -163.450 92.610 ;
        RECT -161.090 92.610 -159.150 92.760 ;
        RECT -161.090 92.460 -160.750 92.610 ;
        RECT -163.770 92.260 -163.450 92.290 ;
        RECT -166.050 91.680 -165.230 91.820 ;
        RECT -164.270 92.120 -163.450 92.260 ;
        RECT -166.050 91.650 -165.730 91.680 ;
        RECT -168.750 91.330 -168.410 91.480 ;
        RECT -170.350 91.180 -168.410 91.330 ;
        RECT -166.050 91.330 -165.710 91.480 ;
        RECT -164.270 91.330 -164.110 92.120 ;
        RECT -163.770 92.010 -163.450 92.120 ;
        RECT -161.090 92.260 -160.770 92.290 ;
        RECT -161.090 92.120 -160.270 92.260 ;
        RECT -161.090 92.010 -160.770 92.120 ;
        RECT -166.050 91.180 -164.110 91.330 ;
        RECT -160.430 91.330 -160.270 92.120 ;
        RECT -159.310 91.820 -159.150 92.610 ;
        RECT -155.470 92.610 -153.530 92.760 ;
        RECT -158.810 91.820 -158.490 91.930 ;
        RECT -159.310 91.680 -158.490 91.820 ;
        RECT -158.810 91.650 -158.490 91.680 ;
        RECT -156.130 91.820 -155.810 91.930 ;
        RECT -155.470 91.820 -155.310 92.610 ;
        RECT -153.870 92.460 -153.530 92.610 ;
        RECT -151.170 92.610 -149.230 92.760 ;
        RECT -151.170 92.460 -150.830 92.610 ;
        RECT -153.850 92.260 -153.530 92.290 ;
        RECT -156.130 91.680 -155.310 91.820 ;
        RECT -154.350 92.120 -153.530 92.260 ;
        RECT -156.130 91.650 -155.810 91.680 ;
        RECT -158.830 91.330 -158.490 91.480 ;
        RECT -160.430 91.180 -158.490 91.330 ;
        RECT -156.130 91.330 -155.790 91.480 ;
        RECT -154.350 91.330 -154.190 92.120 ;
        RECT -153.850 92.010 -153.530 92.120 ;
        RECT -151.170 92.260 -150.850 92.290 ;
        RECT -151.170 92.120 -150.350 92.260 ;
        RECT -151.170 92.010 -150.850 92.120 ;
        RECT -156.130 91.180 -154.190 91.330 ;
        RECT -150.510 91.330 -150.350 92.120 ;
        RECT -149.390 91.820 -149.230 92.610 ;
        RECT -145.550 92.610 -143.610 92.760 ;
        RECT -148.890 91.820 -148.570 91.930 ;
        RECT -149.390 91.680 -148.570 91.820 ;
        RECT -148.890 91.650 -148.570 91.680 ;
        RECT -146.210 91.820 -145.890 91.930 ;
        RECT -145.550 91.820 -145.390 92.610 ;
        RECT -143.950 92.460 -143.610 92.610 ;
        RECT -141.250 92.610 -139.310 92.760 ;
        RECT -141.250 92.460 -140.910 92.610 ;
        RECT -143.930 92.260 -143.610 92.290 ;
        RECT -146.210 91.680 -145.390 91.820 ;
        RECT -144.430 92.120 -143.610 92.260 ;
        RECT -146.210 91.650 -145.890 91.680 ;
        RECT -148.910 91.330 -148.570 91.480 ;
        RECT -150.510 91.180 -148.570 91.330 ;
        RECT -146.210 91.330 -145.870 91.480 ;
        RECT -144.430 91.330 -144.270 92.120 ;
        RECT -143.930 92.010 -143.610 92.120 ;
        RECT -141.250 92.260 -140.930 92.290 ;
        RECT -141.250 92.120 -140.430 92.260 ;
        RECT -141.250 92.010 -140.930 92.120 ;
        RECT -146.210 91.180 -144.270 91.330 ;
        RECT -140.590 91.330 -140.430 92.120 ;
        RECT -139.470 91.820 -139.310 92.610 ;
        RECT -135.630 92.610 -133.690 92.760 ;
        RECT -138.970 91.820 -138.650 91.930 ;
        RECT -139.470 91.680 -138.650 91.820 ;
        RECT -138.970 91.650 -138.650 91.680 ;
        RECT -136.290 91.820 -135.970 91.930 ;
        RECT -135.630 91.820 -135.470 92.610 ;
        RECT -134.030 92.460 -133.690 92.610 ;
        RECT -131.330 92.610 -129.390 92.760 ;
        RECT -131.330 92.460 -130.990 92.610 ;
        RECT -134.010 92.260 -133.690 92.290 ;
        RECT -136.290 91.680 -135.470 91.820 ;
        RECT -134.510 92.120 -133.690 92.260 ;
        RECT -136.290 91.650 -135.970 91.680 ;
        RECT -138.990 91.330 -138.650 91.480 ;
        RECT -140.590 91.180 -138.650 91.330 ;
        RECT -136.290 91.330 -135.950 91.480 ;
        RECT -134.510 91.330 -134.350 92.120 ;
        RECT -134.010 92.010 -133.690 92.120 ;
        RECT -131.330 92.260 -131.010 92.290 ;
        RECT -131.330 92.120 -130.510 92.260 ;
        RECT -131.330 92.010 -131.010 92.120 ;
        RECT -136.290 91.180 -134.350 91.330 ;
        RECT -130.670 91.330 -130.510 92.120 ;
        RECT -129.550 91.820 -129.390 92.610 ;
        RECT -125.710 92.610 -123.770 92.760 ;
        RECT -129.050 91.820 -128.730 91.930 ;
        RECT -129.550 91.680 -128.730 91.820 ;
        RECT -129.050 91.650 -128.730 91.680 ;
        RECT -126.370 91.820 -126.050 91.930 ;
        RECT -125.710 91.820 -125.550 92.610 ;
        RECT -124.110 92.460 -123.770 92.610 ;
        RECT -121.410 92.610 -119.470 92.760 ;
        RECT -121.410 92.460 -121.070 92.610 ;
        RECT -124.090 92.260 -123.770 92.290 ;
        RECT -126.370 91.680 -125.550 91.820 ;
        RECT -124.590 92.120 -123.770 92.260 ;
        RECT -126.370 91.650 -126.050 91.680 ;
        RECT -129.070 91.330 -128.730 91.480 ;
        RECT -130.670 91.180 -128.730 91.330 ;
        RECT -126.370 91.330 -126.030 91.480 ;
        RECT -124.590 91.330 -124.430 92.120 ;
        RECT -124.090 92.010 -123.770 92.120 ;
        RECT -121.410 92.260 -121.090 92.290 ;
        RECT -121.410 92.120 -120.590 92.260 ;
        RECT -121.410 92.010 -121.090 92.120 ;
        RECT -126.370 91.180 -124.430 91.330 ;
        RECT -120.750 91.330 -120.590 92.120 ;
        RECT -119.630 91.820 -119.470 92.610 ;
        RECT -115.790 92.610 -113.850 92.760 ;
        RECT -119.130 91.820 -118.810 91.930 ;
        RECT -119.630 91.680 -118.810 91.820 ;
        RECT -119.130 91.650 -118.810 91.680 ;
        RECT -116.450 91.820 -116.130 91.930 ;
        RECT -115.790 91.820 -115.630 92.610 ;
        RECT -114.190 92.460 -113.850 92.610 ;
        RECT -111.490 92.610 -109.550 92.760 ;
        RECT -111.490 92.460 -111.150 92.610 ;
        RECT -114.170 92.260 -113.850 92.290 ;
        RECT -116.450 91.680 -115.630 91.820 ;
        RECT -114.670 92.120 -113.850 92.260 ;
        RECT -116.450 91.650 -116.130 91.680 ;
        RECT -119.150 91.330 -118.810 91.480 ;
        RECT -120.750 91.180 -118.810 91.330 ;
        RECT -116.450 91.330 -116.110 91.480 ;
        RECT -114.670 91.330 -114.510 92.120 ;
        RECT -114.170 92.010 -113.850 92.120 ;
        RECT -111.490 92.260 -111.170 92.290 ;
        RECT -111.490 92.120 -110.670 92.260 ;
        RECT -111.490 92.010 -111.170 92.120 ;
        RECT -116.450 91.180 -114.510 91.330 ;
        RECT -110.830 91.330 -110.670 92.120 ;
        RECT -109.710 91.820 -109.550 92.610 ;
        RECT -105.870 92.610 -103.930 92.760 ;
        RECT -109.210 91.820 -108.890 91.930 ;
        RECT -109.710 91.680 -108.890 91.820 ;
        RECT -109.210 91.650 -108.890 91.680 ;
        RECT -106.530 91.820 -106.210 91.930 ;
        RECT -105.870 91.820 -105.710 92.610 ;
        RECT -104.270 92.460 -103.930 92.610 ;
        RECT -101.570 92.610 -99.630 92.760 ;
        RECT -101.570 92.460 -101.230 92.610 ;
        RECT -104.250 92.260 -103.930 92.290 ;
        RECT -106.530 91.680 -105.710 91.820 ;
        RECT -104.750 92.120 -103.930 92.260 ;
        RECT -106.530 91.650 -106.210 91.680 ;
        RECT -109.230 91.330 -108.890 91.480 ;
        RECT -110.830 91.180 -108.890 91.330 ;
        RECT -106.530 91.330 -106.190 91.480 ;
        RECT -104.750 91.330 -104.590 92.120 ;
        RECT -104.250 92.010 -103.930 92.120 ;
        RECT -101.570 92.260 -101.250 92.290 ;
        RECT -101.570 92.120 -100.750 92.260 ;
        RECT -101.570 92.010 -101.250 92.120 ;
        RECT -106.530 91.180 -104.590 91.330 ;
        RECT -100.910 91.330 -100.750 92.120 ;
        RECT -99.790 91.820 -99.630 92.610 ;
        RECT -95.950 92.610 -94.010 92.760 ;
        RECT -99.290 91.820 -98.970 91.930 ;
        RECT -99.790 91.680 -98.970 91.820 ;
        RECT -99.290 91.650 -98.970 91.680 ;
        RECT -96.610 91.820 -96.290 91.930 ;
        RECT -95.950 91.820 -95.790 92.610 ;
        RECT -94.350 92.460 -94.010 92.610 ;
        RECT -91.650 92.610 -89.710 92.760 ;
        RECT -91.650 92.460 -91.310 92.610 ;
        RECT -94.330 92.260 -94.010 92.290 ;
        RECT -96.610 91.680 -95.790 91.820 ;
        RECT -94.830 92.120 -94.010 92.260 ;
        RECT -96.610 91.650 -96.290 91.680 ;
        RECT -99.310 91.330 -98.970 91.480 ;
        RECT -100.910 91.180 -98.970 91.330 ;
        RECT -96.610 91.330 -96.270 91.480 ;
        RECT -94.830 91.330 -94.670 92.120 ;
        RECT -94.330 92.010 -94.010 92.120 ;
        RECT -91.650 92.260 -91.330 92.290 ;
        RECT -91.650 92.120 -90.830 92.260 ;
        RECT -91.650 92.010 -91.330 92.120 ;
        RECT -96.610 91.180 -94.670 91.330 ;
        RECT -90.990 91.330 -90.830 92.120 ;
        RECT -89.870 91.820 -89.710 92.610 ;
        RECT -86.030 92.610 -84.090 92.760 ;
        RECT -89.370 91.820 -89.050 91.930 ;
        RECT -89.870 91.680 -89.050 91.820 ;
        RECT -89.370 91.650 -89.050 91.680 ;
        RECT -86.690 91.820 -86.370 91.930 ;
        RECT -86.030 91.820 -85.870 92.610 ;
        RECT -84.430 92.460 -84.090 92.610 ;
        RECT -81.730 92.610 -79.790 92.760 ;
        RECT -81.730 92.460 -81.390 92.610 ;
        RECT -84.410 92.260 -84.090 92.290 ;
        RECT -86.690 91.680 -85.870 91.820 ;
        RECT -84.910 92.120 -84.090 92.260 ;
        RECT -86.690 91.650 -86.370 91.680 ;
        RECT -89.390 91.330 -89.050 91.480 ;
        RECT -90.990 91.180 -89.050 91.330 ;
        RECT -86.690 91.330 -86.350 91.480 ;
        RECT -84.910 91.330 -84.750 92.120 ;
        RECT -84.410 92.010 -84.090 92.120 ;
        RECT -81.730 92.260 -81.410 92.290 ;
        RECT -81.730 92.120 -80.910 92.260 ;
        RECT -81.730 92.010 -81.410 92.120 ;
        RECT -86.690 91.180 -84.750 91.330 ;
        RECT -81.070 91.330 -80.910 92.120 ;
        RECT -79.950 91.820 -79.790 92.610 ;
        RECT -76.110 92.610 -74.170 92.760 ;
        RECT -79.450 91.820 -79.130 91.930 ;
        RECT -79.950 91.680 -79.130 91.820 ;
        RECT -79.450 91.650 -79.130 91.680 ;
        RECT -76.770 91.820 -76.450 91.930 ;
        RECT -76.110 91.820 -75.950 92.610 ;
        RECT -74.510 92.460 -74.170 92.610 ;
        RECT -71.810 92.610 -69.870 92.760 ;
        RECT -71.810 92.460 -71.470 92.610 ;
        RECT -74.490 92.260 -74.170 92.290 ;
        RECT -76.770 91.680 -75.950 91.820 ;
        RECT -74.990 92.120 -74.170 92.260 ;
        RECT -76.770 91.650 -76.450 91.680 ;
        RECT -79.470 91.330 -79.130 91.480 ;
        RECT -81.070 91.180 -79.130 91.330 ;
        RECT -76.770 91.330 -76.430 91.480 ;
        RECT -74.990 91.330 -74.830 92.120 ;
        RECT -74.490 92.010 -74.170 92.120 ;
        RECT -71.810 92.260 -71.490 92.290 ;
        RECT -71.810 92.120 -70.990 92.260 ;
        RECT -71.810 92.010 -71.490 92.120 ;
        RECT -76.770 91.180 -74.830 91.330 ;
        RECT -71.150 91.330 -70.990 92.120 ;
        RECT -70.030 91.820 -69.870 92.610 ;
        RECT -66.190 92.610 -64.250 92.760 ;
        RECT -69.530 91.820 -69.210 91.930 ;
        RECT -70.030 91.680 -69.210 91.820 ;
        RECT -69.530 91.650 -69.210 91.680 ;
        RECT -66.850 91.820 -66.530 91.930 ;
        RECT -66.190 91.820 -66.030 92.610 ;
        RECT -64.590 92.460 -64.250 92.610 ;
        RECT -61.890 92.610 -59.950 92.760 ;
        RECT -61.890 92.460 -61.550 92.610 ;
        RECT -64.570 92.260 -64.250 92.290 ;
        RECT -66.850 91.680 -66.030 91.820 ;
        RECT -65.070 92.120 -64.250 92.260 ;
        RECT -66.850 91.650 -66.530 91.680 ;
        RECT -69.550 91.330 -69.210 91.480 ;
        RECT -71.150 91.180 -69.210 91.330 ;
        RECT -66.850 91.330 -66.510 91.480 ;
        RECT -65.070 91.330 -64.910 92.120 ;
        RECT -64.570 92.010 -64.250 92.120 ;
        RECT -61.890 92.260 -61.570 92.290 ;
        RECT -61.890 92.120 -61.070 92.260 ;
        RECT -61.890 92.010 -61.570 92.120 ;
        RECT -66.850 91.180 -64.910 91.330 ;
        RECT -61.230 91.330 -61.070 92.120 ;
        RECT -60.110 91.820 -59.950 92.610 ;
        RECT -56.270 92.610 -54.330 92.760 ;
        RECT -59.610 91.820 -59.290 91.930 ;
        RECT -60.110 91.680 -59.290 91.820 ;
        RECT -59.610 91.650 -59.290 91.680 ;
        RECT -56.930 91.820 -56.610 91.930 ;
        RECT -56.270 91.820 -56.110 92.610 ;
        RECT -54.670 92.460 -54.330 92.610 ;
        RECT -51.970 92.610 -50.030 92.760 ;
        RECT -51.970 92.460 -51.630 92.610 ;
        RECT -54.650 92.260 -54.330 92.290 ;
        RECT -56.930 91.680 -56.110 91.820 ;
        RECT -55.150 92.120 -54.330 92.260 ;
        RECT -56.930 91.650 -56.610 91.680 ;
        RECT -59.630 91.330 -59.290 91.480 ;
        RECT -61.230 91.180 -59.290 91.330 ;
        RECT -56.930 91.330 -56.590 91.480 ;
        RECT -55.150 91.330 -54.990 92.120 ;
        RECT -54.650 92.010 -54.330 92.120 ;
        RECT -51.970 92.260 -51.650 92.290 ;
        RECT -51.970 92.120 -51.150 92.260 ;
        RECT -51.970 92.010 -51.650 92.120 ;
        RECT -56.930 91.180 -54.990 91.330 ;
        RECT -51.310 91.330 -51.150 92.120 ;
        RECT -50.190 91.820 -50.030 92.610 ;
        RECT -46.350 92.610 -44.410 92.760 ;
        RECT -49.690 91.820 -49.370 91.930 ;
        RECT -50.190 91.680 -49.370 91.820 ;
        RECT -49.690 91.650 -49.370 91.680 ;
        RECT -47.010 91.820 -46.690 91.930 ;
        RECT -46.350 91.820 -46.190 92.610 ;
        RECT -44.750 92.460 -44.410 92.610 ;
        RECT -42.050 92.610 -40.110 92.760 ;
        RECT -42.050 92.460 -41.710 92.610 ;
        RECT -44.730 92.260 -44.410 92.290 ;
        RECT -47.010 91.680 -46.190 91.820 ;
        RECT -45.230 92.120 -44.410 92.260 ;
        RECT -47.010 91.650 -46.690 91.680 ;
        RECT -49.710 91.330 -49.370 91.480 ;
        RECT -51.310 91.180 -49.370 91.330 ;
        RECT -47.010 91.330 -46.670 91.480 ;
        RECT -45.230 91.330 -45.070 92.120 ;
        RECT -44.730 92.010 -44.410 92.120 ;
        RECT -42.050 92.260 -41.730 92.290 ;
        RECT -42.050 92.120 -41.230 92.260 ;
        RECT -42.050 92.010 -41.730 92.120 ;
        RECT -47.010 91.180 -45.070 91.330 ;
        RECT -41.390 91.330 -41.230 92.120 ;
        RECT -40.270 91.820 -40.110 92.610 ;
        RECT -36.430 92.610 -34.490 92.760 ;
        RECT -39.770 91.820 -39.450 91.930 ;
        RECT -40.270 91.680 -39.450 91.820 ;
        RECT -39.770 91.650 -39.450 91.680 ;
        RECT -37.090 91.820 -36.770 91.930 ;
        RECT -36.430 91.820 -36.270 92.610 ;
        RECT -34.830 92.460 -34.490 92.610 ;
        RECT -32.130 92.610 -30.190 92.760 ;
        RECT -32.130 92.460 -31.790 92.610 ;
        RECT -34.810 92.260 -34.490 92.290 ;
        RECT -37.090 91.680 -36.270 91.820 ;
        RECT -35.310 92.120 -34.490 92.260 ;
        RECT -37.090 91.650 -36.770 91.680 ;
        RECT -39.790 91.330 -39.450 91.480 ;
        RECT -41.390 91.180 -39.450 91.330 ;
        RECT -37.090 91.330 -36.750 91.480 ;
        RECT -35.310 91.330 -35.150 92.120 ;
        RECT -34.810 92.010 -34.490 92.120 ;
        RECT -32.130 92.260 -31.810 92.290 ;
        RECT -32.130 92.120 -31.310 92.260 ;
        RECT -32.130 92.010 -31.810 92.120 ;
        RECT -37.090 91.180 -35.150 91.330 ;
        RECT -31.470 91.330 -31.310 92.120 ;
        RECT -30.350 91.820 -30.190 92.610 ;
        RECT -26.510 92.610 -24.570 92.760 ;
        RECT -29.850 91.820 -29.530 91.930 ;
        RECT -30.350 91.680 -29.530 91.820 ;
        RECT -29.850 91.650 -29.530 91.680 ;
        RECT -27.170 91.820 -26.850 91.930 ;
        RECT -26.510 91.820 -26.350 92.610 ;
        RECT -24.910 92.460 -24.570 92.610 ;
        RECT -22.210 92.610 -20.270 92.760 ;
        RECT -22.210 92.460 -21.870 92.610 ;
        RECT -24.890 92.260 -24.570 92.290 ;
        RECT -27.170 91.680 -26.350 91.820 ;
        RECT -25.390 92.120 -24.570 92.260 ;
        RECT -27.170 91.650 -26.850 91.680 ;
        RECT -29.870 91.330 -29.530 91.480 ;
        RECT -31.470 91.180 -29.530 91.330 ;
        RECT -27.170 91.330 -26.830 91.480 ;
        RECT -25.390 91.330 -25.230 92.120 ;
        RECT -24.890 92.010 -24.570 92.120 ;
        RECT -22.210 92.260 -21.890 92.290 ;
        RECT -22.210 92.120 -21.390 92.260 ;
        RECT -22.210 92.010 -21.890 92.120 ;
        RECT -27.170 91.180 -25.230 91.330 ;
        RECT -21.550 91.330 -21.390 92.120 ;
        RECT -20.430 91.820 -20.270 92.610 ;
        RECT -16.590 92.610 -14.650 92.760 ;
        RECT -19.930 91.820 -19.610 91.930 ;
        RECT -20.430 91.680 -19.610 91.820 ;
        RECT -19.930 91.650 -19.610 91.680 ;
        RECT -17.250 91.820 -16.930 91.930 ;
        RECT -16.590 91.820 -16.430 92.610 ;
        RECT -14.990 92.460 -14.650 92.610 ;
        RECT -12.290 92.610 -10.350 92.760 ;
        RECT -12.290 92.460 -11.950 92.610 ;
        RECT -14.970 92.260 -14.650 92.290 ;
        RECT -17.250 91.680 -16.430 91.820 ;
        RECT -15.470 92.120 -14.650 92.260 ;
        RECT -17.250 91.650 -16.930 91.680 ;
        RECT -19.950 91.330 -19.610 91.480 ;
        RECT -21.550 91.180 -19.610 91.330 ;
        RECT -17.250 91.330 -16.910 91.480 ;
        RECT -15.470 91.330 -15.310 92.120 ;
        RECT -14.970 92.010 -14.650 92.120 ;
        RECT -12.290 92.260 -11.970 92.290 ;
        RECT -12.290 92.120 -11.470 92.260 ;
        RECT -12.290 92.010 -11.970 92.120 ;
        RECT -17.250 91.180 -15.310 91.330 ;
        RECT -11.630 91.330 -11.470 92.120 ;
        RECT -10.510 91.820 -10.350 92.610 ;
        RECT -6.670 92.610 -4.730 92.760 ;
        RECT -10.010 91.820 -9.690 91.930 ;
        RECT -10.510 91.680 -9.690 91.820 ;
        RECT -10.010 91.650 -9.690 91.680 ;
        RECT -7.330 91.820 -7.010 91.930 ;
        RECT -6.670 91.820 -6.510 92.610 ;
        RECT -5.070 92.460 -4.730 92.610 ;
        RECT -2.370 92.610 -0.430 92.760 ;
        RECT -2.370 92.460 -2.030 92.610 ;
        RECT -5.050 92.260 -4.730 92.290 ;
        RECT -7.330 91.680 -6.510 91.820 ;
        RECT -5.550 92.120 -4.730 92.260 ;
        RECT -7.330 91.650 -7.010 91.680 ;
        RECT -10.030 91.330 -9.690 91.480 ;
        RECT -11.630 91.180 -9.690 91.330 ;
        RECT -7.330 91.330 -6.990 91.480 ;
        RECT -5.550 91.330 -5.390 92.120 ;
        RECT -5.050 92.010 -4.730 92.120 ;
        RECT -2.370 92.260 -2.050 92.290 ;
        RECT -2.370 92.120 -1.550 92.260 ;
        RECT -2.370 92.010 -2.050 92.120 ;
        RECT -7.330 91.180 -5.390 91.330 ;
        RECT -1.710 91.330 -1.550 92.120 ;
        RECT -0.590 91.820 -0.430 92.610 ;
        RECT 3.250 92.610 5.190 92.760 ;
        RECT -0.090 91.820 0.230 91.930 ;
        RECT -0.590 91.680 0.230 91.820 ;
        RECT -0.090 91.650 0.230 91.680 ;
        RECT 2.590 91.820 2.910 91.930 ;
        RECT 3.250 91.820 3.410 92.610 ;
        RECT 4.850 92.460 5.190 92.610 ;
        RECT 7.550 92.610 9.490 92.760 ;
        RECT 7.550 92.460 7.890 92.610 ;
        RECT 4.870 92.260 5.190 92.290 ;
        RECT 2.590 91.680 3.410 91.820 ;
        RECT 4.370 92.120 5.190 92.260 ;
        RECT 2.590 91.650 2.910 91.680 ;
        RECT -0.110 91.330 0.230 91.480 ;
        RECT -1.710 91.180 0.230 91.330 ;
        RECT 2.590 91.330 2.930 91.480 ;
        RECT 4.370 91.330 4.530 92.120 ;
        RECT 4.870 92.010 5.190 92.120 ;
        RECT 7.550 92.260 7.870 92.290 ;
        RECT 7.550 92.120 8.370 92.260 ;
        RECT 7.550 92.010 7.870 92.120 ;
        RECT 2.590 91.180 4.530 91.330 ;
        RECT 8.210 91.330 8.370 92.120 ;
        RECT 9.330 91.820 9.490 92.610 ;
        RECT 13.170 92.610 15.110 92.760 ;
        RECT 9.830 91.820 10.150 91.930 ;
        RECT 9.330 91.680 10.150 91.820 ;
        RECT 9.830 91.650 10.150 91.680 ;
        RECT 12.510 91.820 12.830 91.930 ;
        RECT 13.170 91.820 13.330 92.610 ;
        RECT 14.770 92.460 15.110 92.610 ;
        RECT 17.470 92.610 19.410 92.760 ;
        RECT 17.470 92.460 17.810 92.610 ;
        RECT 14.790 92.260 15.110 92.290 ;
        RECT 12.510 91.680 13.330 91.820 ;
        RECT 14.290 92.120 15.110 92.260 ;
        RECT 12.510 91.650 12.830 91.680 ;
        RECT 9.810 91.330 10.150 91.480 ;
        RECT 8.210 91.180 10.150 91.330 ;
        RECT 12.510 91.330 12.850 91.480 ;
        RECT 14.290 91.330 14.450 92.120 ;
        RECT 14.790 92.010 15.110 92.120 ;
        RECT 17.470 92.260 17.790 92.290 ;
        RECT 17.470 92.120 18.290 92.260 ;
        RECT 17.470 92.010 17.790 92.120 ;
        RECT 12.510 91.180 14.450 91.330 ;
        RECT 18.130 91.330 18.290 92.120 ;
        RECT 19.250 91.820 19.410 92.610 ;
        RECT 23.090 92.610 25.030 92.760 ;
        RECT 19.750 91.820 20.070 91.930 ;
        RECT 19.250 91.680 20.070 91.820 ;
        RECT 19.750 91.650 20.070 91.680 ;
        RECT 22.430 91.820 22.750 91.930 ;
        RECT 23.090 91.820 23.250 92.610 ;
        RECT 24.690 92.460 25.030 92.610 ;
        RECT 24.710 92.260 25.030 92.290 ;
        RECT 22.430 91.680 23.250 91.820 ;
        RECT 24.210 92.120 25.030 92.260 ;
        RECT 22.430 91.650 22.750 91.680 ;
        RECT 19.730 91.330 20.070 91.480 ;
        RECT 18.130 91.180 20.070 91.330 ;
        RECT 22.430 91.330 22.770 91.480 ;
        RECT 24.210 91.330 24.370 92.120 ;
        RECT 24.710 92.010 25.030 92.120 ;
        RECT 22.430 91.180 24.370 91.330 ;
        RECT -291.460 90.370 -289.620 90.850 ;
        RECT -289.700 89.280 -289.220 90.180 ;
        RECT -288.400 90.050 -288.210 91.180 ;
        RECT -284.330 90.050 -284.140 91.180 ;
        RECT -278.480 90.050 -278.290 91.180 ;
        RECT -274.410 90.050 -274.220 91.180 ;
        RECT -268.560 90.050 -268.370 91.180 ;
        RECT -264.490 90.050 -264.300 91.180 ;
        RECT -258.640 90.050 -258.450 91.180 ;
        RECT -254.570 90.050 -254.380 91.180 ;
        RECT -248.720 90.050 -248.530 91.180 ;
        RECT -244.650 90.050 -244.460 91.180 ;
        RECT -238.800 90.050 -238.610 91.180 ;
        RECT -234.730 90.050 -234.540 91.180 ;
        RECT -228.880 90.050 -228.690 91.180 ;
        RECT -224.810 90.050 -224.620 91.180 ;
        RECT -218.960 90.050 -218.770 91.180 ;
        RECT -214.890 90.050 -214.700 91.180 ;
        RECT -209.040 90.050 -208.850 91.180 ;
        RECT -204.970 90.050 -204.780 91.180 ;
        RECT -199.120 90.050 -198.930 91.180 ;
        RECT -195.050 90.050 -194.860 91.180 ;
        RECT -189.200 90.050 -189.010 91.180 ;
        RECT -185.130 90.050 -184.940 91.180 ;
        RECT -179.280 90.050 -179.090 91.180 ;
        RECT -175.210 90.050 -175.020 91.180 ;
        RECT -169.360 90.050 -169.170 91.180 ;
        RECT -165.290 90.050 -165.100 91.180 ;
        RECT -159.440 90.050 -159.250 91.180 ;
        RECT -155.370 90.050 -155.180 91.180 ;
        RECT -149.520 90.050 -149.330 91.180 ;
        RECT -145.450 90.050 -145.260 91.180 ;
        RECT -139.600 90.050 -139.410 91.180 ;
        RECT -135.530 90.050 -135.340 91.180 ;
        RECT -129.680 90.050 -129.490 91.180 ;
        RECT -125.610 90.050 -125.420 91.180 ;
        RECT -119.760 90.050 -119.570 91.180 ;
        RECT -115.690 90.050 -115.500 91.180 ;
        RECT -109.840 90.050 -109.650 91.180 ;
        RECT -105.770 90.050 -105.580 91.180 ;
        RECT -99.920 90.050 -99.730 91.180 ;
        RECT -95.850 90.050 -95.660 91.180 ;
        RECT -90.000 90.050 -89.810 91.180 ;
        RECT -85.930 90.050 -85.740 91.180 ;
        RECT -80.080 90.050 -79.890 91.180 ;
        RECT -76.010 90.050 -75.820 91.180 ;
        RECT -70.160 90.050 -69.970 91.180 ;
        RECT -66.090 90.050 -65.900 91.180 ;
        RECT -60.240 90.050 -60.050 91.180 ;
        RECT -56.170 90.050 -55.980 91.180 ;
        RECT -50.320 90.050 -50.130 91.180 ;
        RECT -46.250 90.050 -46.060 91.180 ;
        RECT -40.400 90.050 -40.210 91.180 ;
        RECT -36.330 90.050 -36.140 91.180 ;
        RECT -30.480 90.050 -30.290 91.180 ;
        RECT -26.410 90.050 -26.220 91.180 ;
        RECT -20.560 90.050 -20.370 91.180 ;
        RECT -16.490 90.050 -16.300 91.180 ;
        RECT -10.640 90.050 -10.450 91.180 ;
        RECT -6.570 90.050 -6.380 91.180 ;
        RECT -0.720 90.050 -0.530 91.180 ;
        RECT 3.350 90.050 3.540 91.180 ;
        RECT 9.200 90.050 9.390 91.180 ;
        RECT 13.270 90.050 13.460 91.180 ;
        RECT 19.120 90.050 19.310 91.180 ;
        RECT 23.190 90.050 23.380 91.180 ;
        RECT -288.450 89.760 -288.130 90.050 ;
        RECT -284.410 89.760 -284.090 90.050 ;
        RECT -278.530 89.760 -278.210 90.050 ;
        RECT -274.490 89.760 -274.170 90.050 ;
        RECT -268.610 89.760 -268.290 90.050 ;
        RECT -264.570 89.760 -264.250 90.050 ;
        RECT -258.690 89.760 -258.370 90.050 ;
        RECT -254.650 89.760 -254.330 90.050 ;
        RECT -248.770 89.760 -248.450 90.050 ;
        RECT -244.730 89.760 -244.410 90.050 ;
        RECT -238.850 89.760 -238.530 90.050 ;
        RECT -234.810 89.760 -234.490 90.050 ;
        RECT -228.930 89.760 -228.610 90.050 ;
        RECT -224.890 89.760 -224.570 90.050 ;
        RECT -219.010 89.760 -218.690 90.050 ;
        RECT -214.970 89.760 -214.650 90.050 ;
        RECT -209.090 89.760 -208.770 90.050 ;
        RECT -205.050 89.760 -204.730 90.050 ;
        RECT -199.170 89.760 -198.850 90.050 ;
        RECT -195.130 89.760 -194.810 90.050 ;
        RECT -189.250 89.760 -188.930 90.050 ;
        RECT -185.210 89.760 -184.890 90.050 ;
        RECT -179.330 89.760 -179.010 90.050 ;
        RECT -175.290 89.760 -174.970 90.050 ;
        RECT -169.410 89.760 -169.090 90.050 ;
        RECT -165.370 89.760 -165.050 90.050 ;
        RECT -159.490 89.760 -159.170 90.050 ;
        RECT -155.450 89.760 -155.130 90.050 ;
        RECT -149.570 89.760 -149.250 90.050 ;
        RECT -145.530 89.760 -145.210 90.050 ;
        RECT -139.650 89.760 -139.330 90.050 ;
        RECT -135.610 89.760 -135.290 90.050 ;
        RECT -129.730 89.760 -129.410 90.050 ;
        RECT -125.690 89.760 -125.370 90.050 ;
        RECT -119.810 89.760 -119.490 90.050 ;
        RECT -115.770 89.760 -115.450 90.050 ;
        RECT -109.890 89.760 -109.570 90.050 ;
        RECT -105.850 89.760 -105.530 90.050 ;
        RECT -99.970 89.760 -99.650 90.050 ;
        RECT -95.930 89.760 -95.610 90.050 ;
        RECT -90.050 89.760 -89.730 90.050 ;
        RECT -86.010 89.760 -85.690 90.050 ;
        RECT -80.130 89.760 -79.810 90.050 ;
        RECT -76.090 89.760 -75.770 90.050 ;
        RECT -70.210 89.760 -69.890 90.050 ;
        RECT -66.170 89.760 -65.850 90.050 ;
        RECT -60.290 89.760 -59.970 90.050 ;
        RECT -56.250 89.760 -55.930 90.050 ;
        RECT -50.370 89.760 -50.050 90.050 ;
        RECT -46.330 89.760 -46.010 90.050 ;
        RECT -40.450 89.760 -40.130 90.050 ;
        RECT -36.410 89.760 -36.090 90.050 ;
        RECT -30.530 89.760 -30.210 90.050 ;
        RECT -26.490 89.760 -26.170 90.050 ;
        RECT -20.610 89.760 -20.290 90.050 ;
        RECT -16.570 89.760 -16.250 90.050 ;
        RECT -10.690 89.760 -10.370 90.050 ;
        RECT -6.650 89.760 -6.330 90.050 ;
        RECT -0.770 89.760 -0.450 90.050 ;
        RECT 3.270 89.760 3.590 90.050 ;
        RECT 9.150 89.760 9.470 90.050 ;
        RECT 13.190 89.760 13.510 90.050 ;
        RECT 19.070 89.760 19.390 90.050 ;
        RECT 23.110 89.760 23.430 90.050 ;
        RECT -290.160 88.800 -289.220 89.280 ;
        RECT 24.200 89.280 24.680 90.180 ;
        RECT -285.150 88.880 -283.460 89.180 ;
        RECT -275.230 88.880 -273.540 89.180 ;
        RECT -265.310 88.880 -263.620 89.180 ;
        RECT -255.390 88.880 -253.700 89.180 ;
        RECT -245.470 88.880 -243.780 89.180 ;
        RECT -235.550 88.880 -233.860 89.180 ;
        RECT -225.630 88.880 -223.940 89.180 ;
        RECT -215.710 88.880 -214.020 89.180 ;
        RECT -205.790 88.880 -204.100 89.180 ;
        RECT -195.870 88.880 -194.180 89.180 ;
        RECT -185.950 88.880 -184.260 89.180 ;
        RECT -176.030 88.880 -174.340 89.180 ;
        RECT -166.110 88.880 -164.420 89.180 ;
        RECT -156.190 88.880 -154.500 89.180 ;
        RECT -146.270 88.880 -144.580 89.180 ;
        RECT -136.350 88.880 -134.660 89.180 ;
        RECT -126.430 88.880 -124.740 89.180 ;
        RECT -116.510 88.880 -114.820 89.180 ;
        RECT -106.590 88.880 -104.900 89.180 ;
        RECT -96.670 88.880 -94.980 89.180 ;
        RECT -86.750 88.880 -85.060 89.180 ;
        RECT -76.830 88.880 -75.140 89.180 ;
        RECT -66.910 88.880 -65.220 89.180 ;
        RECT -56.990 88.880 -55.300 89.180 ;
        RECT -47.070 88.880 -45.380 89.180 ;
        RECT -37.150 88.880 -35.460 89.180 ;
        RECT -27.230 88.880 -25.540 89.180 ;
        RECT -17.310 88.880 -15.620 89.180 ;
        RECT -7.390 88.880 -5.700 89.180 ;
        RECT 2.530 88.880 4.220 89.180 ;
        RECT 12.450 88.880 14.140 89.180 ;
        RECT 22.370 88.880 24.060 89.180 ;
        RECT -284.640 88.180 -283.640 88.880 ;
        RECT -274.720 88.180 -273.720 88.880 ;
        RECT -264.800 88.180 -263.800 88.880 ;
        RECT -254.880 88.180 -253.880 88.880 ;
        RECT -244.960 88.180 -243.960 88.880 ;
        RECT -235.040 88.180 -234.040 88.880 ;
        RECT -225.120 88.180 -224.120 88.880 ;
        RECT -215.200 88.180 -214.200 88.880 ;
        RECT -205.280 88.180 -204.280 88.880 ;
        RECT -195.360 88.180 -194.360 88.880 ;
        RECT -185.440 88.180 -184.440 88.880 ;
        RECT -175.520 88.180 -174.520 88.880 ;
        RECT -165.600 88.180 -164.600 88.880 ;
        RECT -155.680 88.180 -154.680 88.880 ;
        RECT -145.760 88.180 -144.760 88.880 ;
        RECT -135.840 88.180 -134.840 88.880 ;
        RECT -125.920 88.180 -124.920 88.880 ;
        RECT -116.000 88.180 -115.000 88.880 ;
        RECT -106.080 88.180 -105.080 88.880 ;
        RECT -96.160 88.180 -95.160 88.880 ;
        RECT -86.240 88.180 -85.240 88.880 ;
        RECT -76.320 88.180 -75.320 88.880 ;
        RECT -66.400 88.180 -65.400 88.880 ;
        RECT -56.480 88.180 -55.480 88.880 ;
        RECT -46.560 88.180 -45.560 88.880 ;
        RECT -36.640 88.180 -35.640 88.880 ;
        RECT -26.720 88.180 -25.720 88.880 ;
        RECT -16.800 88.180 -15.800 88.880 ;
        RECT -6.880 88.180 -5.880 88.880 ;
        RECT 3.040 88.180 4.040 88.880 ;
        RECT 12.960 88.180 13.960 88.880 ;
        RECT 22.880 88.180 23.880 88.880 ;
        RECT 24.200 88.800 25.140 89.280 ;
  END
END meta_srlatch_array_row
END LIBRARY

