VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO meta_srlatch_set
  CLASS BLOCK ;
  FOREIGN meta_srlatch_set ;
  ORIGIN 367.230 196.620 ;
  SIZE 533.840 BY 306.490 ;
  SITE unithd ;
  PIN o_ranQ[1]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 18.315 89.065 18.820 89.145 ;
        RECT 19.620 89.065 20.525 89.155 ;
        RECT 18.315 88.885 20.525 89.065 ;
      LAYER mcon ;
        RECT 18.505 88.975 18.675 89.145 ;
        RECT 19.870 88.975 20.040 89.145 ;
      LAYER met1 ;
        RECT 18.440 88.880 20.130 89.180 ;
        RECT 18.620 88.180 19.620 88.880 ;
    END
  END o_ranQ[1]
  PIN o_ranQ[2]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 13.355 94.875 15.565 95.055 ;
        RECT 13.355 94.795 13.860 94.875 ;
        RECT 14.660 94.785 15.565 94.875 ;
      LAYER mcon ;
        RECT 13.545 94.795 13.715 94.965 ;
        RECT 14.910 94.795 15.080 94.965 ;
      LAYER met1 ;
        RECT 13.660 95.060 14.660 95.760 ;
        RECT 13.480 94.760 15.170 95.060 ;
    END
  END o_ranQ[2]
  PIN o_ranQ[3]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 8.395 89.065 8.900 89.145 ;
        RECT 9.700 89.065 10.605 89.155 ;
        RECT 8.395 88.885 10.605 89.065 ;
      LAYER mcon ;
        RECT 8.585 88.975 8.755 89.145 ;
        RECT 9.950 88.975 10.120 89.145 ;
      LAYER met1 ;
        RECT 8.520 88.880 10.210 89.180 ;
        RECT 8.700 88.180 9.700 88.880 ;
    END
  END o_ranQ[3]
  PIN o_ranQ[0]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 23.275 94.875 25.485 95.055 ;
        RECT 23.275 94.795 23.780 94.875 ;
        RECT 24.580 94.785 25.485 94.875 ;
      LAYER mcon ;
        RECT 23.465 94.795 23.635 94.965 ;
        RECT 24.830 94.795 25.000 94.965 ;
      LAYER met1 ;
        RECT 23.580 95.060 24.580 95.760 ;
        RECT 23.400 94.760 25.090 95.060 ;
    END
  END o_ranQ[0]
  PIN o_ranQ[4]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 3.435 94.875 5.645 95.055 ;
        RECT 3.435 94.795 3.940 94.875 ;
        RECT 4.740 94.785 5.645 94.875 ;
      LAYER mcon ;
        RECT 3.625 94.795 3.795 94.965 ;
        RECT 4.990 94.795 5.160 94.965 ;
      LAYER met1 ;
        RECT 3.740 95.060 4.740 95.760 ;
        RECT 3.560 94.760 5.250 95.060 ;
    END
  END o_ranQ[4]
  PIN o_ranQ[5]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -1.525 89.065 -1.020 89.145 ;
        RECT -0.220 89.065 0.685 89.155 ;
        RECT -1.525 88.885 0.685 89.065 ;
      LAYER mcon ;
        RECT -1.335 88.975 -1.165 89.145 ;
        RECT 0.030 88.975 0.200 89.145 ;
      LAYER met1 ;
        RECT -1.400 88.880 0.290 89.180 ;
        RECT -1.220 88.180 -0.220 88.880 ;
    END
  END o_ranQ[5]
  PIN o_ranQ[6]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -6.485 94.875 -4.275 95.055 ;
        RECT -6.485 94.795 -5.980 94.875 ;
        RECT -5.180 94.785 -4.275 94.875 ;
      LAYER mcon ;
        RECT -6.295 94.795 -6.125 94.965 ;
        RECT -4.930 94.795 -4.760 94.965 ;
      LAYER met1 ;
        RECT -6.180 95.060 -5.180 95.760 ;
        RECT -6.360 94.760 -4.670 95.060 ;
    END
  END o_ranQ[6]
  PIN o_ranQ[7]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -11.445 89.065 -10.940 89.145 ;
        RECT -10.140 89.065 -9.235 89.155 ;
        RECT -11.445 88.885 -9.235 89.065 ;
      LAYER mcon ;
        RECT -11.255 88.975 -11.085 89.145 ;
        RECT -9.890 88.975 -9.720 89.145 ;
      LAYER met1 ;
        RECT -11.320 88.880 -9.630 89.180 ;
        RECT -11.140 88.180 -10.140 88.880 ;
    END
  END o_ranQ[7]
  PIN o_ranQ[8]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -16.405 94.875 -14.195 95.055 ;
        RECT -16.405 94.795 -15.900 94.875 ;
        RECT -15.100 94.785 -14.195 94.875 ;
      LAYER mcon ;
        RECT -16.215 94.795 -16.045 94.965 ;
        RECT -14.850 94.795 -14.680 94.965 ;
      LAYER met1 ;
        RECT -16.100 95.060 -15.100 95.760 ;
        RECT -16.280 94.760 -14.590 95.060 ;
    END
  END o_ranQ[8]
  PIN o_ranQ[9]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -21.365 89.065 -20.860 89.145 ;
        RECT -20.060 89.065 -19.155 89.155 ;
        RECT -21.365 88.885 -19.155 89.065 ;
      LAYER mcon ;
        RECT -21.175 88.975 -21.005 89.145 ;
        RECT -19.810 88.975 -19.640 89.145 ;
      LAYER met1 ;
        RECT -21.240 88.880 -19.550 89.180 ;
        RECT -21.060 88.180 -20.060 88.880 ;
    END
  END o_ranQ[9]
  PIN o_ranQ[10]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -26.325 94.875 -24.115 95.055 ;
        RECT -26.325 94.795 -25.820 94.875 ;
        RECT -25.020 94.785 -24.115 94.875 ;
      LAYER mcon ;
        RECT -26.135 94.795 -25.965 94.965 ;
        RECT -24.770 94.795 -24.600 94.965 ;
      LAYER met1 ;
        RECT -26.020 95.060 -25.020 95.760 ;
        RECT -26.200 94.760 -24.510 95.060 ;
    END
  END o_ranQ[10]
  PIN o_ranQ[11]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -31.285 89.065 -30.780 89.145 ;
        RECT -29.980 89.065 -29.075 89.155 ;
        RECT -31.285 88.885 -29.075 89.065 ;
      LAYER mcon ;
        RECT -31.095 88.975 -30.925 89.145 ;
        RECT -29.730 88.975 -29.560 89.145 ;
      LAYER met1 ;
        RECT -31.160 88.880 -29.470 89.180 ;
        RECT -30.980 88.180 -29.980 88.880 ;
    END
  END o_ranQ[11]
  PIN o_ranQ[12]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -36.245 94.875 -34.035 95.055 ;
        RECT -36.245 94.795 -35.740 94.875 ;
        RECT -34.940 94.785 -34.035 94.875 ;
      LAYER mcon ;
        RECT -36.055 94.795 -35.885 94.965 ;
        RECT -34.690 94.795 -34.520 94.965 ;
      LAYER met1 ;
        RECT -35.940 95.060 -34.940 95.760 ;
        RECT -36.120 94.760 -34.430 95.060 ;
    END
  END o_ranQ[12]
  PIN o_ranQ[13]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -41.205 89.065 -40.700 89.145 ;
        RECT -39.900 89.065 -38.995 89.155 ;
        RECT -41.205 88.885 -38.995 89.065 ;
      LAYER mcon ;
        RECT -41.015 88.975 -40.845 89.145 ;
        RECT -39.650 88.975 -39.480 89.145 ;
      LAYER met1 ;
        RECT -41.080 88.880 -39.390 89.180 ;
        RECT -40.900 88.180 -39.900 88.880 ;
    END
  END o_ranQ[13]
  PIN o_ranQ[14]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -46.165 94.875 -43.955 95.055 ;
        RECT -46.165 94.795 -45.660 94.875 ;
        RECT -44.860 94.785 -43.955 94.875 ;
      LAYER mcon ;
        RECT -45.975 94.795 -45.805 94.965 ;
        RECT -44.610 94.795 -44.440 94.965 ;
      LAYER met1 ;
        RECT -45.860 95.060 -44.860 95.760 ;
        RECT -46.040 94.760 -44.350 95.060 ;
    END
  END o_ranQ[14]
  PIN o_ranQ[15]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -51.125 89.065 -50.620 89.145 ;
        RECT -49.820 89.065 -48.915 89.155 ;
        RECT -51.125 88.885 -48.915 89.065 ;
      LAYER mcon ;
        RECT -50.935 88.975 -50.765 89.145 ;
        RECT -49.570 88.975 -49.400 89.145 ;
      LAYER met1 ;
        RECT -51.000 88.880 -49.310 89.180 ;
        RECT -50.820 88.180 -49.820 88.880 ;
    END
  END o_ranQ[15]
  PIN o_ranQ[17]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -61.045 89.065 -60.540 89.145 ;
        RECT -59.740 89.065 -58.835 89.155 ;
        RECT -61.045 88.885 -58.835 89.065 ;
      LAYER mcon ;
        RECT -60.855 88.975 -60.685 89.145 ;
        RECT -59.490 88.975 -59.320 89.145 ;
      LAYER met1 ;
        RECT -60.920 88.880 -59.230 89.180 ;
        RECT -60.740 88.180 -59.740 88.880 ;
    END
  END o_ranQ[17]
  PIN o_ranQ[18]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -66.005 94.875 -63.795 95.055 ;
        RECT -66.005 94.795 -65.500 94.875 ;
        RECT -64.700 94.785 -63.795 94.875 ;
      LAYER mcon ;
        RECT -65.815 94.795 -65.645 94.965 ;
        RECT -64.450 94.795 -64.280 94.965 ;
      LAYER met1 ;
        RECT -65.700 95.060 -64.700 95.760 ;
        RECT -65.880 94.760 -64.190 95.060 ;
    END
  END o_ranQ[18]
  PIN o_ranQ[19]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -70.965 89.065 -70.460 89.145 ;
        RECT -69.660 89.065 -68.755 89.155 ;
        RECT -70.965 88.885 -68.755 89.065 ;
      LAYER mcon ;
        RECT -70.775 88.975 -70.605 89.145 ;
        RECT -69.410 88.975 -69.240 89.145 ;
      LAYER met1 ;
        RECT -70.840 88.880 -69.150 89.180 ;
        RECT -70.660 88.180 -69.660 88.880 ;
    END
  END o_ranQ[19]
  PIN o_ranQ[16]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -56.085 94.875 -53.875 95.055 ;
        RECT -56.085 94.795 -55.580 94.875 ;
        RECT -54.780 94.785 -53.875 94.875 ;
      LAYER mcon ;
        RECT -55.895 94.795 -55.725 94.965 ;
        RECT -54.530 94.795 -54.360 94.965 ;
      LAYER met1 ;
        RECT -55.780 95.060 -54.780 95.760 ;
        RECT -55.960 94.760 -54.270 95.060 ;
    END
  END o_ranQ[16]
  PIN o_ranQ[20]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -75.925 94.875 -73.715 95.055 ;
        RECT -75.925 94.795 -75.420 94.875 ;
        RECT -74.620 94.785 -73.715 94.875 ;
      LAYER mcon ;
        RECT -75.735 94.795 -75.565 94.965 ;
        RECT -74.370 94.795 -74.200 94.965 ;
      LAYER met1 ;
        RECT -75.620 95.060 -74.620 95.760 ;
        RECT -75.800 94.760 -74.110 95.060 ;
    END
  END o_ranQ[20]
  PIN o_ranQ[21]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -80.885 89.065 -80.380 89.145 ;
        RECT -79.580 89.065 -78.675 89.155 ;
        RECT -80.885 88.885 -78.675 89.065 ;
      LAYER mcon ;
        RECT -80.695 88.975 -80.525 89.145 ;
        RECT -79.330 88.975 -79.160 89.145 ;
      LAYER met1 ;
        RECT -80.760 88.880 -79.070 89.180 ;
        RECT -80.580 88.180 -79.580 88.880 ;
    END
  END o_ranQ[21]
  PIN o_ranQ[22]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -85.845 94.875 -83.635 95.055 ;
        RECT -85.845 94.795 -85.340 94.875 ;
        RECT -84.540 94.785 -83.635 94.875 ;
      LAYER mcon ;
        RECT -85.655 94.795 -85.485 94.965 ;
        RECT -84.290 94.795 -84.120 94.965 ;
      LAYER met1 ;
        RECT -85.540 95.060 -84.540 95.760 ;
        RECT -85.720 94.760 -84.030 95.060 ;
    END
  END o_ranQ[22]
  PIN o_ranQ[23]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -90.805 89.065 -90.300 89.145 ;
        RECT -89.500 89.065 -88.595 89.155 ;
        RECT -90.805 88.885 -88.595 89.065 ;
      LAYER mcon ;
        RECT -90.615 88.975 -90.445 89.145 ;
        RECT -89.250 88.975 -89.080 89.145 ;
      LAYER met1 ;
        RECT -90.680 88.880 -88.990 89.180 ;
        RECT -90.500 88.180 -89.500 88.880 ;
    END
  END o_ranQ[23]
  PIN o_ranQ[24]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -95.765 94.875 -93.555 95.055 ;
        RECT -95.765 94.795 -95.260 94.875 ;
        RECT -94.460 94.785 -93.555 94.875 ;
      LAYER mcon ;
        RECT -95.575 94.795 -95.405 94.965 ;
        RECT -94.210 94.795 -94.040 94.965 ;
      LAYER met1 ;
        RECT -95.460 95.060 -94.460 95.760 ;
        RECT -95.640 94.760 -93.950 95.060 ;
    END
  END o_ranQ[24]
  PIN o_ranQ[25]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -100.725 89.065 -100.220 89.145 ;
        RECT -99.420 89.065 -98.515 89.155 ;
        RECT -100.725 88.885 -98.515 89.065 ;
      LAYER mcon ;
        RECT -100.535 88.975 -100.365 89.145 ;
        RECT -99.170 88.975 -99.000 89.145 ;
      LAYER met1 ;
        RECT -100.600 88.880 -98.910 89.180 ;
        RECT -100.420 88.180 -99.420 88.880 ;
    END
  END o_ranQ[25]
  PIN o_ranQ[26]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -105.685 94.875 -103.475 95.055 ;
        RECT -105.685 94.795 -105.180 94.875 ;
        RECT -104.380 94.785 -103.475 94.875 ;
      LAYER mcon ;
        RECT -105.495 94.795 -105.325 94.965 ;
        RECT -104.130 94.795 -103.960 94.965 ;
      LAYER met1 ;
        RECT -105.380 95.060 -104.380 95.760 ;
        RECT -105.560 94.760 -103.870 95.060 ;
    END
  END o_ranQ[26]
  PIN o_ranQ[27]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -110.645 89.065 -110.140 89.145 ;
        RECT -109.340 89.065 -108.435 89.155 ;
        RECT -110.645 88.885 -108.435 89.065 ;
      LAYER mcon ;
        RECT -110.455 88.975 -110.285 89.145 ;
        RECT -109.090 88.975 -108.920 89.145 ;
      LAYER met1 ;
        RECT -110.520 88.880 -108.830 89.180 ;
        RECT -110.340 88.180 -109.340 88.880 ;
    END
  END o_ranQ[27]
  PIN o_ranQ[28]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -115.605 94.875 -113.395 95.055 ;
        RECT -115.605 94.795 -115.100 94.875 ;
        RECT -114.300 94.785 -113.395 94.875 ;
      LAYER mcon ;
        RECT -115.415 94.795 -115.245 94.965 ;
        RECT -114.050 94.795 -113.880 94.965 ;
      LAYER met1 ;
        RECT -115.300 95.060 -114.300 95.760 ;
        RECT -115.480 94.760 -113.790 95.060 ;
    END
  END o_ranQ[28]
  PIN o_ranQ[29]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -120.565 89.065 -120.060 89.145 ;
        RECT -119.260 89.065 -118.355 89.155 ;
        RECT -120.565 88.885 -118.355 89.065 ;
      LAYER mcon ;
        RECT -120.375 88.975 -120.205 89.145 ;
        RECT -119.010 88.975 -118.840 89.145 ;
      LAYER met1 ;
        RECT -120.440 88.880 -118.750 89.180 ;
        RECT -120.260 88.180 -119.260 88.880 ;
    END
  END o_ranQ[29]
  PIN o_ranQ[30]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -125.525 94.875 -123.315 95.055 ;
        RECT -125.525 94.795 -125.020 94.875 ;
        RECT -124.220 94.785 -123.315 94.875 ;
      LAYER mcon ;
        RECT -125.335 94.795 -125.165 94.965 ;
        RECT -123.970 94.795 -123.800 94.965 ;
      LAYER met1 ;
        RECT -125.220 95.060 -124.220 95.760 ;
        RECT -125.400 94.760 -123.710 95.060 ;
    END
  END o_ranQ[30]
  PIN o_ranQ[31]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -130.485 89.065 -129.980 89.145 ;
        RECT -129.180 89.065 -128.275 89.155 ;
        RECT -130.485 88.885 -128.275 89.065 ;
      LAYER mcon ;
        RECT -130.295 88.975 -130.125 89.145 ;
        RECT -128.930 88.975 -128.760 89.145 ;
      LAYER met1 ;
        RECT -130.360 88.880 -128.670 89.180 ;
        RECT -130.180 88.180 -129.180 88.880 ;
    END
  END o_ranQ[31]
  PIN o_ranQ[33]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -140.405 89.065 -139.900 89.145 ;
        RECT -139.100 89.065 -138.195 89.155 ;
        RECT -140.405 88.885 -138.195 89.065 ;
      LAYER mcon ;
        RECT -140.215 88.975 -140.045 89.145 ;
        RECT -138.850 88.975 -138.680 89.145 ;
      LAYER met1 ;
        RECT -140.280 88.880 -138.590 89.180 ;
        RECT -140.100 88.180 -139.100 88.880 ;
    END
  END o_ranQ[33]
  PIN o_ranQ[34]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -145.365 94.875 -143.155 95.055 ;
        RECT -145.365 94.795 -144.860 94.875 ;
        RECT -144.060 94.785 -143.155 94.875 ;
      LAYER mcon ;
        RECT -145.175 94.795 -145.005 94.965 ;
        RECT -143.810 94.795 -143.640 94.965 ;
      LAYER met1 ;
        RECT -145.060 95.060 -144.060 95.760 ;
        RECT -145.240 94.760 -143.550 95.060 ;
    END
  END o_ranQ[34]
  PIN o_ranQ[35]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -150.325 89.065 -149.820 89.145 ;
        RECT -149.020 89.065 -148.115 89.155 ;
        RECT -150.325 88.885 -148.115 89.065 ;
      LAYER mcon ;
        RECT -150.135 88.975 -149.965 89.145 ;
        RECT -148.770 88.975 -148.600 89.145 ;
      LAYER met1 ;
        RECT -150.200 88.880 -148.510 89.180 ;
        RECT -150.020 88.180 -149.020 88.880 ;
    END
  END o_ranQ[35]
  PIN o_ranQ[32]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -135.445 94.875 -133.235 95.055 ;
        RECT -135.445 94.795 -134.940 94.875 ;
        RECT -134.140 94.785 -133.235 94.875 ;
      LAYER mcon ;
        RECT -135.255 94.795 -135.085 94.965 ;
        RECT -133.890 94.795 -133.720 94.965 ;
      LAYER met1 ;
        RECT -135.140 95.060 -134.140 95.760 ;
        RECT -135.320 94.760 -133.630 95.060 ;
    END
  END o_ranQ[32]
  PIN o_ranQ[36]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -155.285 94.875 -153.075 95.055 ;
        RECT -155.285 94.795 -154.780 94.875 ;
        RECT -153.980 94.785 -153.075 94.875 ;
      LAYER mcon ;
        RECT -155.095 94.795 -154.925 94.965 ;
        RECT -153.730 94.795 -153.560 94.965 ;
      LAYER met1 ;
        RECT -154.980 95.060 -153.980 95.760 ;
        RECT -155.160 94.760 -153.470 95.060 ;
    END
  END o_ranQ[36]
  PIN o_ranQ[37]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -160.245 89.065 -159.740 89.145 ;
        RECT -158.940 89.065 -158.035 89.155 ;
        RECT -160.245 88.885 -158.035 89.065 ;
      LAYER mcon ;
        RECT -160.055 88.975 -159.885 89.145 ;
        RECT -158.690 88.975 -158.520 89.145 ;
      LAYER met1 ;
        RECT -160.120 88.880 -158.430 89.180 ;
        RECT -159.940 88.180 -158.940 88.880 ;
    END
  END o_ranQ[37]
  PIN o_ranQ[38]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -165.205 94.875 -162.995 95.055 ;
        RECT -165.205 94.795 -164.700 94.875 ;
        RECT -163.900 94.785 -162.995 94.875 ;
      LAYER mcon ;
        RECT -165.015 94.795 -164.845 94.965 ;
        RECT -163.650 94.795 -163.480 94.965 ;
      LAYER met1 ;
        RECT -164.900 95.060 -163.900 95.760 ;
        RECT -165.080 94.760 -163.390 95.060 ;
    END
  END o_ranQ[38]
  PIN o_ranQ[39]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -170.165 89.065 -169.660 89.145 ;
        RECT -168.860 89.065 -167.955 89.155 ;
        RECT -170.165 88.885 -167.955 89.065 ;
      LAYER mcon ;
        RECT -169.975 88.975 -169.805 89.145 ;
        RECT -168.610 88.975 -168.440 89.145 ;
      LAYER met1 ;
        RECT -170.040 88.880 -168.350 89.180 ;
        RECT -169.860 88.180 -168.860 88.880 ;
    END
  END o_ranQ[39]
  PIN o_ranQ[40]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -175.125 94.875 -172.915 95.055 ;
        RECT -175.125 94.795 -174.620 94.875 ;
        RECT -173.820 94.785 -172.915 94.875 ;
      LAYER mcon ;
        RECT -174.935 94.795 -174.765 94.965 ;
        RECT -173.570 94.795 -173.400 94.965 ;
      LAYER met1 ;
        RECT -174.820 95.060 -173.820 95.760 ;
        RECT -175.000 94.760 -173.310 95.060 ;
    END
  END o_ranQ[40]
  PIN o_ranQ[41]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -180.085 89.065 -179.580 89.145 ;
        RECT -178.780 89.065 -177.875 89.155 ;
        RECT -180.085 88.885 -177.875 89.065 ;
      LAYER mcon ;
        RECT -179.895 88.975 -179.725 89.145 ;
        RECT -178.530 88.975 -178.360 89.145 ;
      LAYER met1 ;
        RECT -179.960 88.880 -178.270 89.180 ;
        RECT -179.780 88.180 -178.780 88.880 ;
    END
  END o_ranQ[41]
  PIN o_ranQ[42]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -185.045 94.875 -182.835 95.055 ;
        RECT -185.045 94.795 -184.540 94.875 ;
        RECT -183.740 94.785 -182.835 94.875 ;
      LAYER mcon ;
        RECT -184.855 94.795 -184.685 94.965 ;
        RECT -183.490 94.795 -183.320 94.965 ;
      LAYER met1 ;
        RECT -184.740 95.060 -183.740 95.760 ;
        RECT -184.920 94.760 -183.230 95.060 ;
    END
  END o_ranQ[42]
  PIN o_ranQ[43]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -190.005 89.065 -189.500 89.145 ;
        RECT -188.700 89.065 -187.795 89.155 ;
        RECT -190.005 88.885 -187.795 89.065 ;
      LAYER mcon ;
        RECT -189.815 88.975 -189.645 89.145 ;
        RECT -188.450 88.975 -188.280 89.145 ;
      LAYER met1 ;
        RECT -189.880 88.880 -188.190 89.180 ;
        RECT -189.700 88.180 -188.700 88.880 ;
    END
  END o_ranQ[43]
  PIN o_ranQ[44]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -194.965 94.875 -192.755 95.055 ;
        RECT -194.965 94.795 -194.460 94.875 ;
        RECT -193.660 94.785 -192.755 94.875 ;
      LAYER mcon ;
        RECT -194.775 94.795 -194.605 94.965 ;
        RECT -193.410 94.795 -193.240 94.965 ;
      LAYER met1 ;
        RECT -194.660 95.060 -193.660 95.760 ;
        RECT -194.840 94.760 -193.150 95.060 ;
    END
  END o_ranQ[44]
  PIN o_ranQ[45]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -199.925 89.065 -199.420 89.145 ;
        RECT -198.620 89.065 -197.715 89.155 ;
        RECT -199.925 88.885 -197.715 89.065 ;
      LAYER mcon ;
        RECT -199.735 88.975 -199.565 89.145 ;
        RECT -198.370 88.975 -198.200 89.145 ;
      LAYER met1 ;
        RECT -199.800 88.880 -198.110 89.180 ;
        RECT -199.620 88.180 -198.620 88.880 ;
    END
  END o_ranQ[45]
  PIN o_ranQ[46]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -204.885 94.875 -202.675 95.055 ;
        RECT -204.885 94.795 -204.380 94.875 ;
        RECT -203.580 94.785 -202.675 94.875 ;
      LAYER mcon ;
        RECT -204.695 94.795 -204.525 94.965 ;
        RECT -203.330 94.795 -203.160 94.965 ;
      LAYER met1 ;
        RECT -204.580 95.060 -203.580 95.760 ;
        RECT -204.760 94.760 -203.070 95.060 ;
    END
  END o_ranQ[46]
  PIN o_ranQ[47]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -209.845 89.065 -209.340 89.145 ;
        RECT -208.540 89.065 -207.635 89.155 ;
        RECT -209.845 88.885 -207.635 89.065 ;
      LAYER mcon ;
        RECT -209.655 88.975 -209.485 89.145 ;
        RECT -208.290 88.975 -208.120 89.145 ;
      LAYER met1 ;
        RECT -209.720 88.880 -208.030 89.180 ;
        RECT -209.540 88.180 -208.540 88.880 ;
    END
  END o_ranQ[47]
  PIN o_ranQ[49]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -219.765 89.065 -219.260 89.145 ;
        RECT -218.460 89.065 -217.555 89.155 ;
        RECT -219.765 88.885 -217.555 89.065 ;
      LAYER mcon ;
        RECT -219.575 88.975 -219.405 89.145 ;
        RECT -218.210 88.975 -218.040 89.145 ;
      LAYER met1 ;
        RECT -219.640 88.880 -217.950 89.180 ;
        RECT -219.460 88.180 -218.460 88.880 ;
    END
  END o_ranQ[49]
  PIN o_ranQ[50]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -224.725 94.875 -222.515 95.055 ;
        RECT -224.725 94.795 -224.220 94.875 ;
        RECT -223.420 94.785 -222.515 94.875 ;
      LAYER mcon ;
        RECT -224.535 94.795 -224.365 94.965 ;
        RECT -223.170 94.795 -223.000 94.965 ;
      LAYER met1 ;
        RECT -224.420 95.060 -223.420 95.760 ;
        RECT -224.600 94.760 -222.910 95.060 ;
    END
  END o_ranQ[50]
  PIN o_ranQ[51]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -229.685 89.065 -229.180 89.145 ;
        RECT -228.380 89.065 -227.475 89.155 ;
        RECT -229.685 88.885 -227.475 89.065 ;
      LAYER mcon ;
        RECT -229.495 88.975 -229.325 89.145 ;
        RECT -228.130 88.975 -227.960 89.145 ;
      LAYER met1 ;
        RECT -229.560 88.880 -227.870 89.180 ;
        RECT -229.380 88.180 -228.380 88.880 ;
    END
  END o_ranQ[51]
  PIN o_ranQ[48]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -214.805 94.875 -212.595 95.055 ;
        RECT -214.805 94.795 -214.300 94.875 ;
        RECT -213.500 94.785 -212.595 94.875 ;
      LAYER mcon ;
        RECT -214.615 94.795 -214.445 94.965 ;
        RECT -213.250 94.795 -213.080 94.965 ;
      LAYER met1 ;
        RECT -214.500 95.060 -213.500 95.760 ;
        RECT -214.680 94.760 -212.990 95.060 ;
    END
  END o_ranQ[48]
  PIN o_ranQ[52]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -234.645 94.875 -232.435 95.055 ;
        RECT -234.645 94.795 -234.140 94.875 ;
        RECT -233.340 94.785 -232.435 94.875 ;
      LAYER mcon ;
        RECT -234.455 94.795 -234.285 94.965 ;
        RECT -233.090 94.795 -232.920 94.965 ;
      LAYER met1 ;
        RECT -234.340 95.060 -233.340 95.760 ;
        RECT -234.520 94.760 -232.830 95.060 ;
    END
  END o_ranQ[52]
  PIN o_ranQ[53]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -239.605 89.065 -239.100 89.145 ;
        RECT -238.300 89.065 -237.395 89.155 ;
        RECT -239.605 88.885 -237.395 89.065 ;
      LAYER mcon ;
        RECT -239.415 88.975 -239.245 89.145 ;
        RECT -238.050 88.975 -237.880 89.145 ;
      LAYER met1 ;
        RECT -239.480 88.880 -237.790 89.180 ;
        RECT -239.300 88.180 -238.300 88.880 ;
    END
  END o_ranQ[53]
  PIN o_ranQ[54]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -244.565 94.875 -242.355 95.055 ;
        RECT -244.565 94.795 -244.060 94.875 ;
        RECT -243.260 94.785 -242.355 94.875 ;
      LAYER mcon ;
        RECT -244.375 94.795 -244.205 94.965 ;
        RECT -243.010 94.795 -242.840 94.965 ;
      LAYER met1 ;
        RECT -244.260 95.060 -243.260 95.760 ;
        RECT -244.440 94.760 -242.750 95.060 ;
    END
  END o_ranQ[54]
  PIN o_ranQ[55]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -249.525 89.065 -249.020 89.145 ;
        RECT -248.220 89.065 -247.315 89.155 ;
        RECT -249.525 88.885 -247.315 89.065 ;
      LAYER mcon ;
        RECT -249.335 88.975 -249.165 89.145 ;
        RECT -247.970 88.975 -247.800 89.145 ;
      LAYER met1 ;
        RECT -249.400 88.880 -247.710 89.180 ;
        RECT -249.220 88.180 -248.220 88.880 ;
    END
  END o_ranQ[55]
  PIN o_ranQ[56]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -254.485 94.875 -252.275 95.055 ;
        RECT -254.485 94.795 -253.980 94.875 ;
        RECT -253.180 94.785 -252.275 94.875 ;
      LAYER mcon ;
        RECT -254.295 94.795 -254.125 94.965 ;
        RECT -252.930 94.795 -252.760 94.965 ;
      LAYER met1 ;
        RECT -254.180 95.060 -253.180 95.760 ;
        RECT -254.360 94.760 -252.670 95.060 ;
    END
  END o_ranQ[56]
  PIN o_ranQ[57]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -259.445 89.065 -258.940 89.145 ;
        RECT -258.140 89.065 -257.235 89.155 ;
        RECT -259.445 88.885 -257.235 89.065 ;
      LAYER mcon ;
        RECT -259.255 88.975 -259.085 89.145 ;
        RECT -257.890 88.975 -257.720 89.145 ;
      LAYER met1 ;
        RECT -259.320 88.880 -257.630 89.180 ;
        RECT -259.140 88.180 -258.140 88.880 ;
    END
  END o_ranQ[57]
  PIN o_ranQ[58]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -264.405 94.875 -262.195 95.055 ;
        RECT -264.405 94.795 -263.900 94.875 ;
        RECT -263.100 94.785 -262.195 94.875 ;
      LAYER mcon ;
        RECT -264.215 94.795 -264.045 94.965 ;
        RECT -262.850 94.795 -262.680 94.965 ;
      LAYER met1 ;
        RECT -264.100 95.060 -263.100 95.760 ;
        RECT -264.280 94.760 -262.590 95.060 ;
    END
  END o_ranQ[58]
  PIN o_ranQ[59]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -269.365 89.065 -268.860 89.145 ;
        RECT -268.060 89.065 -267.155 89.155 ;
        RECT -269.365 88.885 -267.155 89.065 ;
      LAYER mcon ;
        RECT -269.175 88.975 -269.005 89.145 ;
        RECT -267.810 88.975 -267.640 89.145 ;
      LAYER met1 ;
        RECT -269.240 88.880 -267.550 89.180 ;
        RECT -269.060 88.180 -268.060 88.880 ;
    END
  END o_ranQ[59]
  PIN o_ranQ[61]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -279.285 89.065 -278.780 89.145 ;
        RECT -277.980 89.065 -277.075 89.155 ;
        RECT -279.285 88.885 -277.075 89.065 ;
      LAYER mcon ;
        RECT -279.095 88.975 -278.925 89.145 ;
        RECT -277.730 88.975 -277.560 89.145 ;
      LAYER met1 ;
        RECT -279.160 88.880 -277.470 89.180 ;
        RECT -278.980 88.180 -277.980 88.880 ;
    END
  END o_ranQ[61]
  PIN o_ranQ[62]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -284.245 94.875 -282.035 95.055 ;
        RECT -284.245 94.795 -283.740 94.875 ;
        RECT -282.940 94.785 -282.035 94.875 ;
      LAYER mcon ;
        RECT -284.055 94.795 -283.885 94.965 ;
        RECT -282.690 94.795 -282.520 94.965 ;
      LAYER met1 ;
        RECT -283.940 95.060 -282.940 95.760 ;
        RECT -284.120 94.760 -282.430 95.060 ;
    END
  END o_ranQ[62]
  PIN o_ranQ[63]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -289.205 89.065 -288.700 89.145 ;
        RECT -287.900 89.065 -286.995 89.155 ;
        RECT -289.205 88.885 -286.995 89.065 ;
      LAYER mcon ;
        RECT -289.015 88.975 -288.845 89.145 ;
        RECT -287.650 88.975 -287.480 89.145 ;
      LAYER met1 ;
        RECT -289.080 88.880 -287.390 89.180 ;
        RECT -288.900 88.180 -287.900 88.880 ;
    END
  END o_ranQ[63]
  PIN i_srclk
    ANTENNAGATEAREA 126.719994 ;
    PORT
      LAYER li1 ;
        RECT -290.905 92.005 -290.570 92.275 ;
        RECT -281.970 92.005 -281.635 92.275 ;
        RECT -280.985 92.005 -280.650 92.275 ;
        RECT -272.050 92.005 -271.715 92.275 ;
        RECT -271.065 92.005 -270.730 92.275 ;
        RECT -262.130 92.005 -261.795 92.275 ;
        RECT -261.145 92.005 -260.810 92.275 ;
        RECT -252.210 92.005 -251.875 92.275 ;
        RECT -251.225 92.005 -250.890 92.275 ;
        RECT -242.290 92.005 -241.955 92.275 ;
        RECT -241.305 92.005 -240.970 92.275 ;
        RECT -232.370 92.005 -232.035 92.275 ;
        RECT -231.385 92.005 -231.050 92.275 ;
        RECT -222.450 92.005 -222.115 92.275 ;
        RECT -221.465 92.005 -221.130 92.275 ;
        RECT -212.530 92.005 -212.195 92.275 ;
        RECT -211.545 92.005 -211.210 92.275 ;
        RECT -202.610 92.005 -202.275 92.275 ;
        RECT -201.625 92.005 -201.290 92.275 ;
        RECT -192.690 92.005 -192.355 92.275 ;
        RECT -191.705 92.005 -191.370 92.275 ;
        RECT -182.770 92.005 -182.435 92.275 ;
        RECT -181.785 92.005 -181.450 92.275 ;
        RECT -172.850 92.005 -172.515 92.275 ;
        RECT -171.865 92.005 -171.530 92.275 ;
        RECT -162.930 92.005 -162.595 92.275 ;
        RECT -161.945 92.005 -161.610 92.275 ;
        RECT -153.010 92.005 -152.675 92.275 ;
        RECT -152.025 92.005 -151.690 92.275 ;
        RECT -143.090 92.005 -142.755 92.275 ;
        RECT -142.105 92.005 -141.770 92.275 ;
        RECT -133.170 92.005 -132.835 92.275 ;
        RECT -132.185 92.005 -131.850 92.275 ;
        RECT -123.250 92.005 -122.915 92.275 ;
        RECT -122.265 92.005 -121.930 92.275 ;
        RECT -113.330 92.005 -112.995 92.275 ;
        RECT -112.345 92.005 -112.010 92.275 ;
        RECT -103.410 92.005 -103.075 92.275 ;
        RECT -102.425 92.005 -102.090 92.275 ;
        RECT -93.490 92.005 -93.155 92.275 ;
        RECT -92.505 92.005 -92.170 92.275 ;
        RECT -83.570 92.005 -83.235 92.275 ;
        RECT -82.585 92.005 -82.250 92.275 ;
        RECT -73.650 92.005 -73.315 92.275 ;
        RECT -72.665 92.005 -72.330 92.275 ;
        RECT -63.730 92.005 -63.395 92.275 ;
        RECT -62.745 92.005 -62.410 92.275 ;
        RECT -53.810 92.005 -53.475 92.275 ;
        RECT -52.825 92.005 -52.490 92.275 ;
        RECT -43.890 92.005 -43.555 92.275 ;
        RECT -42.905 92.005 -42.570 92.275 ;
        RECT -33.970 92.005 -33.635 92.275 ;
        RECT -32.985 92.005 -32.650 92.275 ;
        RECT -24.050 92.005 -23.715 92.275 ;
        RECT -23.065 92.005 -22.730 92.275 ;
        RECT -14.130 92.005 -13.795 92.275 ;
        RECT -13.145 92.005 -12.810 92.275 ;
        RECT -4.210 92.005 -3.875 92.275 ;
        RECT -3.225 92.005 -2.890 92.275 ;
        RECT 5.710 92.005 6.045 92.275 ;
        RECT 6.695 92.005 7.030 92.275 ;
        RECT 15.630 92.005 15.965 92.275 ;
        RECT 16.615 92.005 16.950 92.275 ;
        RECT 25.550 92.005 25.885 92.275 ;
        RECT -286.930 91.665 -286.595 91.935 ;
        RECT -285.945 91.665 -285.610 91.935 ;
        RECT -277.010 91.665 -276.675 91.935 ;
        RECT -276.025 91.665 -275.690 91.935 ;
        RECT -267.090 91.665 -266.755 91.935 ;
        RECT -266.105 91.665 -265.770 91.935 ;
        RECT -257.170 91.665 -256.835 91.935 ;
        RECT -256.185 91.665 -255.850 91.935 ;
        RECT -247.250 91.665 -246.915 91.935 ;
        RECT -246.265 91.665 -245.930 91.935 ;
        RECT -237.330 91.665 -236.995 91.935 ;
        RECT -236.345 91.665 -236.010 91.935 ;
        RECT -227.410 91.665 -227.075 91.935 ;
        RECT -226.425 91.665 -226.090 91.935 ;
        RECT -217.490 91.665 -217.155 91.935 ;
        RECT -216.505 91.665 -216.170 91.935 ;
        RECT -207.570 91.665 -207.235 91.935 ;
        RECT -206.585 91.665 -206.250 91.935 ;
        RECT -197.650 91.665 -197.315 91.935 ;
        RECT -196.665 91.665 -196.330 91.935 ;
        RECT -187.730 91.665 -187.395 91.935 ;
        RECT -186.745 91.665 -186.410 91.935 ;
        RECT -177.810 91.665 -177.475 91.935 ;
        RECT -176.825 91.665 -176.490 91.935 ;
        RECT -167.890 91.665 -167.555 91.935 ;
        RECT -166.905 91.665 -166.570 91.935 ;
        RECT -157.970 91.665 -157.635 91.935 ;
        RECT -156.985 91.665 -156.650 91.935 ;
        RECT -148.050 91.665 -147.715 91.935 ;
        RECT -147.065 91.665 -146.730 91.935 ;
        RECT -138.130 91.665 -137.795 91.935 ;
        RECT -137.145 91.665 -136.810 91.935 ;
        RECT -128.210 91.665 -127.875 91.935 ;
        RECT -127.225 91.665 -126.890 91.935 ;
        RECT -118.290 91.665 -117.955 91.935 ;
        RECT -117.305 91.665 -116.970 91.935 ;
        RECT -108.370 91.665 -108.035 91.935 ;
        RECT -107.385 91.665 -107.050 91.935 ;
        RECT -98.450 91.665 -98.115 91.935 ;
        RECT -97.465 91.665 -97.130 91.935 ;
        RECT -88.530 91.665 -88.195 91.935 ;
        RECT -87.545 91.665 -87.210 91.935 ;
        RECT -78.610 91.665 -78.275 91.935 ;
        RECT -77.625 91.665 -77.290 91.935 ;
        RECT -68.690 91.665 -68.355 91.935 ;
        RECT -67.705 91.665 -67.370 91.935 ;
        RECT -58.770 91.665 -58.435 91.935 ;
        RECT -57.785 91.665 -57.450 91.935 ;
        RECT -48.850 91.665 -48.515 91.935 ;
        RECT -47.865 91.665 -47.530 91.935 ;
        RECT -38.930 91.665 -38.595 91.935 ;
        RECT -37.945 91.665 -37.610 91.935 ;
        RECT -29.010 91.665 -28.675 91.935 ;
        RECT -28.025 91.665 -27.690 91.935 ;
        RECT -19.090 91.665 -18.755 91.935 ;
        RECT -18.105 91.665 -17.770 91.935 ;
        RECT -9.170 91.665 -8.835 91.935 ;
        RECT -8.185 91.665 -7.850 91.935 ;
        RECT 0.750 91.665 1.085 91.935 ;
        RECT 1.735 91.665 2.070 91.935 ;
        RECT 10.670 91.665 11.005 91.935 ;
        RECT 11.655 91.665 11.990 91.935 ;
        RECT 20.590 91.665 20.925 91.935 ;
        RECT 21.575 91.665 21.910 91.935 ;
        RECT -290.655 4.295 -290.320 4.565 ;
        RECT -281.720 4.295 -281.385 4.565 ;
        RECT -280.735 4.295 -280.400 4.565 ;
        RECT -271.800 4.295 -271.465 4.565 ;
        RECT -270.815 4.295 -270.480 4.565 ;
        RECT -261.880 4.295 -261.545 4.565 ;
        RECT -260.895 4.295 -260.560 4.565 ;
        RECT -251.960 4.295 -251.625 4.565 ;
        RECT -250.975 4.295 -250.640 4.565 ;
        RECT -242.040 4.295 -241.705 4.565 ;
        RECT -241.055 4.295 -240.720 4.565 ;
        RECT -232.120 4.295 -231.785 4.565 ;
        RECT -231.135 4.295 -230.800 4.565 ;
        RECT -222.200 4.295 -221.865 4.565 ;
        RECT -221.215 4.295 -220.880 4.565 ;
        RECT -212.280 4.295 -211.945 4.565 ;
        RECT -211.295 4.295 -210.960 4.565 ;
        RECT -202.360 4.295 -202.025 4.565 ;
        RECT -201.375 4.295 -201.040 4.565 ;
        RECT -192.440 4.295 -192.105 4.565 ;
        RECT -191.455 4.295 -191.120 4.565 ;
        RECT -182.520 4.295 -182.185 4.565 ;
        RECT -181.535 4.295 -181.200 4.565 ;
        RECT -172.600 4.295 -172.265 4.565 ;
        RECT -171.615 4.295 -171.280 4.565 ;
        RECT -162.680 4.295 -162.345 4.565 ;
        RECT -161.695 4.295 -161.360 4.565 ;
        RECT -152.760 4.295 -152.425 4.565 ;
        RECT -151.775 4.295 -151.440 4.565 ;
        RECT -142.840 4.295 -142.505 4.565 ;
        RECT -141.855 4.295 -141.520 4.565 ;
        RECT -132.920 4.295 -132.585 4.565 ;
        RECT -131.935 4.295 -131.600 4.565 ;
        RECT -123.000 4.295 -122.665 4.565 ;
        RECT -122.015 4.295 -121.680 4.565 ;
        RECT -113.080 4.295 -112.745 4.565 ;
        RECT -112.095 4.295 -111.760 4.565 ;
        RECT -103.160 4.295 -102.825 4.565 ;
        RECT -102.175 4.295 -101.840 4.565 ;
        RECT -93.240 4.295 -92.905 4.565 ;
        RECT -92.255 4.295 -91.920 4.565 ;
        RECT -83.320 4.295 -82.985 4.565 ;
        RECT -82.335 4.295 -82.000 4.565 ;
        RECT -73.400 4.295 -73.065 4.565 ;
        RECT -72.415 4.295 -72.080 4.565 ;
        RECT -63.480 4.295 -63.145 4.565 ;
        RECT -62.495 4.295 -62.160 4.565 ;
        RECT -53.560 4.295 -53.225 4.565 ;
        RECT -52.575 4.295 -52.240 4.565 ;
        RECT -43.640 4.295 -43.305 4.565 ;
        RECT -42.655 4.295 -42.320 4.565 ;
        RECT -33.720 4.295 -33.385 4.565 ;
        RECT -32.735 4.295 -32.400 4.565 ;
        RECT -23.800 4.295 -23.465 4.565 ;
        RECT -22.815 4.295 -22.480 4.565 ;
        RECT -13.880 4.295 -13.545 4.565 ;
        RECT -12.895 4.295 -12.560 4.565 ;
        RECT -3.960 4.295 -3.625 4.565 ;
        RECT -2.975 4.295 -2.640 4.565 ;
        RECT 5.960 4.295 6.295 4.565 ;
        RECT 6.945 4.295 7.280 4.565 ;
        RECT 15.880 4.295 16.215 4.565 ;
        RECT 16.865 4.295 17.200 4.565 ;
        RECT 25.800 4.295 26.135 4.565 ;
        RECT -286.680 3.955 -286.345 4.225 ;
        RECT -285.695 3.955 -285.360 4.225 ;
        RECT -276.760 3.955 -276.425 4.225 ;
        RECT -275.775 3.955 -275.440 4.225 ;
        RECT -266.840 3.955 -266.505 4.225 ;
        RECT -265.855 3.955 -265.520 4.225 ;
        RECT -256.920 3.955 -256.585 4.225 ;
        RECT -255.935 3.955 -255.600 4.225 ;
        RECT -247.000 3.955 -246.665 4.225 ;
        RECT -246.015 3.955 -245.680 4.225 ;
        RECT -237.080 3.955 -236.745 4.225 ;
        RECT -236.095 3.955 -235.760 4.225 ;
        RECT -227.160 3.955 -226.825 4.225 ;
        RECT -226.175 3.955 -225.840 4.225 ;
        RECT -217.240 3.955 -216.905 4.225 ;
        RECT -216.255 3.955 -215.920 4.225 ;
        RECT -207.320 3.955 -206.985 4.225 ;
        RECT -206.335 3.955 -206.000 4.225 ;
        RECT -197.400 3.955 -197.065 4.225 ;
        RECT -196.415 3.955 -196.080 4.225 ;
        RECT -187.480 3.955 -187.145 4.225 ;
        RECT -186.495 3.955 -186.160 4.225 ;
        RECT -177.560 3.955 -177.225 4.225 ;
        RECT -176.575 3.955 -176.240 4.225 ;
        RECT -167.640 3.955 -167.305 4.225 ;
        RECT -166.655 3.955 -166.320 4.225 ;
        RECT -157.720 3.955 -157.385 4.225 ;
        RECT -156.735 3.955 -156.400 4.225 ;
        RECT -147.800 3.955 -147.465 4.225 ;
        RECT -146.815 3.955 -146.480 4.225 ;
        RECT -137.880 3.955 -137.545 4.225 ;
        RECT -136.895 3.955 -136.560 4.225 ;
        RECT -127.960 3.955 -127.625 4.225 ;
        RECT -126.975 3.955 -126.640 4.225 ;
        RECT -118.040 3.955 -117.705 4.225 ;
        RECT -117.055 3.955 -116.720 4.225 ;
        RECT -108.120 3.955 -107.785 4.225 ;
        RECT -107.135 3.955 -106.800 4.225 ;
        RECT -98.200 3.955 -97.865 4.225 ;
        RECT -97.215 3.955 -96.880 4.225 ;
        RECT -88.280 3.955 -87.945 4.225 ;
        RECT -87.295 3.955 -86.960 4.225 ;
        RECT -78.360 3.955 -78.025 4.225 ;
        RECT -77.375 3.955 -77.040 4.225 ;
        RECT -68.440 3.955 -68.105 4.225 ;
        RECT -67.455 3.955 -67.120 4.225 ;
        RECT -58.520 3.955 -58.185 4.225 ;
        RECT -57.535 3.955 -57.200 4.225 ;
        RECT -48.600 3.955 -48.265 4.225 ;
        RECT -47.615 3.955 -47.280 4.225 ;
        RECT -38.680 3.955 -38.345 4.225 ;
        RECT -37.695 3.955 -37.360 4.225 ;
        RECT -28.760 3.955 -28.425 4.225 ;
        RECT -27.775 3.955 -27.440 4.225 ;
        RECT -18.840 3.955 -18.505 4.225 ;
        RECT -17.855 3.955 -17.520 4.225 ;
        RECT -8.920 3.955 -8.585 4.225 ;
        RECT -7.935 3.955 -7.600 4.225 ;
        RECT 1.000 3.955 1.335 4.225 ;
        RECT 1.985 3.955 2.320 4.225 ;
        RECT 10.920 3.955 11.255 4.225 ;
        RECT 11.905 3.955 12.240 4.225 ;
        RECT 20.840 3.955 21.175 4.225 ;
        RECT 21.825 3.955 22.160 4.225 ;
        RECT -288.895 -89.055 -288.560 -88.785 ;
        RECT -279.960 -89.055 -279.625 -88.785 ;
        RECT -278.975 -89.055 -278.640 -88.785 ;
        RECT -270.040 -89.055 -269.705 -88.785 ;
        RECT -269.055 -89.055 -268.720 -88.785 ;
        RECT -260.120 -89.055 -259.785 -88.785 ;
        RECT -259.135 -89.055 -258.800 -88.785 ;
        RECT -250.200 -89.055 -249.865 -88.785 ;
        RECT -249.215 -89.055 -248.880 -88.785 ;
        RECT -240.280 -89.055 -239.945 -88.785 ;
        RECT -239.295 -89.055 -238.960 -88.785 ;
        RECT -230.360 -89.055 -230.025 -88.785 ;
        RECT -229.375 -89.055 -229.040 -88.785 ;
        RECT -220.440 -89.055 -220.105 -88.785 ;
        RECT -219.455 -89.055 -219.120 -88.785 ;
        RECT -210.520 -89.055 -210.185 -88.785 ;
        RECT -209.535 -89.055 -209.200 -88.785 ;
        RECT -200.600 -89.055 -200.265 -88.785 ;
        RECT -199.615 -89.055 -199.280 -88.785 ;
        RECT -190.680 -89.055 -190.345 -88.785 ;
        RECT -189.695 -89.055 -189.360 -88.785 ;
        RECT -180.760 -89.055 -180.425 -88.785 ;
        RECT -179.775 -89.055 -179.440 -88.785 ;
        RECT -170.840 -89.055 -170.505 -88.785 ;
        RECT -169.855 -89.055 -169.520 -88.785 ;
        RECT -160.920 -89.055 -160.585 -88.785 ;
        RECT -159.935 -89.055 -159.600 -88.785 ;
        RECT -151.000 -89.055 -150.665 -88.785 ;
        RECT -150.015 -89.055 -149.680 -88.785 ;
        RECT -141.080 -89.055 -140.745 -88.785 ;
        RECT -140.095 -89.055 -139.760 -88.785 ;
        RECT -131.160 -89.055 -130.825 -88.785 ;
        RECT -130.175 -89.055 -129.840 -88.785 ;
        RECT -121.240 -89.055 -120.905 -88.785 ;
        RECT -120.255 -89.055 -119.920 -88.785 ;
        RECT -111.320 -89.055 -110.985 -88.785 ;
        RECT -110.335 -89.055 -110.000 -88.785 ;
        RECT -101.400 -89.055 -101.065 -88.785 ;
        RECT -100.415 -89.055 -100.080 -88.785 ;
        RECT -91.480 -89.055 -91.145 -88.785 ;
        RECT -90.495 -89.055 -90.160 -88.785 ;
        RECT -81.560 -89.055 -81.225 -88.785 ;
        RECT -80.575 -89.055 -80.240 -88.785 ;
        RECT -71.640 -89.055 -71.305 -88.785 ;
        RECT -70.655 -89.055 -70.320 -88.785 ;
        RECT -61.720 -89.055 -61.385 -88.785 ;
        RECT -60.735 -89.055 -60.400 -88.785 ;
        RECT -51.800 -89.055 -51.465 -88.785 ;
        RECT -50.815 -89.055 -50.480 -88.785 ;
        RECT -41.880 -89.055 -41.545 -88.785 ;
        RECT -40.895 -89.055 -40.560 -88.785 ;
        RECT -31.960 -89.055 -31.625 -88.785 ;
        RECT -30.975 -89.055 -30.640 -88.785 ;
        RECT -22.040 -89.055 -21.705 -88.785 ;
        RECT -21.055 -89.055 -20.720 -88.785 ;
        RECT -12.120 -89.055 -11.785 -88.785 ;
        RECT -11.135 -89.055 -10.800 -88.785 ;
        RECT -2.200 -89.055 -1.865 -88.785 ;
        RECT -1.215 -89.055 -0.880 -88.785 ;
        RECT 7.720 -89.055 8.055 -88.785 ;
        RECT 8.705 -89.055 9.040 -88.785 ;
        RECT 17.640 -89.055 17.975 -88.785 ;
        RECT 18.625 -89.055 18.960 -88.785 ;
        RECT 27.560 -89.055 27.895 -88.785 ;
        RECT -284.920 -89.395 -284.585 -89.125 ;
        RECT -283.935 -89.395 -283.600 -89.125 ;
        RECT -275.000 -89.395 -274.665 -89.125 ;
        RECT -274.015 -89.395 -273.680 -89.125 ;
        RECT -265.080 -89.395 -264.745 -89.125 ;
        RECT -264.095 -89.395 -263.760 -89.125 ;
        RECT -255.160 -89.395 -254.825 -89.125 ;
        RECT -254.175 -89.395 -253.840 -89.125 ;
        RECT -245.240 -89.395 -244.905 -89.125 ;
        RECT -244.255 -89.395 -243.920 -89.125 ;
        RECT -235.320 -89.395 -234.985 -89.125 ;
        RECT -234.335 -89.395 -234.000 -89.125 ;
        RECT -225.400 -89.395 -225.065 -89.125 ;
        RECT -224.415 -89.395 -224.080 -89.125 ;
        RECT -215.480 -89.395 -215.145 -89.125 ;
        RECT -214.495 -89.395 -214.160 -89.125 ;
        RECT -205.560 -89.395 -205.225 -89.125 ;
        RECT -204.575 -89.395 -204.240 -89.125 ;
        RECT -195.640 -89.395 -195.305 -89.125 ;
        RECT -194.655 -89.395 -194.320 -89.125 ;
        RECT -185.720 -89.395 -185.385 -89.125 ;
        RECT -184.735 -89.395 -184.400 -89.125 ;
        RECT -175.800 -89.395 -175.465 -89.125 ;
        RECT -174.815 -89.395 -174.480 -89.125 ;
        RECT -165.880 -89.395 -165.545 -89.125 ;
        RECT -164.895 -89.395 -164.560 -89.125 ;
        RECT -155.960 -89.395 -155.625 -89.125 ;
        RECT -154.975 -89.395 -154.640 -89.125 ;
        RECT -146.040 -89.395 -145.705 -89.125 ;
        RECT -145.055 -89.395 -144.720 -89.125 ;
        RECT -136.120 -89.395 -135.785 -89.125 ;
        RECT -135.135 -89.395 -134.800 -89.125 ;
        RECT -126.200 -89.395 -125.865 -89.125 ;
        RECT -125.215 -89.395 -124.880 -89.125 ;
        RECT -116.280 -89.395 -115.945 -89.125 ;
        RECT -115.295 -89.395 -114.960 -89.125 ;
        RECT -106.360 -89.395 -106.025 -89.125 ;
        RECT -105.375 -89.395 -105.040 -89.125 ;
        RECT -96.440 -89.395 -96.105 -89.125 ;
        RECT -95.455 -89.395 -95.120 -89.125 ;
        RECT -86.520 -89.395 -86.185 -89.125 ;
        RECT -85.535 -89.395 -85.200 -89.125 ;
        RECT -76.600 -89.395 -76.265 -89.125 ;
        RECT -75.615 -89.395 -75.280 -89.125 ;
        RECT -66.680 -89.395 -66.345 -89.125 ;
        RECT -65.695 -89.395 -65.360 -89.125 ;
        RECT -56.760 -89.395 -56.425 -89.125 ;
        RECT -55.775 -89.395 -55.440 -89.125 ;
        RECT -46.840 -89.395 -46.505 -89.125 ;
        RECT -45.855 -89.395 -45.520 -89.125 ;
        RECT -36.920 -89.395 -36.585 -89.125 ;
        RECT -35.935 -89.395 -35.600 -89.125 ;
        RECT -27.000 -89.395 -26.665 -89.125 ;
        RECT -26.015 -89.395 -25.680 -89.125 ;
        RECT -17.080 -89.395 -16.745 -89.125 ;
        RECT -16.095 -89.395 -15.760 -89.125 ;
        RECT -7.160 -89.395 -6.825 -89.125 ;
        RECT -6.175 -89.395 -5.840 -89.125 ;
        RECT 2.760 -89.395 3.095 -89.125 ;
        RECT 3.745 -89.395 4.080 -89.125 ;
        RECT 12.680 -89.395 13.015 -89.125 ;
        RECT 13.665 -89.395 14.000 -89.125 ;
        RECT 22.600 -89.395 22.935 -89.125 ;
        RECT 23.585 -89.395 23.920 -89.125 ;
        RECT -288.645 -176.765 -288.310 -176.495 ;
        RECT -279.710 -176.765 -279.375 -176.495 ;
        RECT -278.725 -176.765 -278.390 -176.495 ;
        RECT -269.790 -176.765 -269.455 -176.495 ;
        RECT -268.805 -176.765 -268.470 -176.495 ;
        RECT -259.870 -176.765 -259.535 -176.495 ;
        RECT -258.885 -176.765 -258.550 -176.495 ;
        RECT -249.950 -176.765 -249.615 -176.495 ;
        RECT -248.965 -176.765 -248.630 -176.495 ;
        RECT -240.030 -176.765 -239.695 -176.495 ;
        RECT -239.045 -176.765 -238.710 -176.495 ;
        RECT -230.110 -176.765 -229.775 -176.495 ;
        RECT -229.125 -176.765 -228.790 -176.495 ;
        RECT -220.190 -176.765 -219.855 -176.495 ;
        RECT -219.205 -176.765 -218.870 -176.495 ;
        RECT -210.270 -176.765 -209.935 -176.495 ;
        RECT -209.285 -176.765 -208.950 -176.495 ;
        RECT -200.350 -176.765 -200.015 -176.495 ;
        RECT -199.365 -176.765 -199.030 -176.495 ;
        RECT -190.430 -176.765 -190.095 -176.495 ;
        RECT -189.445 -176.765 -189.110 -176.495 ;
        RECT -180.510 -176.765 -180.175 -176.495 ;
        RECT -179.525 -176.765 -179.190 -176.495 ;
        RECT -170.590 -176.765 -170.255 -176.495 ;
        RECT -169.605 -176.765 -169.270 -176.495 ;
        RECT -160.670 -176.765 -160.335 -176.495 ;
        RECT -159.685 -176.765 -159.350 -176.495 ;
        RECT -150.750 -176.765 -150.415 -176.495 ;
        RECT -149.765 -176.765 -149.430 -176.495 ;
        RECT -140.830 -176.765 -140.495 -176.495 ;
        RECT -139.845 -176.765 -139.510 -176.495 ;
        RECT -130.910 -176.765 -130.575 -176.495 ;
        RECT -129.925 -176.765 -129.590 -176.495 ;
        RECT -120.990 -176.765 -120.655 -176.495 ;
        RECT -120.005 -176.765 -119.670 -176.495 ;
        RECT -111.070 -176.765 -110.735 -176.495 ;
        RECT -110.085 -176.765 -109.750 -176.495 ;
        RECT -101.150 -176.765 -100.815 -176.495 ;
        RECT -100.165 -176.765 -99.830 -176.495 ;
        RECT -91.230 -176.765 -90.895 -176.495 ;
        RECT -90.245 -176.765 -89.910 -176.495 ;
        RECT -81.310 -176.765 -80.975 -176.495 ;
        RECT -80.325 -176.765 -79.990 -176.495 ;
        RECT -71.390 -176.765 -71.055 -176.495 ;
        RECT -70.405 -176.765 -70.070 -176.495 ;
        RECT -61.470 -176.765 -61.135 -176.495 ;
        RECT -60.485 -176.765 -60.150 -176.495 ;
        RECT -51.550 -176.765 -51.215 -176.495 ;
        RECT -50.565 -176.765 -50.230 -176.495 ;
        RECT -41.630 -176.765 -41.295 -176.495 ;
        RECT -40.645 -176.765 -40.310 -176.495 ;
        RECT -31.710 -176.765 -31.375 -176.495 ;
        RECT -30.725 -176.765 -30.390 -176.495 ;
        RECT -21.790 -176.765 -21.455 -176.495 ;
        RECT -20.805 -176.765 -20.470 -176.495 ;
        RECT -11.870 -176.765 -11.535 -176.495 ;
        RECT -10.885 -176.765 -10.550 -176.495 ;
        RECT -1.950 -176.765 -1.615 -176.495 ;
        RECT -0.965 -176.765 -0.630 -176.495 ;
        RECT 7.970 -176.765 8.305 -176.495 ;
        RECT 8.955 -176.765 9.290 -176.495 ;
        RECT 17.890 -176.765 18.225 -176.495 ;
        RECT 18.875 -176.765 19.210 -176.495 ;
        RECT 27.810 -176.765 28.145 -176.495 ;
        RECT -284.670 -177.105 -284.335 -176.835 ;
        RECT -283.685 -177.105 -283.350 -176.835 ;
        RECT -274.750 -177.105 -274.415 -176.835 ;
        RECT -273.765 -177.105 -273.430 -176.835 ;
        RECT -264.830 -177.105 -264.495 -176.835 ;
        RECT -263.845 -177.105 -263.510 -176.835 ;
        RECT -254.910 -177.105 -254.575 -176.835 ;
        RECT -253.925 -177.105 -253.590 -176.835 ;
        RECT -244.990 -177.105 -244.655 -176.835 ;
        RECT -244.005 -177.105 -243.670 -176.835 ;
        RECT -235.070 -177.105 -234.735 -176.835 ;
        RECT -234.085 -177.105 -233.750 -176.835 ;
        RECT -225.150 -177.105 -224.815 -176.835 ;
        RECT -224.165 -177.105 -223.830 -176.835 ;
        RECT -215.230 -177.105 -214.895 -176.835 ;
        RECT -214.245 -177.105 -213.910 -176.835 ;
        RECT -205.310 -177.105 -204.975 -176.835 ;
        RECT -204.325 -177.105 -203.990 -176.835 ;
        RECT -195.390 -177.105 -195.055 -176.835 ;
        RECT -194.405 -177.105 -194.070 -176.835 ;
        RECT -185.470 -177.105 -185.135 -176.835 ;
        RECT -184.485 -177.105 -184.150 -176.835 ;
        RECT -175.550 -177.105 -175.215 -176.835 ;
        RECT -174.565 -177.105 -174.230 -176.835 ;
        RECT -165.630 -177.105 -165.295 -176.835 ;
        RECT -164.645 -177.105 -164.310 -176.835 ;
        RECT -155.710 -177.105 -155.375 -176.835 ;
        RECT -154.725 -177.105 -154.390 -176.835 ;
        RECT -145.790 -177.105 -145.455 -176.835 ;
        RECT -144.805 -177.105 -144.470 -176.835 ;
        RECT -135.870 -177.105 -135.535 -176.835 ;
        RECT -134.885 -177.105 -134.550 -176.835 ;
        RECT -125.950 -177.105 -125.615 -176.835 ;
        RECT -124.965 -177.105 -124.630 -176.835 ;
        RECT -116.030 -177.105 -115.695 -176.835 ;
        RECT -115.045 -177.105 -114.710 -176.835 ;
        RECT -106.110 -177.105 -105.775 -176.835 ;
        RECT -105.125 -177.105 -104.790 -176.835 ;
        RECT -96.190 -177.105 -95.855 -176.835 ;
        RECT -95.205 -177.105 -94.870 -176.835 ;
        RECT -86.270 -177.105 -85.935 -176.835 ;
        RECT -85.285 -177.105 -84.950 -176.835 ;
        RECT -76.350 -177.105 -76.015 -176.835 ;
        RECT -75.365 -177.105 -75.030 -176.835 ;
        RECT -66.430 -177.105 -66.095 -176.835 ;
        RECT -65.445 -177.105 -65.110 -176.835 ;
        RECT -56.510 -177.105 -56.175 -176.835 ;
        RECT -55.525 -177.105 -55.190 -176.835 ;
        RECT -46.590 -177.105 -46.255 -176.835 ;
        RECT -45.605 -177.105 -45.270 -176.835 ;
        RECT -36.670 -177.105 -36.335 -176.835 ;
        RECT -35.685 -177.105 -35.350 -176.835 ;
        RECT -26.750 -177.105 -26.415 -176.835 ;
        RECT -25.765 -177.105 -25.430 -176.835 ;
        RECT -16.830 -177.105 -16.495 -176.835 ;
        RECT -15.845 -177.105 -15.510 -176.835 ;
        RECT -6.910 -177.105 -6.575 -176.835 ;
        RECT -5.925 -177.105 -5.590 -176.835 ;
        RECT 3.010 -177.105 3.345 -176.835 ;
        RECT 3.995 -177.105 4.330 -176.835 ;
        RECT 12.930 -177.105 13.265 -176.835 ;
        RECT 13.915 -177.105 14.250 -176.835 ;
        RECT 22.850 -177.105 23.185 -176.835 ;
        RECT 23.835 -177.105 24.170 -176.835 ;
      LAYER mcon ;
        RECT -290.820 92.085 -290.650 92.255 ;
        RECT -281.890 92.085 -281.720 92.255 ;
        RECT -280.900 92.085 -280.730 92.255 ;
        RECT -271.970 92.085 -271.800 92.255 ;
        RECT -270.980 92.085 -270.810 92.255 ;
        RECT -262.050 92.085 -261.880 92.255 ;
        RECT -261.060 92.085 -260.890 92.255 ;
        RECT -252.130 92.085 -251.960 92.255 ;
        RECT -251.140 92.085 -250.970 92.255 ;
        RECT -242.210 92.085 -242.040 92.255 ;
        RECT -241.220 92.085 -241.050 92.255 ;
        RECT -232.290 92.085 -232.120 92.255 ;
        RECT -231.300 92.085 -231.130 92.255 ;
        RECT -222.370 92.085 -222.200 92.255 ;
        RECT -221.380 92.085 -221.210 92.255 ;
        RECT -212.450 92.085 -212.280 92.255 ;
        RECT -211.460 92.085 -211.290 92.255 ;
        RECT -202.530 92.085 -202.360 92.255 ;
        RECT -201.540 92.085 -201.370 92.255 ;
        RECT -192.610 92.085 -192.440 92.255 ;
        RECT -191.620 92.085 -191.450 92.255 ;
        RECT -182.690 92.085 -182.520 92.255 ;
        RECT -181.700 92.085 -181.530 92.255 ;
        RECT -172.770 92.085 -172.600 92.255 ;
        RECT -171.780 92.085 -171.610 92.255 ;
        RECT -162.850 92.085 -162.680 92.255 ;
        RECT -161.860 92.085 -161.690 92.255 ;
        RECT -152.930 92.085 -152.760 92.255 ;
        RECT -151.940 92.085 -151.770 92.255 ;
        RECT -143.010 92.085 -142.840 92.255 ;
        RECT -142.020 92.085 -141.850 92.255 ;
        RECT -133.090 92.085 -132.920 92.255 ;
        RECT -132.100 92.085 -131.930 92.255 ;
        RECT -123.170 92.085 -123.000 92.255 ;
        RECT -122.180 92.085 -122.010 92.255 ;
        RECT -113.250 92.085 -113.080 92.255 ;
        RECT -112.260 92.085 -112.090 92.255 ;
        RECT -103.330 92.085 -103.160 92.255 ;
        RECT -102.340 92.085 -102.170 92.255 ;
        RECT -93.410 92.085 -93.240 92.255 ;
        RECT -92.420 92.085 -92.250 92.255 ;
        RECT -83.490 92.085 -83.320 92.255 ;
        RECT -82.500 92.085 -82.330 92.255 ;
        RECT -73.570 92.085 -73.400 92.255 ;
        RECT -72.580 92.085 -72.410 92.255 ;
        RECT -63.650 92.085 -63.480 92.255 ;
        RECT -62.660 92.085 -62.490 92.255 ;
        RECT -53.730 92.085 -53.560 92.255 ;
        RECT -52.740 92.085 -52.570 92.255 ;
        RECT -43.810 92.085 -43.640 92.255 ;
        RECT -42.820 92.085 -42.650 92.255 ;
        RECT -33.890 92.085 -33.720 92.255 ;
        RECT -32.900 92.085 -32.730 92.255 ;
        RECT -23.970 92.085 -23.800 92.255 ;
        RECT -22.980 92.085 -22.810 92.255 ;
        RECT -14.050 92.085 -13.880 92.255 ;
        RECT -13.060 92.085 -12.890 92.255 ;
        RECT -4.130 92.085 -3.960 92.255 ;
        RECT -3.140 92.085 -2.970 92.255 ;
        RECT 5.790 92.085 5.960 92.255 ;
        RECT 6.780 92.085 6.950 92.255 ;
        RECT 15.710 92.085 15.880 92.255 ;
        RECT 16.700 92.085 16.870 92.255 ;
        RECT 25.630 92.085 25.800 92.255 ;
        RECT -286.850 91.685 -286.680 91.855 ;
        RECT -285.860 91.685 -285.690 91.855 ;
        RECT -276.930 91.685 -276.760 91.855 ;
        RECT -275.940 91.685 -275.770 91.855 ;
        RECT -267.010 91.685 -266.840 91.855 ;
        RECT -266.020 91.685 -265.850 91.855 ;
        RECT -257.090 91.685 -256.920 91.855 ;
        RECT -256.100 91.685 -255.930 91.855 ;
        RECT -247.170 91.685 -247.000 91.855 ;
        RECT -246.180 91.685 -246.010 91.855 ;
        RECT -237.250 91.685 -237.080 91.855 ;
        RECT -236.260 91.685 -236.090 91.855 ;
        RECT -227.330 91.685 -227.160 91.855 ;
        RECT -226.340 91.685 -226.170 91.855 ;
        RECT -217.410 91.685 -217.240 91.855 ;
        RECT -216.420 91.685 -216.250 91.855 ;
        RECT -207.490 91.685 -207.320 91.855 ;
        RECT -206.500 91.685 -206.330 91.855 ;
        RECT -197.570 91.685 -197.400 91.855 ;
        RECT -196.580 91.685 -196.410 91.855 ;
        RECT -187.650 91.685 -187.480 91.855 ;
        RECT -186.660 91.685 -186.490 91.855 ;
        RECT -177.730 91.685 -177.560 91.855 ;
        RECT -176.740 91.685 -176.570 91.855 ;
        RECT -167.810 91.685 -167.640 91.855 ;
        RECT -166.820 91.685 -166.650 91.855 ;
        RECT -157.890 91.685 -157.720 91.855 ;
        RECT -156.900 91.685 -156.730 91.855 ;
        RECT -147.970 91.685 -147.800 91.855 ;
        RECT -146.980 91.685 -146.810 91.855 ;
        RECT -138.050 91.685 -137.880 91.855 ;
        RECT -137.060 91.685 -136.890 91.855 ;
        RECT -128.130 91.685 -127.960 91.855 ;
        RECT -127.140 91.685 -126.970 91.855 ;
        RECT -118.210 91.685 -118.040 91.855 ;
        RECT -117.220 91.685 -117.050 91.855 ;
        RECT -108.290 91.685 -108.120 91.855 ;
        RECT -107.300 91.685 -107.130 91.855 ;
        RECT -98.370 91.685 -98.200 91.855 ;
        RECT -97.380 91.685 -97.210 91.855 ;
        RECT -88.450 91.685 -88.280 91.855 ;
        RECT -87.460 91.685 -87.290 91.855 ;
        RECT -78.530 91.685 -78.360 91.855 ;
        RECT -77.540 91.685 -77.370 91.855 ;
        RECT -68.610 91.685 -68.440 91.855 ;
        RECT -67.620 91.685 -67.450 91.855 ;
        RECT -58.690 91.685 -58.520 91.855 ;
        RECT -57.700 91.685 -57.530 91.855 ;
        RECT -48.770 91.685 -48.600 91.855 ;
        RECT -47.780 91.685 -47.610 91.855 ;
        RECT -38.850 91.685 -38.680 91.855 ;
        RECT -37.860 91.685 -37.690 91.855 ;
        RECT -28.930 91.685 -28.760 91.855 ;
        RECT -27.940 91.685 -27.770 91.855 ;
        RECT -19.010 91.685 -18.840 91.855 ;
        RECT -18.020 91.685 -17.850 91.855 ;
        RECT -9.090 91.685 -8.920 91.855 ;
        RECT -8.100 91.685 -7.930 91.855 ;
        RECT 0.830 91.685 1.000 91.855 ;
        RECT 1.820 91.685 1.990 91.855 ;
        RECT 10.750 91.685 10.920 91.855 ;
        RECT 11.740 91.685 11.910 91.855 ;
        RECT 20.670 91.685 20.840 91.855 ;
        RECT 21.660 91.685 21.830 91.855 ;
        RECT -290.570 4.375 -290.400 4.545 ;
        RECT -281.640 4.375 -281.470 4.545 ;
        RECT -280.650 4.375 -280.480 4.545 ;
        RECT -271.720 4.375 -271.550 4.545 ;
        RECT -270.730 4.375 -270.560 4.545 ;
        RECT -261.800 4.375 -261.630 4.545 ;
        RECT -260.810 4.375 -260.640 4.545 ;
        RECT -251.880 4.375 -251.710 4.545 ;
        RECT -250.890 4.375 -250.720 4.545 ;
        RECT -241.960 4.375 -241.790 4.545 ;
        RECT -240.970 4.375 -240.800 4.545 ;
        RECT -232.040 4.375 -231.870 4.545 ;
        RECT -231.050 4.375 -230.880 4.545 ;
        RECT -222.120 4.375 -221.950 4.545 ;
        RECT -221.130 4.375 -220.960 4.545 ;
        RECT -212.200 4.375 -212.030 4.545 ;
        RECT -211.210 4.375 -211.040 4.545 ;
        RECT -202.280 4.375 -202.110 4.545 ;
        RECT -201.290 4.375 -201.120 4.545 ;
        RECT -192.360 4.375 -192.190 4.545 ;
        RECT -191.370 4.375 -191.200 4.545 ;
        RECT -182.440 4.375 -182.270 4.545 ;
        RECT -181.450 4.375 -181.280 4.545 ;
        RECT -172.520 4.375 -172.350 4.545 ;
        RECT -171.530 4.375 -171.360 4.545 ;
        RECT -162.600 4.375 -162.430 4.545 ;
        RECT -161.610 4.375 -161.440 4.545 ;
        RECT -152.680 4.375 -152.510 4.545 ;
        RECT -151.690 4.375 -151.520 4.545 ;
        RECT -142.760 4.375 -142.590 4.545 ;
        RECT -141.770 4.375 -141.600 4.545 ;
        RECT -132.840 4.375 -132.670 4.545 ;
        RECT -131.850 4.375 -131.680 4.545 ;
        RECT -122.920 4.375 -122.750 4.545 ;
        RECT -121.930 4.375 -121.760 4.545 ;
        RECT -113.000 4.375 -112.830 4.545 ;
        RECT -112.010 4.375 -111.840 4.545 ;
        RECT -103.080 4.375 -102.910 4.545 ;
        RECT -102.090 4.375 -101.920 4.545 ;
        RECT -93.160 4.375 -92.990 4.545 ;
        RECT -92.170 4.375 -92.000 4.545 ;
        RECT -83.240 4.375 -83.070 4.545 ;
        RECT -82.250 4.375 -82.080 4.545 ;
        RECT -73.320 4.375 -73.150 4.545 ;
        RECT -72.330 4.375 -72.160 4.545 ;
        RECT -63.400 4.375 -63.230 4.545 ;
        RECT -62.410 4.375 -62.240 4.545 ;
        RECT -53.480 4.375 -53.310 4.545 ;
        RECT -52.490 4.375 -52.320 4.545 ;
        RECT -43.560 4.375 -43.390 4.545 ;
        RECT -42.570 4.375 -42.400 4.545 ;
        RECT -33.640 4.375 -33.470 4.545 ;
        RECT -32.650 4.375 -32.480 4.545 ;
        RECT -23.720 4.375 -23.550 4.545 ;
        RECT -22.730 4.375 -22.560 4.545 ;
        RECT -13.800 4.375 -13.630 4.545 ;
        RECT -12.810 4.375 -12.640 4.545 ;
        RECT -3.880 4.375 -3.710 4.545 ;
        RECT -2.890 4.375 -2.720 4.545 ;
        RECT 6.040 4.375 6.210 4.545 ;
        RECT 7.030 4.375 7.200 4.545 ;
        RECT 15.960 4.375 16.130 4.545 ;
        RECT 16.950 4.375 17.120 4.545 ;
        RECT 25.880 4.375 26.050 4.545 ;
        RECT -286.600 3.975 -286.430 4.145 ;
        RECT -285.610 3.975 -285.440 4.145 ;
        RECT -276.680 3.975 -276.510 4.145 ;
        RECT -275.690 3.975 -275.520 4.145 ;
        RECT -266.760 3.975 -266.590 4.145 ;
        RECT -265.770 3.975 -265.600 4.145 ;
        RECT -256.840 3.975 -256.670 4.145 ;
        RECT -255.850 3.975 -255.680 4.145 ;
        RECT -246.920 3.975 -246.750 4.145 ;
        RECT -245.930 3.975 -245.760 4.145 ;
        RECT -237.000 3.975 -236.830 4.145 ;
        RECT -236.010 3.975 -235.840 4.145 ;
        RECT -227.080 3.975 -226.910 4.145 ;
        RECT -226.090 3.975 -225.920 4.145 ;
        RECT -217.160 3.975 -216.990 4.145 ;
        RECT -216.170 3.975 -216.000 4.145 ;
        RECT -207.240 3.975 -207.070 4.145 ;
        RECT -206.250 3.975 -206.080 4.145 ;
        RECT -197.320 3.975 -197.150 4.145 ;
        RECT -196.330 3.975 -196.160 4.145 ;
        RECT -187.400 3.975 -187.230 4.145 ;
        RECT -186.410 3.975 -186.240 4.145 ;
        RECT -177.480 3.975 -177.310 4.145 ;
        RECT -176.490 3.975 -176.320 4.145 ;
        RECT -167.560 3.975 -167.390 4.145 ;
        RECT -166.570 3.975 -166.400 4.145 ;
        RECT -157.640 3.975 -157.470 4.145 ;
        RECT -156.650 3.975 -156.480 4.145 ;
        RECT -147.720 3.975 -147.550 4.145 ;
        RECT -146.730 3.975 -146.560 4.145 ;
        RECT -137.800 3.975 -137.630 4.145 ;
        RECT -136.810 3.975 -136.640 4.145 ;
        RECT -127.880 3.975 -127.710 4.145 ;
        RECT -126.890 3.975 -126.720 4.145 ;
        RECT -117.960 3.975 -117.790 4.145 ;
        RECT -116.970 3.975 -116.800 4.145 ;
        RECT -108.040 3.975 -107.870 4.145 ;
        RECT -107.050 3.975 -106.880 4.145 ;
        RECT -98.120 3.975 -97.950 4.145 ;
        RECT -97.130 3.975 -96.960 4.145 ;
        RECT -88.200 3.975 -88.030 4.145 ;
        RECT -87.210 3.975 -87.040 4.145 ;
        RECT -78.280 3.975 -78.110 4.145 ;
        RECT -77.290 3.975 -77.120 4.145 ;
        RECT -68.360 3.975 -68.190 4.145 ;
        RECT -67.370 3.975 -67.200 4.145 ;
        RECT -58.440 3.975 -58.270 4.145 ;
        RECT -57.450 3.975 -57.280 4.145 ;
        RECT -48.520 3.975 -48.350 4.145 ;
        RECT -47.530 3.975 -47.360 4.145 ;
        RECT -38.600 3.975 -38.430 4.145 ;
        RECT -37.610 3.975 -37.440 4.145 ;
        RECT -28.680 3.975 -28.510 4.145 ;
        RECT -27.690 3.975 -27.520 4.145 ;
        RECT -18.760 3.975 -18.590 4.145 ;
        RECT -17.770 3.975 -17.600 4.145 ;
        RECT -8.840 3.975 -8.670 4.145 ;
        RECT -7.850 3.975 -7.680 4.145 ;
        RECT 1.080 3.975 1.250 4.145 ;
        RECT 2.070 3.975 2.240 4.145 ;
        RECT 11.000 3.975 11.170 4.145 ;
        RECT 11.990 3.975 12.160 4.145 ;
        RECT 20.920 3.975 21.090 4.145 ;
        RECT 21.910 3.975 22.080 4.145 ;
        RECT -288.810 -88.975 -288.640 -88.805 ;
        RECT -279.880 -88.975 -279.710 -88.805 ;
        RECT -278.890 -88.975 -278.720 -88.805 ;
        RECT -269.960 -88.975 -269.790 -88.805 ;
        RECT -268.970 -88.975 -268.800 -88.805 ;
        RECT -260.040 -88.975 -259.870 -88.805 ;
        RECT -259.050 -88.975 -258.880 -88.805 ;
        RECT -250.120 -88.975 -249.950 -88.805 ;
        RECT -249.130 -88.975 -248.960 -88.805 ;
        RECT -240.200 -88.975 -240.030 -88.805 ;
        RECT -239.210 -88.975 -239.040 -88.805 ;
        RECT -230.280 -88.975 -230.110 -88.805 ;
        RECT -229.290 -88.975 -229.120 -88.805 ;
        RECT -220.360 -88.975 -220.190 -88.805 ;
        RECT -219.370 -88.975 -219.200 -88.805 ;
        RECT -210.440 -88.975 -210.270 -88.805 ;
        RECT -209.450 -88.975 -209.280 -88.805 ;
        RECT -200.520 -88.975 -200.350 -88.805 ;
        RECT -199.530 -88.975 -199.360 -88.805 ;
        RECT -190.600 -88.975 -190.430 -88.805 ;
        RECT -189.610 -88.975 -189.440 -88.805 ;
        RECT -180.680 -88.975 -180.510 -88.805 ;
        RECT -179.690 -88.975 -179.520 -88.805 ;
        RECT -170.760 -88.975 -170.590 -88.805 ;
        RECT -169.770 -88.975 -169.600 -88.805 ;
        RECT -160.840 -88.975 -160.670 -88.805 ;
        RECT -159.850 -88.975 -159.680 -88.805 ;
        RECT -150.920 -88.975 -150.750 -88.805 ;
        RECT -149.930 -88.975 -149.760 -88.805 ;
        RECT -141.000 -88.975 -140.830 -88.805 ;
        RECT -140.010 -88.975 -139.840 -88.805 ;
        RECT -131.080 -88.975 -130.910 -88.805 ;
        RECT -130.090 -88.975 -129.920 -88.805 ;
        RECT -121.160 -88.975 -120.990 -88.805 ;
        RECT -120.170 -88.975 -120.000 -88.805 ;
        RECT -111.240 -88.975 -111.070 -88.805 ;
        RECT -110.250 -88.975 -110.080 -88.805 ;
        RECT -101.320 -88.975 -101.150 -88.805 ;
        RECT -100.330 -88.975 -100.160 -88.805 ;
        RECT -91.400 -88.975 -91.230 -88.805 ;
        RECT -90.410 -88.975 -90.240 -88.805 ;
        RECT -81.480 -88.975 -81.310 -88.805 ;
        RECT -80.490 -88.975 -80.320 -88.805 ;
        RECT -71.560 -88.975 -71.390 -88.805 ;
        RECT -70.570 -88.975 -70.400 -88.805 ;
        RECT -61.640 -88.975 -61.470 -88.805 ;
        RECT -60.650 -88.975 -60.480 -88.805 ;
        RECT -51.720 -88.975 -51.550 -88.805 ;
        RECT -50.730 -88.975 -50.560 -88.805 ;
        RECT -41.800 -88.975 -41.630 -88.805 ;
        RECT -40.810 -88.975 -40.640 -88.805 ;
        RECT -31.880 -88.975 -31.710 -88.805 ;
        RECT -30.890 -88.975 -30.720 -88.805 ;
        RECT -21.960 -88.975 -21.790 -88.805 ;
        RECT -20.970 -88.975 -20.800 -88.805 ;
        RECT -12.040 -88.975 -11.870 -88.805 ;
        RECT -11.050 -88.975 -10.880 -88.805 ;
        RECT -2.120 -88.975 -1.950 -88.805 ;
        RECT -1.130 -88.975 -0.960 -88.805 ;
        RECT 7.800 -88.975 7.970 -88.805 ;
        RECT 8.790 -88.975 8.960 -88.805 ;
        RECT 17.720 -88.975 17.890 -88.805 ;
        RECT 18.710 -88.975 18.880 -88.805 ;
        RECT 27.640 -88.975 27.810 -88.805 ;
        RECT -284.840 -89.375 -284.670 -89.205 ;
        RECT -283.850 -89.375 -283.680 -89.205 ;
        RECT -274.920 -89.375 -274.750 -89.205 ;
        RECT -273.930 -89.375 -273.760 -89.205 ;
        RECT -265.000 -89.375 -264.830 -89.205 ;
        RECT -264.010 -89.375 -263.840 -89.205 ;
        RECT -255.080 -89.375 -254.910 -89.205 ;
        RECT -254.090 -89.375 -253.920 -89.205 ;
        RECT -245.160 -89.375 -244.990 -89.205 ;
        RECT -244.170 -89.375 -244.000 -89.205 ;
        RECT -235.240 -89.375 -235.070 -89.205 ;
        RECT -234.250 -89.375 -234.080 -89.205 ;
        RECT -225.320 -89.375 -225.150 -89.205 ;
        RECT -224.330 -89.375 -224.160 -89.205 ;
        RECT -215.400 -89.375 -215.230 -89.205 ;
        RECT -214.410 -89.375 -214.240 -89.205 ;
        RECT -205.480 -89.375 -205.310 -89.205 ;
        RECT -204.490 -89.375 -204.320 -89.205 ;
        RECT -195.560 -89.375 -195.390 -89.205 ;
        RECT -194.570 -89.375 -194.400 -89.205 ;
        RECT -185.640 -89.375 -185.470 -89.205 ;
        RECT -184.650 -89.375 -184.480 -89.205 ;
        RECT -175.720 -89.375 -175.550 -89.205 ;
        RECT -174.730 -89.375 -174.560 -89.205 ;
        RECT -165.800 -89.375 -165.630 -89.205 ;
        RECT -164.810 -89.375 -164.640 -89.205 ;
        RECT -155.880 -89.375 -155.710 -89.205 ;
        RECT -154.890 -89.375 -154.720 -89.205 ;
        RECT -145.960 -89.375 -145.790 -89.205 ;
        RECT -144.970 -89.375 -144.800 -89.205 ;
        RECT -136.040 -89.375 -135.870 -89.205 ;
        RECT -135.050 -89.375 -134.880 -89.205 ;
        RECT -126.120 -89.375 -125.950 -89.205 ;
        RECT -125.130 -89.375 -124.960 -89.205 ;
        RECT -116.200 -89.375 -116.030 -89.205 ;
        RECT -115.210 -89.375 -115.040 -89.205 ;
        RECT -106.280 -89.375 -106.110 -89.205 ;
        RECT -105.290 -89.375 -105.120 -89.205 ;
        RECT -96.360 -89.375 -96.190 -89.205 ;
        RECT -95.370 -89.375 -95.200 -89.205 ;
        RECT -86.440 -89.375 -86.270 -89.205 ;
        RECT -85.450 -89.375 -85.280 -89.205 ;
        RECT -76.520 -89.375 -76.350 -89.205 ;
        RECT -75.530 -89.375 -75.360 -89.205 ;
        RECT -66.600 -89.375 -66.430 -89.205 ;
        RECT -65.610 -89.375 -65.440 -89.205 ;
        RECT -56.680 -89.375 -56.510 -89.205 ;
        RECT -55.690 -89.375 -55.520 -89.205 ;
        RECT -46.760 -89.375 -46.590 -89.205 ;
        RECT -45.770 -89.375 -45.600 -89.205 ;
        RECT -36.840 -89.375 -36.670 -89.205 ;
        RECT -35.850 -89.375 -35.680 -89.205 ;
        RECT -26.920 -89.375 -26.750 -89.205 ;
        RECT -25.930 -89.375 -25.760 -89.205 ;
        RECT -17.000 -89.375 -16.830 -89.205 ;
        RECT -16.010 -89.375 -15.840 -89.205 ;
        RECT -7.080 -89.375 -6.910 -89.205 ;
        RECT -6.090 -89.375 -5.920 -89.205 ;
        RECT 2.840 -89.375 3.010 -89.205 ;
        RECT 3.830 -89.375 4.000 -89.205 ;
        RECT 12.760 -89.375 12.930 -89.205 ;
        RECT 13.750 -89.375 13.920 -89.205 ;
        RECT 22.680 -89.375 22.850 -89.205 ;
        RECT 23.670 -89.375 23.840 -89.205 ;
        RECT -288.560 -176.685 -288.390 -176.515 ;
        RECT -279.630 -176.685 -279.460 -176.515 ;
        RECT -278.640 -176.685 -278.470 -176.515 ;
        RECT -269.710 -176.685 -269.540 -176.515 ;
        RECT -268.720 -176.685 -268.550 -176.515 ;
        RECT -259.790 -176.685 -259.620 -176.515 ;
        RECT -258.800 -176.685 -258.630 -176.515 ;
        RECT -249.870 -176.685 -249.700 -176.515 ;
        RECT -248.880 -176.685 -248.710 -176.515 ;
        RECT -239.950 -176.685 -239.780 -176.515 ;
        RECT -238.960 -176.685 -238.790 -176.515 ;
        RECT -230.030 -176.685 -229.860 -176.515 ;
        RECT -229.040 -176.685 -228.870 -176.515 ;
        RECT -220.110 -176.685 -219.940 -176.515 ;
        RECT -219.120 -176.685 -218.950 -176.515 ;
        RECT -210.190 -176.685 -210.020 -176.515 ;
        RECT -209.200 -176.685 -209.030 -176.515 ;
        RECT -200.270 -176.685 -200.100 -176.515 ;
        RECT -199.280 -176.685 -199.110 -176.515 ;
        RECT -190.350 -176.685 -190.180 -176.515 ;
        RECT -189.360 -176.685 -189.190 -176.515 ;
        RECT -180.430 -176.685 -180.260 -176.515 ;
        RECT -179.440 -176.685 -179.270 -176.515 ;
        RECT -170.510 -176.685 -170.340 -176.515 ;
        RECT -169.520 -176.685 -169.350 -176.515 ;
        RECT -160.590 -176.685 -160.420 -176.515 ;
        RECT -159.600 -176.685 -159.430 -176.515 ;
        RECT -150.670 -176.685 -150.500 -176.515 ;
        RECT -149.680 -176.685 -149.510 -176.515 ;
        RECT -140.750 -176.685 -140.580 -176.515 ;
        RECT -139.760 -176.685 -139.590 -176.515 ;
        RECT -130.830 -176.685 -130.660 -176.515 ;
        RECT -129.840 -176.685 -129.670 -176.515 ;
        RECT -120.910 -176.685 -120.740 -176.515 ;
        RECT -119.920 -176.685 -119.750 -176.515 ;
        RECT -110.990 -176.685 -110.820 -176.515 ;
        RECT -110.000 -176.685 -109.830 -176.515 ;
        RECT -101.070 -176.685 -100.900 -176.515 ;
        RECT -100.080 -176.685 -99.910 -176.515 ;
        RECT -91.150 -176.685 -90.980 -176.515 ;
        RECT -90.160 -176.685 -89.990 -176.515 ;
        RECT -81.230 -176.685 -81.060 -176.515 ;
        RECT -80.240 -176.685 -80.070 -176.515 ;
        RECT -71.310 -176.685 -71.140 -176.515 ;
        RECT -70.320 -176.685 -70.150 -176.515 ;
        RECT -61.390 -176.685 -61.220 -176.515 ;
        RECT -60.400 -176.685 -60.230 -176.515 ;
        RECT -51.470 -176.685 -51.300 -176.515 ;
        RECT -50.480 -176.685 -50.310 -176.515 ;
        RECT -41.550 -176.685 -41.380 -176.515 ;
        RECT -40.560 -176.685 -40.390 -176.515 ;
        RECT -31.630 -176.685 -31.460 -176.515 ;
        RECT -30.640 -176.685 -30.470 -176.515 ;
        RECT -21.710 -176.685 -21.540 -176.515 ;
        RECT -20.720 -176.685 -20.550 -176.515 ;
        RECT -11.790 -176.685 -11.620 -176.515 ;
        RECT -10.800 -176.685 -10.630 -176.515 ;
        RECT -1.870 -176.685 -1.700 -176.515 ;
        RECT -0.880 -176.685 -0.710 -176.515 ;
        RECT 8.050 -176.685 8.220 -176.515 ;
        RECT 9.040 -176.685 9.210 -176.515 ;
        RECT 17.970 -176.685 18.140 -176.515 ;
        RECT 18.960 -176.685 19.130 -176.515 ;
        RECT 27.890 -176.685 28.060 -176.515 ;
        RECT -284.590 -177.085 -284.420 -176.915 ;
        RECT -283.600 -177.085 -283.430 -176.915 ;
        RECT -274.670 -177.085 -274.500 -176.915 ;
        RECT -273.680 -177.085 -273.510 -176.915 ;
        RECT -264.750 -177.085 -264.580 -176.915 ;
        RECT -263.760 -177.085 -263.590 -176.915 ;
        RECT -254.830 -177.085 -254.660 -176.915 ;
        RECT -253.840 -177.085 -253.670 -176.915 ;
        RECT -244.910 -177.085 -244.740 -176.915 ;
        RECT -243.920 -177.085 -243.750 -176.915 ;
        RECT -234.990 -177.085 -234.820 -176.915 ;
        RECT -234.000 -177.085 -233.830 -176.915 ;
        RECT -225.070 -177.085 -224.900 -176.915 ;
        RECT -224.080 -177.085 -223.910 -176.915 ;
        RECT -215.150 -177.085 -214.980 -176.915 ;
        RECT -214.160 -177.085 -213.990 -176.915 ;
        RECT -205.230 -177.085 -205.060 -176.915 ;
        RECT -204.240 -177.085 -204.070 -176.915 ;
        RECT -195.310 -177.085 -195.140 -176.915 ;
        RECT -194.320 -177.085 -194.150 -176.915 ;
        RECT -185.390 -177.085 -185.220 -176.915 ;
        RECT -184.400 -177.085 -184.230 -176.915 ;
        RECT -175.470 -177.085 -175.300 -176.915 ;
        RECT -174.480 -177.085 -174.310 -176.915 ;
        RECT -165.550 -177.085 -165.380 -176.915 ;
        RECT -164.560 -177.085 -164.390 -176.915 ;
        RECT -155.630 -177.085 -155.460 -176.915 ;
        RECT -154.640 -177.085 -154.470 -176.915 ;
        RECT -145.710 -177.085 -145.540 -176.915 ;
        RECT -144.720 -177.085 -144.550 -176.915 ;
        RECT -135.790 -177.085 -135.620 -176.915 ;
        RECT -134.800 -177.085 -134.630 -176.915 ;
        RECT -125.870 -177.085 -125.700 -176.915 ;
        RECT -124.880 -177.085 -124.710 -176.915 ;
        RECT -115.950 -177.085 -115.780 -176.915 ;
        RECT -114.960 -177.085 -114.790 -176.915 ;
        RECT -106.030 -177.085 -105.860 -176.915 ;
        RECT -105.040 -177.085 -104.870 -176.915 ;
        RECT -96.110 -177.085 -95.940 -176.915 ;
        RECT -95.120 -177.085 -94.950 -176.915 ;
        RECT -86.190 -177.085 -86.020 -176.915 ;
        RECT -85.200 -177.085 -85.030 -176.915 ;
        RECT -76.270 -177.085 -76.100 -176.915 ;
        RECT -75.280 -177.085 -75.110 -176.915 ;
        RECT -66.350 -177.085 -66.180 -176.915 ;
        RECT -65.360 -177.085 -65.190 -176.915 ;
        RECT -56.430 -177.085 -56.260 -176.915 ;
        RECT -55.440 -177.085 -55.270 -176.915 ;
        RECT -46.510 -177.085 -46.340 -176.915 ;
        RECT -45.520 -177.085 -45.350 -176.915 ;
        RECT -36.590 -177.085 -36.420 -176.915 ;
        RECT -35.600 -177.085 -35.430 -176.915 ;
        RECT -26.670 -177.085 -26.500 -176.915 ;
        RECT -25.680 -177.085 -25.510 -176.915 ;
        RECT -16.750 -177.085 -16.580 -176.915 ;
        RECT -15.760 -177.085 -15.590 -176.915 ;
        RECT -6.830 -177.085 -6.660 -176.915 ;
        RECT -5.840 -177.085 -5.670 -176.915 ;
        RECT 3.090 -177.085 3.260 -176.915 ;
        RECT 4.080 -177.085 4.250 -176.915 ;
        RECT 13.010 -177.085 13.180 -176.915 ;
        RECT 14.000 -177.085 14.170 -176.915 ;
        RECT 22.930 -177.085 23.100 -176.915 ;
        RECT 23.920 -177.085 24.090 -176.915 ;
      LAYER met1 ;
        RECT -291.010 91.900 -290.550 92.350 ;
        RECT -286.950 91.590 -286.490 92.040 ;
        RECT -286.050 91.590 -285.590 92.040 ;
        RECT -281.990 91.900 -281.530 92.350 ;
        RECT -281.090 91.900 -280.630 92.350 ;
        RECT -277.030 91.590 -276.570 92.040 ;
        RECT -276.130 91.590 -275.670 92.040 ;
        RECT -272.070 91.900 -271.610 92.350 ;
        RECT -271.170 91.900 -270.710 92.350 ;
        RECT -267.110 91.590 -266.650 92.040 ;
        RECT -266.210 91.590 -265.750 92.040 ;
        RECT -262.150 91.900 -261.690 92.350 ;
        RECT -261.250 91.900 -260.790 92.350 ;
        RECT -257.190 91.590 -256.730 92.040 ;
        RECT -256.290 91.590 -255.830 92.040 ;
        RECT -252.230 91.900 -251.770 92.350 ;
        RECT -251.330 91.900 -250.870 92.350 ;
        RECT -247.270 91.590 -246.810 92.040 ;
        RECT -246.370 91.590 -245.910 92.040 ;
        RECT -242.310 91.900 -241.850 92.350 ;
        RECT -241.410 91.900 -240.950 92.350 ;
        RECT -237.350 91.590 -236.890 92.040 ;
        RECT -236.450 91.590 -235.990 92.040 ;
        RECT -232.390 91.900 -231.930 92.350 ;
        RECT -231.490 91.900 -231.030 92.350 ;
        RECT -227.430 91.590 -226.970 92.040 ;
        RECT -226.530 91.590 -226.070 92.040 ;
        RECT -222.470 91.900 -222.010 92.350 ;
        RECT -221.570 91.900 -221.110 92.350 ;
        RECT -217.510 91.590 -217.050 92.040 ;
        RECT -216.610 91.590 -216.150 92.040 ;
        RECT -212.550 91.900 -212.090 92.350 ;
        RECT -211.650 91.900 -211.190 92.350 ;
        RECT -207.590 91.590 -207.130 92.040 ;
        RECT -206.690 91.590 -206.230 92.040 ;
        RECT -202.630 91.900 -202.170 92.350 ;
        RECT -201.730 91.900 -201.270 92.350 ;
        RECT -197.670 91.590 -197.210 92.040 ;
        RECT -196.770 91.590 -196.310 92.040 ;
        RECT -192.710 91.900 -192.250 92.350 ;
        RECT -191.810 91.900 -191.350 92.350 ;
        RECT -187.750 91.590 -187.290 92.040 ;
        RECT -186.850 91.590 -186.390 92.040 ;
        RECT -182.790 91.900 -182.330 92.350 ;
        RECT -181.890 91.900 -181.430 92.350 ;
        RECT -177.830 91.590 -177.370 92.040 ;
        RECT -176.930 91.590 -176.470 92.040 ;
        RECT -172.870 91.900 -172.410 92.350 ;
        RECT -171.970 91.900 -171.510 92.350 ;
        RECT -167.910 91.590 -167.450 92.040 ;
        RECT -167.010 91.590 -166.550 92.040 ;
        RECT -162.950 91.900 -162.490 92.350 ;
        RECT -162.050 91.900 -161.590 92.350 ;
        RECT -157.990 91.590 -157.530 92.040 ;
        RECT -157.090 91.590 -156.630 92.040 ;
        RECT -153.030 91.900 -152.570 92.350 ;
        RECT -152.130 91.900 -151.670 92.350 ;
        RECT -148.070 91.590 -147.610 92.040 ;
        RECT -147.170 91.590 -146.710 92.040 ;
        RECT -143.110 91.900 -142.650 92.350 ;
        RECT -142.210 91.900 -141.750 92.350 ;
        RECT -138.150 91.590 -137.690 92.040 ;
        RECT -137.250 91.590 -136.790 92.040 ;
        RECT -133.190 91.900 -132.730 92.350 ;
        RECT -132.290 91.900 -131.830 92.350 ;
        RECT -128.230 91.590 -127.770 92.040 ;
        RECT -127.330 91.590 -126.870 92.040 ;
        RECT -123.270 91.900 -122.810 92.350 ;
        RECT -122.370 91.900 -121.910 92.350 ;
        RECT -118.310 91.590 -117.850 92.040 ;
        RECT -117.410 91.590 -116.950 92.040 ;
        RECT -113.350 91.900 -112.890 92.350 ;
        RECT -112.450 91.900 -111.990 92.350 ;
        RECT -108.390 91.590 -107.930 92.040 ;
        RECT -107.490 91.590 -107.030 92.040 ;
        RECT -103.430 91.900 -102.970 92.350 ;
        RECT -102.530 91.900 -102.070 92.350 ;
        RECT -98.470 91.590 -98.010 92.040 ;
        RECT -97.570 91.590 -97.110 92.040 ;
        RECT -93.510 91.900 -93.050 92.350 ;
        RECT -92.610 91.900 -92.150 92.350 ;
        RECT -88.550 91.590 -88.090 92.040 ;
        RECT -87.650 91.590 -87.190 92.040 ;
        RECT -83.590 91.900 -83.130 92.350 ;
        RECT -82.690 91.900 -82.230 92.350 ;
        RECT -78.630 91.590 -78.170 92.040 ;
        RECT -77.730 91.590 -77.270 92.040 ;
        RECT -73.670 91.900 -73.210 92.350 ;
        RECT -72.770 91.900 -72.310 92.350 ;
        RECT -68.710 91.590 -68.250 92.040 ;
        RECT -67.810 91.590 -67.350 92.040 ;
        RECT -63.750 91.900 -63.290 92.350 ;
        RECT -62.850 91.900 -62.390 92.350 ;
        RECT -58.790 91.590 -58.330 92.040 ;
        RECT -57.890 91.590 -57.430 92.040 ;
        RECT -53.830 91.900 -53.370 92.350 ;
        RECT -52.930 91.900 -52.470 92.350 ;
        RECT -48.870 91.590 -48.410 92.040 ;
        RECT -47.970 91.590 -47.510 92.040 ;
        RECT -43.910 91.900 -43.450 92.350 ;
        RECT -43.010 91.900 -42.550 92.350 ;
        RECT -38.950 91.590 -38.490 92.040 ;
        RECT -38.050 91.590 -37.590 92.040 ;
        RECT -33.990 91.900 -33.530 92.350 ;
        RECT -33.090 91.900 -32.630 92.350 ;
        RECT -29.030 91.590 -28.570 92.040 ;
        RECT -28.130 91.590 -27.670 92.040 ;
        RECT -24.070 91.900 -23.610 92.350 ;
        RECT -23.170 91.900 -22.710 92.350 ;
        RECT -19.110 91.590 -18.650 92.040 ;
        RECT -18.210 91.590 -17.750 92.040 ;
        RECT -14.150 91.900 -13.690 92.350 ;
        RECT -13.250 91.900 -12.790 92.350 ;
        RECT -9.190 91.590 -8.730 92.040 ;
        RECT -8.290 91.590 -7.830 92.040 ;
        RECT -4.230 91.900 -3.770 92.350 ;
        RECT -3.330 91.900 -2.870 92.350 ;
        RECT 0.730 91.590 1.190 92.040 ;
        RECT 1.630 91.590 2.090 92.040 ;
        RECT 5.690 91.900 6.150 92.350 ;
        RECT 6.590 91.900 7.050 92.350 ;
        RECT 10.650 91.590 11.110 92.040 ;
        RECT 11.550 91.590 12.010 92.040 ;
        RECT 15.610 91.900 16.070 92.350 ;
        RECT 16.510 91.900 16.970 92.350 ;
        RECT 20.570 91.590 21.030 92.040 ;
        RECT 21.470 91.590 21.930 92.040 ;
        RECT 25.530 91.900 25.990 92.350 ;
        RECT -290.760 4.190 -290.300 4.640 ;
        RECT -286.700 3.880 -286.240 4.330 ;
        RECT -285.800 3.880 -285.340 4.330 ;
        RECT -281.740 4.190 -281.280 4.640 ;
        RECT -280.840 4.190 -280.380 4.640 ;
        RECT -276.780 3.880 -276.320 4.330 ;
        RECT -275.880 3.880 -275.420 4.330 ;
        RECT -271.820 4.190 -271.360 4.640 ;
        RECT -270.920 4.190 -270.460 4.640 ;
        RECT -266.860 3.880 -266.400 4.330 ;
        RECT -265.960 3.880 -265.500 4.330 ;
        RECT -261.900 4.190 -261.440 4.640 ;
        RECT -261.000 4.190 -260.540 4.640 ;
        RECT -256.940 3.880 -256.480 4.330 ;
        RECT -256.040 3.880 -255.580 4.330 ;
        RECT -251.980 4.190 -251.520 4.640 ;
        RECT -251.080 4.190 -250.620 4.640 ;
        RECT -247.020 3.880 -246.560 4.330 ;
        RECT -246.120 3.880 -245.660 4.330 ;
        RECT -242.060 4.190 -241.600 4.640 ;
        RECT -241.160 4.190 -240.700 4.640 ;
        RECT -237.100 3.880 -236.640 4.330 ;
        RECT -236.200 3.880 -235.740 4.330 ;
        RECT -232.140 4.190 -231.680 4.640 ;
        RECT -231.240 4.190 -230.780 4.640 ;
        RECT -227.180 3.880 -226.720 4.330 ;
        RECT -226.280 3.880 -225.820 4.330 ;
        RECT -222.220 4.190 -221.760 4.640 ;
        RECT -221.320 4.190 -220.860 4.640 ;
        RECT -217.260 3.880 -216.800 4.330 ;
        RECT -216.360 3.880 -215.900 4.330 ;
        RECT -212.300 4.190 -211.840 4.640 ;
        RECT -211.400 4.190 -210.940 4.640 ;
        RECT -207.340 3.880 -206.880 4.330 ;
        RECT -206.440 3.880 -205.980 4.330 ;
        RECT -202.380 4.190 -201.920 4.640 ;
        RECT -201.480 4.190 -201.020 4.640 ;
        RECT -197.420 3.880 -196.960 4.330 ;
        RECT -196.520 3.880 -196.060 4.330 ;
        RECT -192.460 4.190 -192.000 4.640 ;
        RECT -191.560 4.190 -191.100 4.640 ;
        RECT -187.500 3.880 -187.040 4.330 ;
        RECT -186.600 3.880 -186.140 4.330 ;
        RECT -182.540 4.190 -182.080 4.640 ;
        RECT -181.640 4.190 -181.180 4.640 ;
        RECT -177.580 3.880 -177.120 4.330 ;
        RECT -176.680 3.880 -176.220 4.330 ;
        RECT -172.620 4.190 -172.160 4.640 ;
        RECT -171.720 4.190 -171.260 4.640 ;
        RECT -167.660 3.880 -167.200 4.330 ;
        RECT -166.760 3.880 -166.300 4.330 ;
        RECT -162.700 4.190 -162.240 4.640 ;
        RECT -161.800 4.190 -161.340 4.640 ;
        RECT -157.740 3.880 -157.280 4.330 ;
        RECT -156.840 3.880 -156.380 4.330 ;
        RECT -152.780 4.190 -152.320 4.640 ;
        RECT -151.880 4.190 -151.420 4.640 ;
        RECT -147.820 3.880 -147.360 4.330 ;
        RECT -146.920 3.880 -146.460 4.330 ;
        RECT -142.860 4.190 -142.400 4.640 ;
        RECT -141.960 4.190 -141.500 4.640 ;
        RECT -137.900 3.880 -137.440 4.330 ;
        RECT -137.000 3.880 -136.540 4.330 ;
        RECT -132.940 4.190 -132.480 4.640 ;
        RECT -132.040 4.190 -131.580 4.640 ;
        RECT -127.980 3.880 -127.520 4.330 ;
        RECT -127.080 3.880 -126.620 4.330 ;
        RECT -123.020 4.190 -122.560 4.640 ;
        RECT -122.120 4.190 -121.660 4.640 ;
        RECT -118.060 3.880 -117.600 4.330 ;
        RECT -117.160 3.880 -116.700 4.330 ;
        RECT -113.100 4.190 -112.640 4.640 ;
        RECT -112.200 4.190 -111.740 4.640 ;
        RECT -108.140 3.880 -107.680 4.330 ;
        RECT -107.240 3.880 -106.780 4.330 ;
        RECT -103.180 4.190 -102.720 4.640 ;
        RECT -102.280 4.190 -101.820 4.640 ;
        RECT -98.220 3.880 -97.760 4.330 ;
        RECT -97.320 3.880 -96.860 4.330 ;
        RECT -93.260 4.190 -92.800 4.640 ;
        RECT -92.360 4.190 -91.900 4.640 ;
        RECT -88.300 3.880 -87.840 4.330 ;
        RECT -87.400 3.880 -86.940 4.330 ;
        RECT -83.340 4.190 -82.880 4.640 ;
        RECT -82.440 4.190 -81.980 4.640 ;
        RECT -78.380 3.880 -77.920 4.330 ;
        RECT -77.480 3.880 -77.020 4.330 ;
        RECT -73.420 4.190 -72.960 4.640 ;
        RECT -72.520 4.190 -72.060 4.640 ;
        RECT -68.460 3.880 -68.000 4.330 ;
        RECT -67.560 3.880 -67.100 4.330 ;
        RECT -63.500 4.190 -63.040 4.640 ;
        RECT -62.600 4.190 -62.140 4.640 ;
        RECT -58.540 3.880 -58.080 4.330 ;
        RECT -57.640 3.880 -57.180 4.330 ;
        RECT -53.580 4.190 -53.120 4.640 ;
        RECT -52.680 4.190 -52.220 4.640 ;
        RECT -48.620 3.880 -48.160 4.330 ;
        RECT -47.720 3.880 -47.260 4.330 ;
        RECT -43.660 4.190 -43.200 4.640 ;
        RECT -42.760 4.190 -42.300 4.640 ;
        RECT -38.700 3.880 -38.240 4.330 ;
        RECT -37.800 3.880 -37.340 4.330 ;
        RECT -33.740 4.190 -33.280 4.640 ;
        RECT -32.840 4.190 -32.380 4.640 ;
        RECT -28.780 3.880 -28.320 4.330 ;
        RECT -27.880 3.880 -27.420 4.330 ;
        RECT -23.820 4.190 -23.360 4.640 ;
        RECT -22.920 4.190 -22.460 4.640 ;
        RECT -18.860 3.880 -18.400 4.330 ;
        RECT -17.960 3.880 -17.500 4.330 ;
        RECT -13.900 4.190 -13.440 4.640 ;
        RECT -13.000 4.190 -12.540 4.640 ;
        RECT -8.940 3.880 -8.480 4.330 ;
        RECT -8.040 3.880 -7.580 4.330 ;
        RECT -3.980 4.190 -3.520 4.640 ;
        RECT -3.080 4.190 -2.620 4.640 ;
        RECT 0.980 3.880 1.440 4.330 ;
        RECT 1.880 3.880 2.340 4.330 ;
        RECT 5.940 4.190 6.400 4.640 ;
        RECT 6.840 4.190 7.300 4.640 ;
        RECT 10.900 3.880 11.360 4.330 ;
        RECT 11.800 3.880 12.260 4.330 ;
        RECT 15.860 4.190 16.320 4.640 ;
        RECT 16.760 4.190 17.220 4.640 ;
        RECT 20.820 3.880 21.280 4.330 ;
        RECT 21.720 3.880 22.180 4.330 ;
        RECT 25.780 4.190 26.240 4.640 ;
        RECT -289.000 -89.160 -288.540 -88.710 ;
        RECT -284.940 -89.470 -284.480 -89.020 ;
        RECT -284.040 -89.470 -283.580 -89.020 ;
        RECT -279.980 -89.160 -279.520 -88.710 ;
        RECT -279.080 -89.160 -278.620 -88.710 ;
        RECT -275.020 -89.470 -274.560 -89.020 ;
        RECT -274.120 -89.470 -273.660 -89.020 ;
        RECT -270.060 -89.160 -269.600 -88.710 ;
        RECT -269.160 -89.160 -268.700 -88.710 ;
        RECT -265.100 -89.470 -264.640 -89.020 ;
        RECT -264.200 -89.470 -263.740 -89.020 ;
        RECT -260.140 -89.160 -259.680 -88.710 ;
        RECT -259.240 -89.160 -258.780 -88.710 ;
        RECT -255.180 -89.470 -254.720 -89.020 ;
        RECT -254.280 -89.470 -253.820 -89.020 ;
        RECT -250.220 -89.160 -249.760 -88.710 ;
        RECT -249.320 -89.160 -248.860 -88.710 ;
        RECT -245.260 -89.470 -244.800 -89.020 ;
        RECT -244.360 -89.470 -243.900 -89.020 ;
        RECT -240.300 -89.160 -239.840 -88.710 ;
        RECT -239.400 -89.160 -238.940 -88.710 ;
        RECT -235.340 -89.470 -234.880 -89.020 ;
        RECT -234.440 -89.470 -233.980 -89.020 ;
        RECT -230.380 -89.160 -229.920 -88.710 ;
        RECT -229.480 -89.160 -229.020 -88.710 ;
        RECT -225.420 -89.470 -224.960 -89.020 ;
        RECT -224.520 -89.470 -224.060 -89.020 ;
        RECT -220.460 -89.160 -220.000 -88.710 ;
        RECT -219.560 -89.160 -219.100 -88.710 ;
        RECT -215.500 -89.470 -215.040 -89.020 ;
        RECT -214.600 -89.470 -214.140 -89.020 ;
        RECT -210.540 -89.160 -210.080 -88.710 ;
        RECT -209.640 -89.160 -209.180 -88.710 ;
        RECT -205.580 -89.470 -205.120 -89.020 ;
        RECT -204.680 -89.470 -204.220 -89.020 ;
        RECT -200.620 -89.160 -200.160 -88.710 ;
        RECT -199.720 -89.160 -199.260 -88.710 ;
        RECT -195.660 -89.470 -195.200 -89.020 ;
        RECT -194.760 -89.470 -194.300 -89.020 ;
        RECT -190.700 -89.160 -190.240 -88.710 ;
        RECT -189.800 -89.160 -189.340 -88.710 ;
        RECT -185.740 -89.470 -185.280 -89.020 ;
        RECT -184.840 -89.470 -184.380 -89.020 ;
        RECT -180.780 -89.160 -180.320 -88.710 ;
        RECT -179.880 -89.160 -179.420 -88.710 ;
        RECT -175.820 -89.470 -175.360 -89.020 ;
        RECT -174.920 -89.470 -174.460 -89.020 ;
        RECT -170.860 -89.160 -170.400 -88.710 ;
        RECT -169.960 -89.160 -169.500 -88.710 ;
        RECT -165.900 -89.470 -165.440 -89.020 ;
        RECT -165.000 -89.470 -164.540 -89.020 ;
        RECT -160.940 -89.160 -160.480 -88.710 ;
        RECT -160.040 -89.160 -159.580 -88.710 ;
        RECT -155.980 -89.470 -155.520 -89.020 ;
        RECT -155.080 -89.470 -154.620 -89.020 ;
        RECT -151.020 -89.160 -150.560 -88.710 ;
        RECT -150.120 -89.160 -149.660 -88.710 ;
        RECT -146.060 -89.470 -145.600 -89.020 ;
        RECT -145.160 -89.470 -144.700 -89.020 ;
        RECT -141.100 -89.160 -140.640 -88.710 ;
        RECT -140.200 -89.160 -139.740 -88.710 ;
        RECT -136.140 -89.470 -135.680 -89.020 ;
        RECT -135.240 -89.470 -134.780 -89.020 ;
        RECT -131.180 -89.160 -130.720 -88.710 ;
        RECT -130.280 -89.160 -129.820 -88.710 ;
        RECT -126.220 -89.470 -125.760 -89.020 ;
        RECT -125.320 -89.470 -124.860 -89.020 ;
        RECT -121.260 -89.160 -120.800 -88.710 ;
        RECT -120.360 -89.160 -119.900 -88.710 ;
        RECT -116.300 -89.470 -115.840 -89.020 ;
        RECT -115.400 -89.470 -114.940 -89.020 ;
        RECT -111.340 -89.160 -110.880 -88.710 ;
        RECT -110.440 -89.160 -109.980 -88.710 ;
        RECT -106.380 -89.470 -105.920 -89.020 ;
        RECT -105.480 -89.470 -105.020 -89.020 ;
        RECT -101.420 -89.160 -100.960 -88.710 ;
        RECT -100.520 -89.160 -100.060 -88.710 ;
        RECT -96.460 -89.470 -96.000 -89.020 ;
        RECT -95.560 -89.470 -95.100 -89.020 ;
        RECT -91.500 -89.160 -91.040 -88.710 ;
        RECT -90.600 -89.160 -90.140 -88.710 ;
        RECT -86.540 -89.470 -86.080 -89.020 ;
        RECT -85.640 -89.470 -85.180 -89.020 ;
        RECT -81.580 -89.160 -81.120 -88.710 ;
        RECT -80.680 -89.160 -80.220 -88.710 ;
        RECT -76.620 -89.470 -76.160 -89.020 ;
        RECT -75.720 -89.470 -75.260 -89.020 ;
        RECT -71.660 -89.160 -71.200 -88.710 ;
        RECT -70.760 -89.160 -70.300 -88.710 ;
        RECT -66.700 -89.470 -66.240 -89.020 ;
        RECT -65.800 -89.470 -65.340 -89.020 ;
        RECT -61.740 -89.160 -61.280 -88.710 ;
        RECT -60.840 -89.160 -60.380 -88.710 ;
        RECT -56.780 -89.470 -56.320 -89.020 ;
        RECT -55.880 -89.470 -55.420 -89.020 ;
        RECT -51.820 -89.160 -51.360 -88.710 ;
        RECT -50.920 -89.160 -50.460 -88.710 ;
        RECT -46.860 -89.470 -46.400 -89.020 ;
        RECT -45.960 -89.470 -45.500 -89.020 ;
        RECT -41.900 -89.160 -41.440 -88.710 ;
        RECT -41.000 -89.160 -40.540 -88.710 ;
        RECT -36.940 -89.470 -36.480 -89.020 ;
        RECT -36.040 -89.470 -35.580 -89.020 ;
        RECT -31.980 -89.160 -31.520 -88.710 ;
        RECT -31.080 -89.160 -30.620 -88.710 ;
        RECT -27.020 -89.470 -26.560 -89.020 ;
        RECT -26.120 -89.470 -25.660 -89.020 ;
        RECT -22.060 -89.160 -21.600 -88.710 ;
        RECT -21.160 -89.160 -20.700 -88.710 ;
        RECT -17.100 -89.470 -16.640 -89.020 ;
        RECT -16.200 -89.470 -15.740 -89.020 ;
        RECT -12.140 -89.160 -11.680 -88.710 ;
        RECT -11.240 -89.160 -10.780 -88.710 ;
        RECT -7.180 -89.470 -6.720 -89.020 ;
        RECT -6.280 -89.470 -5.820 -89.020 ;
        RECT -2.220 -89.160 -1.760 -88.710 ;
        RECT -1.320 -89.160 -0.860 -88.710 ;
        RECT 2.740 -89.470 3.200 -89.020 ;
        RECT 3.640 -89.470 4.100 -89.020 ;
        RECT 7.700 -89.160 8.160 -88.710 ;
        RECT 8.600 -89.160 9.060 -88.710 ;
        RECT 12.660 -89.470 13.120 -89.020 ;
        RECT 13.560 -89.470 14.020 -89.020 ;
        RECT 17.620 -89.160 18.080 -88.710 ;
        RECT 18.520 -89.160 18.980 -88.710 ;
        RECT 22.580 -89.470 23.040 -89.020 ;
        RECT 23.480 -89.470 23.940 -89.020 ;
        RECT 27.540 -89.160 28.000 -88.710 ;
        RECT -288.750 -176.870 -288.290 -176.420 ;
        RECT -284.690 -177.180 -284.230 -176.730 ;
        RECT -283.790 -177.180 -283.330 -176.730 ;
        RECT -279.730 -176.870 -279.270 -176.420 ;
        RECT -278.830 -176.870 -278.370 -176.420 ;
        RECT -274.770 -177.180 -274.310 -176.730 ;
        RECT -273.870 -177.180 -273.410 -176.730 ;
        RECT -269.810 -176.870 -269.350 -176.420 ;
        RECT -268.910 -176.870 -268.450 -176.420 ;
        RECT -264.850 -177.180 -264.390 -176.730 ;
        RECT -263.950 -177.180 -263.490 -176.730 ;
        RECT -259.890 -176.870 -259.430 -176.420 ;
        RECT -258.990 -176.870 -258.530 -176.420 ;
        RECT -254.930 -177.180 -254.470 -176.730 ;
        RECT -254.030 -177.180 -253.570 -176.730 ;
        RECT -249.970 -176.870 -249.510 -176.420 ;
        RECT -249.070 -176.870 -248.610 -176.420 ;
        RECT -245.010 -177.180 -244.550 -176.730 ;
        RECT -244.110 -177.180 -243.650 -176.730 ;
        RECT -240.050 -176.870 -239.590 -176.420 ;
        RECT -239.150 -176.870 -238.690 -176.420 ;
        RECT -235.090 -177.180 -234.630 -176.730 ;
        RECT -234.190 -177.180 -233.730 -176.730 ;
        RECT -230.130 -176.870 -229.670 -176.420 ;
        RECT -229.230 -176.870 -228.770 -176.420 ;
        RECT -225.170 -177.180 -224.710 -176.730 ;
        RECT -224.270 -177.180 -223.810 -176.730 ;
        RECT -220.210 -176.870 -219.750 -176.420 ;
        RECT -219.310 -176.870 -218.850 -176.420 ;
        RECT -215.250 -177.180 -214.790 -176.730 ;
        RECT -214.350 -177.180 -213.890 -176.730 ;
        RECT -210.290 -176.870 -209.830 -176.420 ;
        RECT -209.390 -176.870 -208.930 -176.420 ;
        RECT -205.330 -177.180 -204.870 -176.730 ;
        RECT -204.430 -177.180 -203.970 -176.730 ;
        RECT -200.370 -176.870 -199.910 -176.420 ;
        RECT -199.470 -176.870 -199.010 -176.420 ;
        RECT -195.410 -177.180 -194.950 -176.730 ;
        RECT -194.510 -177.180 -194.050 -176.730 ;
        RECT -190.450 -176.870 -189.990 -176.420 ;
        RECT -189.550 -176.870 -189.090 -176.420 ;
        RECT -185.490 -177.180 -185.030 -176.730 ;
        RECT -184.590 -177.180 -184.130 -176.730 ;
        RECT -180.530 -176.870 -180.070 -176.420 ;
        RECT -179.630 -176.870 -179.170 -176.420 ;
        RECT -175.570 -177.180 -175.110 -176.730 ;
        RECT -174.670 -177.180 -174.210 -176.730 ;
        RECT -170.610 -176.870 -170.150 -176.420 ;
        RECT -169.710 -176.870 -169.250 -176.420 ;
        RECT -165.650 -177.180 -165.190 -176.730 ;
        RECT -164.750 -177.180 -164.290 -176.730 ;
        RECT -160.690 -176.870 -160.230 -176.420 ;
        RECT -159.790 -176.870 -159.330 -176.420 ;
        RECT -155.730 -177.180 -155.270 -176.730 ;
        RECT -154.830 -177.180 -154.370 -176.730 ;
        RECT -150.770 -176.870 -150.310 -176.420 ;
        RECT -149.870 -176.870 -149.410 -176.420 ;
        RECT -145.810 -177.180 -145.350 -176.730 ;
        RECT -144.910 -177.180 -144.450 -176.730 ;
        RECT -140.850 -176.870 -140.390 -176.420 ;
        RECT -139.950 -176.870 -139.490 -176.420 ;
        RECT -135.890 -177.180 -135.430 -176.730 ;
        RECT -134.990 -177.180 -134.530 -176.730 ;
        RECT -130.930 -176.870 -130.470 -176.420 ;
        RECT -130.030 -176.870 -129.570 -176.420 ;
        RECT -125.970 -177.180 -125.510 -176.730 ;
        RECT -125.070 -177.180 -124.610 -176.730 ;
        RECT -121.010 -176.870 -120.550 -176.420 ;
        RECT -120.110 -176.870 -119.650 -176.420 ;
        RECT -116.050 -177.180 -115.590 -176.730 ;
        RECT -115.150 -177.180 -114.690 -176.730 ;
        RECT -111.090 -176.870 -110.630 -176.420 ;
        RECT -110.190 -176.870 -109.730 -176.420 ;
        RECT -106.130 -177.180 -105.670 -176.730 ;
        RECT -105.230 -177.180 -104.770 -176.730 ;
        RECT -101.170 -176.870 -100.710 -176.420 ;
        RECT -100.270 -176.870 -99.810 -176.420 ;
        RECT -96.210 -177.180 -95.750 -176.730 ;
        RECT -95.310 -177.180 -94.850 -176.730 ;
        RECT -91.250 -176.870 -90.790 -176.420 ;
        RECT -90.350 -176.870 -89.890 -176.420 ;
        RECT -86.290 -177.180 -85.830 -176.730 ;
        RECT -85.390 -177.180 -84.930 -176.730 ;
        RECT -81.330 -176.870 -80.870 -176.420 ;
        RECT -80.430 -176.870 -79.970 -176.420 ;
        RECT -76.370 -177.180 -75.910 -176.730 ;
        RECT -75.470 -177.180 -75.010 -176.730 ;
        RECT -71.410 -176.870 -70.950 -176.420 ;
        RECT -70.510 -176.870 -70.050 -176.420 ;
        RECT -66.450 -177.180 -65.990 -176.730 ;
        RECT -65.550 -177.180 -65.090 -176.730 ;
        RECT -61.490 -176.870 -61.030 -176.420 ;
        RECT -60.590 -176.870 -60.130 -176.420 ;
        RECT -56.530 -177.180 -56.070 -176.730 ;
        RECT -55.630 -177.180 -55.170 -176.730 ;
        RECT -51.570 -176.870 -51.110 -176.420 ;
        RECT -50.670 -176.870 -50.210 -176.420 ;
        RECT -46.610 -177.180 -46.150 -176.730 ;
        RECT -45.710 -177.180 -45.250 -176.730 ;
        RECT -41.650 -176.870 -41.190 -176.420 ;
        RECT -40.750 -176.870 -40.290 -176.420 ;
        RECT -36.690 -177.180 -36.230 -176.730 ;
        RECT -35.790 -177.180 -35.330 -176.730 ;
        RECT -31.730 -176.870 -31.270 -176.420 ;
        RECT -30.830 -176.870 -30.370 -176.420 ;
        RECT -26.770 -177.180 -26.310 -176.730 ;
        RECT -25.870 -177.180 -25.410 -176.730 ;
        RECT -21.810 -176.870 -21.350 -176.420 ;
        RECT -20.910 -176.870 -20.450 -176.420 ;
        RECT -16.850 -177.180 -16.390 -176.730 ;
        RECT -15.950 -177.180 -15.490 -176.730 ;
        RECT -11.890 -176.870 -11.430 -176.420 ;
        RECT -10.990 -176.870 -10.530 -176.420 ;
        RECT -6.930 -177.180 -6.470 -176.730 ;
        RECT -6.030 -177.180 -5.570 -176.730 ;
        RECT -1.970 -176.870 -1.510 -176.420 ;
        RECT -1.070 -176.870 -0.610 -176.420 ;
        RECT 2.990 -177.180 3.450 -176.730 ;
        RECT 3.890 -177.180 4.350 -176.730 ;
        RECT 7.950 -176.870 8.410 -176.420 ;
        RECT 8.850 -176.870 9.310 -176.420 ;
        RECT 12.910 -177.180 13.370 -176.730 ;
        RECT 13.810 -177.180 14.270 -176.730 ;
        RECT 17.870 -176.870 18.330 -176.420 ;
        RECT 18.770 -176.870 19.230 -176.420 ;
        RECT 22.830 -177.180 23.290 -176.730 ;
        RECT 23.730 -177.180 24.190 -176.730 ;
        RECT 27.790 -176.870 28.250 -176.420 ;
      LAYER via ;
        RECT -290.920 92.020 -290.660 92.280 ;
        RECT -286.840 91.660 -286.580 91.920 ;
        RECT -285.960 91.660 -285.700 91.920 ;
        RECT -281.880 92.020 -281.620 92.280 ;
        RECT -281.000 92.020 -280.740 92.280 ;
        RECT -276.920 91.660 -276.660 91.920 ;
        RECT -276.040 91.660 -275.780 91.920 ;
        RECT -271.960 92.020 -271.700 92.280 ;
        RECT -271.080 92.020 -270.820 92.280 ;
        RECT -267.000 91.660 -266.740 91.920 ;
        RECT -266.120 91.660 -265.860 91.920 ;
        RECT -262.040 92.020 -261.780 92.280 ;
        RECT -261.160 92.020 -260.900 92.280 ;
        RECT -257.080 91.660 -256.820 91.920 ;
        RECT -256.200 91.660 -255.940 91.920 ;
        RECT -252.120 92.020 -251.860 92.280 ;
        RECT -251.240 92.020 -250.980 92.280 ;
        RECT -247.160 91.660 -246.900 91.920 ;
        RECT -246.280 91.660 -246.020 91.920 ;
        RECT -242.200 92.020 -241.940 92.280 ;
        RECT -241.320 92.020 -241.060 92.280 ;
        RECT -237.240 91.660 -236.980 91.920 ;
        RECT -236.360 91.660 -236.100 91.920 ;
        RECT -232.280 92.020 -232.020 92.280 ;
        RECT -231.400 92.020 -231.140 92.280 ;
        RECT -227.320 91.660 -227.060 91.920 ;
        RECT -226.440 91.660 -226.180 91.920 ;
        RECT -222.360 92.020 -222.100 92.280 ;
        RECT -221.480 92.020 -221.220 92.280 ;
        RECT -217.400 91.660 -217.140 91.920 ;
        RECT -216.520 91.660 -216.260 91.920 ;
        RECT -212.440 92.020 -212.180 92.280 ;
        RECT -211.560 92.020 -211.300 92.280 ;
        RECT -207.480 91.660 -207.220 91.920 ;
        RECT -206.600 91.660 -206.340 91.920 ;
        RECT -202.520 92.020 -202.260 92.280 ;
        RECT -201.640 92.020 -201.380 92.280 ;
        RECT -197.560 91.660 -197.300 91.920 ;
        RECT -196.680 91.660 -196.420 91.920 ;
        RECT -192.600 92.020 -192.340 92.280 ;
        RECT -191.720 92.020 -191.460 92.280 ;
        RECT -187.640 91.660 -187.380 91.920 ;
        RECT -186.760 91.660 -186.500 91.920 ;
        RECT -182.680 92.020 -182.420 92.280 ;
        RECT -181.800 92.020 -181.540 92.280 ;
        RECT -177.720 91.660 -177.460 91.920 ;
        RECT -176.840 91.660 -176.580 91.920 ;
        RECT -172.760 92.020 -172.500 92.280 ;
        RECT -171.880 92.020 -171.620 92.280 ;
        RECT -167.800 91.660 -167.540 91.920 ;
        RECT -166.920 91.660 -166.660 91.920 ;
        RECT -162.840 92.020 -162.580 92.280 ;
        RECT -161.960 92.020 -161.700 92.280 ;
        RECT -157.880 91.660 -157.620 91.920 ;
        RECT -157.000 91.660 -156.740 91.920 ;
        RECT -152.920 92.020 -152.660 92.280 ;
        RECT -152.040 92.020 -151.780 92.280 ;
        RECT -147.960 91.660 -147.700 91.920 ;
        RECT -147.080 91.660 -146.820 91.920 ;
        RECT -143.000 92.020 -142.740 92.280 ;
        RECT -142.120 92.020 -141.860 92.280 ;
        RECT -138.040 91.660 -137.780 91.920 ;
        RECT -137.160 91.660 -136.900 91.920 ;
        RECT -133.080 92.020 -132.820 92.280 ;
        RECT -132.200 92.020 -131.940 92.280 ;
        RECT -128.120 91.660 -127.860 91.920 ;
        RECT -127.240 91.660 -126.980 91.920 ;
        RECT -123.160 92.020 -122.900 92.280 ;
        RECT -122.280 92.020 -122.020 92.280 ;
        RECT -118.200 91.660 -117.940 91.920 ;
        RECT -117.320 91.660 -117.060 91.920 ;
        RECT -113.240 92.020 -112.980 92.280 ;
        RECT -112.360 92.020 -112.100 92.280 ;
        RECT -108.280 91.660 -108.020 91.920 ;
        RECT -107.400 91.660 -107.140 91.920 ;
        RECT -103.320 92.020 -103.060 92.280 ;
        RECT -102.440 92.020 -102.180 92.280 ;
        RECT -98.360 91.660 -98.100 91.920 ;
        RECT -97.480 91.660 -97.220 91.920 ;
        RECT -93.400 92.020 -93.140 92.280 ;
        RECT -92.520 92.020 -92.260 92.280 ;
        RECT -88.440 91.660 -88.180 91.920 ;
        RECT -87.560 91.660 -87.300 91.920 ;
        RECT -83.480 92.020 -83.220 92.280 ;
        RECT -82.600 92.020 -82.340 92.280 ;
        RECT -78.520 91.660 -78.260 91.920 ;
        RECT -77.640 91.660 -77.380 91.920 ;
        RECT -73.560 92.020 -73.300 92.280 ;
        RECT -72.680 92.020 -72.420 92.280 ;
        RECT -68.600 91.660 -68.340 91.920 ;
        RECT -67.720 91.660 -67.460 91.920 ;
        RECT -63.640 92.020 -63.380 92.280 ;
        RECT -62.760 92.020 -62.500 92.280 ;
        RECT -58.680 91.660 -58.420 91.920 ;
        RECT -57.800 91.660 -57.540 91.920 ;
        RECT -53.720 92.020 -53.460 92.280 ;
        RECT -52.840 92.020 -52.580 92.280 ;
        RECT -48.760 91.660 -48.500 91.920 ;
        RECT -47.880 91.660 -47.620 91.920 ;
        RECT -43.800 92.020 -43.540 92.280 ;
        RECT -42.920 92.020 -42.660 92.280 ;
        RECT -38.840 91.660 -38.580 91.920 ;
        RECT -37.960 91.660 -37.700 91.920 ;
        RECT -33.880 92.020 -33.620 92.280 ;
        RECT -33.000 92.020 -32.740 92.280 ;
        RECT -28.920 91.660 -28.660 91.920 ;
        RECT -28.040 91.660 -27.780 91.920 ;
        RECT -23.960 92.020 -23.700 92.280 ;
        RECT -23.080 92.020 -22.820 92.280 ;
        RECT -19.000 91.660 -18.740 91.920 ;
        RECT -18.120 91.660 -17.860 91.920 ;
        RECT -14.040 92.020 -13.780 92.280 ;
        RECT -13.160 92.020 -12.900 92.280 ;
        RECT -9.080 91.660 -8.820 91.920 ;
        RECT -8.200 91.660 -7.940 91.920 ;
        RECT -4.120 92.020 -3.860 92.280 ;
        RECT -3.240 92.020 -2.980 92.280 ;
        RECT 0.840 91.660 1.100 91.920 ;
        RECT 1.720 91.660 1.980 91.920 ;
        RECT 5.800 92.020 6.060 92.280 ;
        RECT 6.680 92.020 6.940 92.280 ;
        RECT 10.760 91.660 11.020 91.920 ;
        RECT 11.640 91.660 11.900 91.920 ;
        RECT 15.720 92.020 15.980 92.280 ;
        RECT 16.600 92.020 16.860 92.280 ;
        RECT 20.680 91.660 20.940 91.920 ;
        RECT 21.560 91.660 21.820 91.920 ;
        RECT 25.640 92.020 25.900 92.280 ;
        RECT -290.670 4.310 -290.410 4.570 ;
        RECT -286.590 3.950 -286.330 4.210 ;
        RECT -285.710 3.950 -285.450 4.210 ;
        RECT -281.630 4.310 -281.370 4.570 ;
        RECT -280.750 4.310 -280.490 4.570 ;
        RECT -276.670 3.950 -276.410 4.210 ;
        RECT -275.790 3.950 -275.530 4.210 ;
        RECT -271.710 4.310 -271.450 4.570 ;
        RECT -270.830 4.310 -270.570 4.570 ;
        RECT -266.750 3.950 -266.490 4.210 ;
        RECT -265.870 3.950 -265.610 4.210 ;
        RECT -261.790 4.310 -261.530 4.570 ;
        RECT -260.910 4.310 -260.650 4.570 ;
        RECT -256.830 3.950 -256.570 4.210 ;
        RECT -255.950 3.950 -255.690 4.210 ;
        RECT -251.870 4.310 -251.610 4.570 ;
        RECT -250.990 4.310 -250.730 4.570 ;
        RECT -246.910 3.950 -246.650 4.210 ;
        RECT -246.030 3.950 -245.770 4.210 ;
        RECT -241.950 4.310 -241.690 4.570 ;
        RECT -241.070 4.310 -240.810 4.570 ;
        RECT -236.990 3.950 -236.730 4.210 ;
        RECT -236.110 3.950 -235.850 4.210 ;
        RECT -232.030 4.310 -231.770 4.570 ;
        RECT -231.150 4.310 -230.890 4.570 ;
        RECT -227.070 3.950 -226.810 4.210 ;
        RECT -226.190 3.950 -225.930 4.210 ;
        RECT -222.110 4.310 -221.850 4.570 ;
        RECT -221.230 4.310 -220.970 4.570 ;
        RECT -217.150 3.950 -216.890 4.210 ;
        RECT -216.270 3.950 -216.010 4.210 ;
        RECT -212.190 4.310 -211.930 4.570 ;
        RECT -211.310 4.310 -211.050 4.570 ;
        RECT -207.230 3.950 -206.970 4.210 ;
        RECT -206.350 3.950 -206.090 4.210 ;
        RECT -202.270 4.310 -202.010 4.570 ;
        RECT -201.390 4.310 -201.130 4.570 ;
        RECT -197.310 3.950 -197.050 4.210 ;
        RECT -196.430 3.950 -196.170 4.210 ;
        RECT -192.350 4.310 -192.090 4.570 ;
        RECT -191.470 4.310 -191.210 4.570 ;
        RECT -187.390 3.950 -187.130 4.210 ;
        RECT -186.510 3.950 -186.250 4.210 ;
        RECT -182.430 4.310 -182.170 4.570 ;
        RECT -181.550 4.310 -181.290 4.570 ;
        RECT -177.470 3.950 -177.210 4.210 ;
        RECT -176.590 3.950 -176.330 4.210 ;
        RECT -172.510 4.310 -172.250 4.570 ;
        RECT -171.630 4.310 -171.370 4.570 ;
        RECT -167.550 3.950 -167.290 4.210 ;
        RECT -166.670 3.950 -166.410 4.210 ;
        RECT -162.590 4.310 -162.330 4.570 ;
        RECT -161.710 4.310 -161.450 4.570 ;
        RECT -157.630 3.950 -157.370 4.210 ;
        RECT -156.750 3.950 -156.490 4.210 ;
        RECT -152.670 4.310 -152.410 4.570 ;
        RECT -151.790 4.310 -151.530 4.570 ;
        RECT -147.710 3.950 -147.450 4.210 ;
        RECT -146.830 3.950 -146.570 4.210 ;
        RECT -142.750 4.310 -142.490 4.570 ;
        RECT -141.870 4.310 -141.610 4.570 ;
        RECT -137.790 3.950 -137.530 4.210 ;
        RECT -136.910 3.950 -136.650 4.210 ;
        RECT -132.830 4.310 -132.570 4.570 ;
        RECT -131.950 4.310 -131.690 4.570 ;
        RECT -127.870 3.950 -127.610 4.210 ;
        RECT -126.990 3.950 -126.730 4.210 ;
        RECT -122.910 4.310 -122.650 4.570 ;
        RECT -122.030 4.310 -121.770 4.570 ;
        RECT -117.950 3.950 -117.690 4.210 ;
        RECT -117.070 3.950 -116.810 4.210 ;
        RECT -112.990 4.310 -112.730 4.570 ;
        RECT -112.110 4.310 -111.850 4.570 ;
        RECT -108.030 3.950 -107.770 4.210 ;
        RECT -107.150 3.950 -106.890 4.210 ;
        RECT -103.070 4.310 -102.810 4.570 ;
        RECT -102.190 4.310 -101.930 4.570 ;
        RECT -98.110 3.950 -97.850 4.210 ;
        RECT -97.230 3.950 -96.970 4.210 ;
        RECT -93.150 4.310 -92.890 4.570 ;
        RECT -92.270 4.310 -92.010 4.570 ;
        RECT -88.190 3.950 -87.930 4.210 ;
        RECT -87.310 3.950 -87.050 4.210 ;
        RECT -83.230 4.310 -82.970 4.570 ;
        RECT -82.350 4.310 -82.090 4.570 ;
        RECT -78.270 3.950 -78.010 4.210 ;
        RECT -77.390 3.950 -77.130 4.210 ;
        RECT -73.310 4.310 -73.050 4.570 ;
        RECT -72.430 4.310 -72.170 4.570 ;
        RECT -68.350 3.950 -68.090 4.210 ;
        RECT -67.470 3.950 -67.210 4.210 ;
        RECT -63.390 4.310 -63.130 4.570 ;
        RECT -62.510 4.310 -62.250 4.570 ;
        RECT -58.430 3.950 -58.170 4.210 ;
        RECT -57.550 3.950 -57.290 4.210 ;
        RECT -53.470 4.310 -53.210 4.570 ;
        RECT -52.590 4.310 -52.330 4.570 ;
        RECT -48.510 3.950 -48.250 4.210 ;
        RECT -47.630 3.950 -47.370 4.210 ;
        RECT -43.550 4.310 -43.290 4.570 ;
        RECT -42.670 4.310 -42.410 4.570 ;
        RECT -38.590 3.950 -38.330 4.210 ;
        RECT -37.710 3.950 -37.450 4.210 ;
        RECT -33.630 4.310 -33.370 4.570 ;
        RECT -32.750 4.310 -32.490 4.570 ;
        RECT -28.670 3.950 -28.410 4.210 ;
        RECT -27.790 3.950 -27.530 4.210 ;
        RECT -23.710 4.310 -23.450 4.570 ;
        RECT -22.830 4.310 -22.570 4.570 ;
        RECT -18.750 3.950 -18.490 4.210 ;
        RECT -17.870 3.950 -17.610 4.210 ;
        RECT -13.790 4.310 -13.530 4.570 ;
        RECT -12.910 4.310 -12.650 4.570 ;
        RECT -8.830 3.950 -8.570 4.210 ;
        RECT -7.950 3.950 -7.690 4.210 ;
        RECT -3.870 4.310 -3.610 4.570 ;
        RECT -2.990 4.310 -2.730 4.570 ;
        RECT 1.090 3.950 1.350 4.210 ;
        RECT 1.970 3.950 2.230 4.210 ;
        RECT 6.050 4.310 6.310 4.570 ;
        RECT 6.930 4.310 7.190 4.570 ;
        RECT 11.010 3.950 11.270 4.210 ;
        RECT 11.890 3.950 12.150 4.210 ;
        RECT 15.970 4.310 16.230 4.570 ;
        RECT 16.850 4.310 17.110 4.570 ;
        RECT 20.930 3.950 21.190 4.210 ;
        RECT 21.810 3.950 22.070 4.210 ;
        RECT 25.890 4.310 26.150 4.570 ;
        RECT -288.910 -89.040 -288.650 -88.780 ;
        RECT -284.830 -89.400 -284.570 -89.140 ;
        RECT -283.950 -89.400 -283.690 -89.140 ;
        RECT -279.870 -89.040 -279.610 -88.780 ;
        RECT -278.990 -89.040 -278.730 -88.780 ;
        RECT -274.910 -89.400 -274.650 -89.140 ;
        RECT -274.030 -89.400 -273.770 -89.140 ;
        RECT -269.950 -89.040 -269.690 -88.780 ;
        RECT -269.070 -89.040 -268.810 -88.780 ;
        RECT -264.990 -89.400 -264.730 -89.140 ;
        RECT -264.110 -89.400 -263.850 -89.140 ;
        RECT -260.030 -89.040 -259.770 -88.780 ;
        RECT -259.150 -89.040 -258.890 -88.780 ;
        RECT -255.070 -89.400 -254.810 -89.140 ;
        RECT -254.190 -89.400 -253.930 -89.140 ;
        RECT -250.110 -89.040 -249.850 -88.780 ;
        RECT -249.230 -89.040 -248.970 -88.780 ;
        RECT -245.150 -89.400 -244.890 -89.140 ;
        RECT -244.270 -89.400 -244.010 -89.140 ;
        RECT -240.190 -89.040 -239.930 -88.780 ;
        RECT -239.310 -89.040 -239.050 -88.780 ;
        RECT -235.230 -89.400 -234.970 -89.140 ;
        RECT -234.350 -89.400 -234.090 -89.140 ;
        RECT -230.270 -89.040 -230.010 -88.780 ;
        RECT -229.390 -89.040 -229.130 -88.780 ;
        RECT -225.310 -89.400 -225.050 -89.140 ;
        RECT -224.430 -89.400 -224.170 -89.140 ;
        RECT -220.350 -89.040 -220.090 -88.780 ;
        RECT -219.470 -89.040 -219.210 -88.780 ;
        RECT -215.390 -89.400 -215.130 -89.140 ;
        RECT -214.510 -89.400 -214.250 -89.140 ;
        RECT -210.430 -89.040 -210.170 -88.780 ;
        RECT -209.550 -89.040 -209.290 -88.780 ;
        RECT -205.470 -89.400 -205.210 -89.140 ;
        RECT -204.590 -89.400 -204.330 -89.140 ;
        RECT -200.510 -89.040 -200.250 -88.780 ;
        RECT -199.630 -89.040 -199.370 -88.780 ;
        RECT -195.550 -89.400 -195.290 -89.140 ;
        RECT -194.670 -89.400 -194.410 -89.140 ;
        RECT -190.590 -89.040 -190.330 -88.780 ;
        RECT -189.710 -89.040 -189.450 -88.780 ;
        RECT -185.630 -89.400 -185.370 -89.140 ;
        RECT -184.750 -89.400 -184.490 -89.140 ;
        RECT -180.670 -89.040 -180.410 -88.780 ;
        RECT -179.790 -89.040 -179.530 -88.780 ;
        RECT -175.710 -89.400 -175.450 -89.140 ;
        RECT -174.830 -89.400 -174.570 -89.140 ;
        RECT -170.750 -89.040 -170.490 -88.780 ;
        RECT -169.870 -89.040 -169.610 -88.780 ;
        RECT -165.790 -89.400 -165.530 -89.140 ;
        RECT -164.910 -89.400 -164.650 -89.140 ;
        RECT -160.830 -89.040 -160.570 -88.780 ;
        RECT -159.950 -89.040 -159.690 -88.780 ;
        RECT -155.870 -89.400 -155.610 -89.140 ;
        RECT -154.990 -89.400 -154.730 -89.140 ;
        RECT -150.910 -89.040 -150.650 -88.780 ;
        RECT -150.030 -89.040 -149.770 -88.780 ;
        RECT -145.950 -89.400 -145.690 -89.140 ;
        RECT -145.070 -89.400 -144.810 -89.140 ;
        RECT -140.990 -89.040 -140.730 -88.780 ;
        RECT -140.110 -89.040 -139.850 -88.780 ;
        RECT -136.030 -89.400 -135.770 -89.140 ;
        RECT -135.150 -89.400 -134.890 -89.140 ;
        RECT -131.070 -89.040 -130.810 -88.780 ;
        RECT -130.190 -89.040 -129.930 -88.780 ;
        RECT -126.110 -89.400 -125.850 -89.140 ;
        RECT -125.230 -89.400 -124.970 -89.140 ;
        RECT -121.150 -89.040 -120.890 -88.780 ;
        RECT -120.270 -89.040 -120.010 -88.780 ;
        RECT -116.190 -89.400 -115.930 -89.140 ;
        RECT -115.310 -89.400 -115.050 -89.140 ;
        RECT -111.230 -89.040 -110.970 -88.780 ;
        RECT -110.350 -89.040 -110.090 -88.780 ;
        RECT -106.270 -89.400 -106.010 -89.140 ;
        RECT -105.390 -89.400 -105.130 -89.140 ;
        RECT -101.310 -89.040 -101.050 -88.780 ;
        RECT -100.430 -89.040 -100.170 -88.780 ;
        RECT -96.350 -89.400 -96.090 -89.140 ;
        RECT -95.470 -89.400 -95.210 -89.140 ;
        RECT -91.390 -89.040 -91.130 -88.780 ;
        RECT -90.510 -89.040 -90.250 -88.780 ;
        RECT -86.430 -89.400 -86.170 -89.140 ;
        RECT -85.550 -89.400 -85.290 -89.140 ;
        RECT -81.470 -89.040 -81.210 -88.780 ;
        RECT -80.590 -89.040 -80.330 -88.780 ;
        RECT -76.510 -89.400 -76.250 -89.140 ;
        RECT -75.630 -89.400 -75.370 -89.140 ;
        RECT -71.550 -89.040 -71.290 -88.780 ;
        RECT -70.670 -89.040 -70.410 -88.780 ;
        RECT -66.590 -89.400 -66.330 -89.140 ;
        RECT -65.710 -89.400 -65.450 -89.140 ;
        RECT -61.630 -89.040 -61.370 -88.780 ;
        RECT -60.750 -89.040 -60.490 -88.780 ;
        RECT -56.670 -89.400 -56.410 -89.140 ;
        RECT -55.790 -89.400 -55.530 -89.140 ;
        RECT -51.710 -89.040 -51.450 -88.780 ;
        RECT -50.830 -89.040 -50.570 -88.780 ;
        RECT -46.750 -89.400 -46.490 -89.140 ;
        RECT -45.870 -89.400 -45.610 -89.140 ;
        RECT -41.790 -89.040 -41.530 -88.780 ;
        RECT -40.910 -89.040 -40.650 -88.780 ;
        RECT -36.830 -89.400 -36.570 -89.140 ;
        RECT -35.950 -89.400 -35.690 -89.140 ;
        RECT -31.870 -89.040 -31.610 -88.780 ;
        RECT -30.990 -89.040 -30.730 -88.780 ;
        RECT -26.910 -89.400 -26.650 -89.140 ;
        RECT -26.030 -89.400 -25.770 -89.140 ;
        RECT -21.950 -89.040 -21.690 -88.780 ;
        RECT -21.070 -89.040 -20.810 -88.780 ;
        RECT -16.990 -89.400 -16.730 -89.140 ;
        RECT -16.110 -89.400 -15.850 -89.140 ;
        RECT -12.030 -89.040 -11.770 -88.780 ;
        RECT -11.150 -89.040 -10.890 -88.780 ;
        RECT -7.070 -89.400 -6.810 -89.140 ;
        RECT -6.190 -89.400 -5.930 -89.140 ;
        RECT -2.110 -89.040 -1.850 -88.780 ;
        RECT -1.230 -89.040 -0.970 -88.780 ;
        RECT 2.850 -89.400 3.110 -89.140 ;
        RECT 3.730 -89.400 3.990 -89.140 ;
        RECT 7.810 -89.040 8.070 -88.780 ;
        RECT 8.690 -89.040 8.950 -88.780 ;
        RECT 12.770 -89.400 13.030 -89.140 ;
        RECT 13.650 -89.400 13.910 -89.140 ;
        RECT 17.730 -89.040 17.990 -88.780 ;
        RECT 18.610 -89.040 18.870 -88.780 ;
        RECT 22.690 -89.400 22.950 -89.140 ;
        RECT 23.570 -89.400 23.830 -89.140 ;
        RECT 27.650 -89.040 27.910 -88.780 ;
        RECT -288.660 -176.750 -288.400 -176.490 ;
        RECT -284.580 -177.110 -284.320 -176.850 ;
        RECT -283.700 -177.110 -283.440 -176.850 ;
        RECT -279.620 -176.750 -279.360 -176.490 ;
        RECT -278.740 -176.750 -278.480 -176.490 ;
        RECT -274.660 -177.110 -274.400 -176.850 ;
        RECT -273.780 -177.110 -273.520 -176.850 ;
        RECT -269.700 -176.750 -269.440 -176.490 ;
        RECT -268.820 -176.750 -268.560 -176.490 ;
        RECT -264.740 -177.110 -264.480 -176.850 ;
        RECT -263.860 -177.110 -263.600 -176.850 ;
        RECT -259.780 -176.750 -259.520 -176.490 ;
        RECT -258.900 -176.750 -258.640 -176.490 ;
        RECT -254.820 -177.110 -254.560 -176.850 ;
        RECT -253.940 -177.110 -253.680 -176.850 ;
        RECT -249.860 -176.750 -249.600 -176.490 ;
        RECT -248.980 -176.750 -248.720 -176.490 ;
        RECT -244.900 -177.110 -244.640 -176.850 ;
        RECT -244.020 -177.110 -243.760 -176.850 ;
        RECT -239.940 -176.750 -239.680 -176.490 ;
        RECT -239.060 -176.750 -238.800 -176.490 ;
        RECT -234.980 -177.110 -234.720 -176.850 ;
        RECT -234.100 -177.110 -233.840 -176.850 ;
        RECT -230.020 -176.750 -229.760 -176.490 ;
        RECT -229.140 -176.750 -228.880 -176.490 ;
        RECT -225.060 -177.110 -224.800 -176.850 ;
        RECT -224.180 -177.110 -223.920 -176.850 ;
        RECT -220.100 -176.750 -219.840 -176.490 ;
        RECT -219.220 -176.750 -218.960 -176.490 ;
        RECT -215.140 -177.110 -214.880 -176.850 ;
        RECT -214.260 -177.110 -214.000 -176.850 ;
        RECT -210.180 -176.750 -209.920 -176.490 ;
        RECT -209.300 -176.750 -209.040 -176.490 ;
        RECT -205.220 -177.110 -204.960 -176.850 ;
        RECT -204.340 -177.110 -204.080 -176.850 ;
        RECT -200.260 -176.750 -200.000 -176.490 ;
        RECT -199.380 -176.750 -199.120 -176.490 ;
        RECT -195.300 -177.110 -195.040 -176.850 ;
        RECT -194.420 -177.110 -194.160 -176.850 ;
        RECT -190.340 -176.750 -190.080 -176.490 ;
        RECT -189.460 -176.750 -189.200 -176.490 ;
        RECT -185.380 -177.110 -185.120 -176.850 ;
        RECT -184.500 -177.110 -184.240 -176.850 ;
        RECT -180.420 -176.750 -180.160 -176.490 ;
        RECT -179.540 -176.750 -179.280 -176.490 ;
        RECT -175.460 -177.110 -175.200 -176.850 ;
        RECT -174.580 -177.110 -174.320 -176.850 ;
        RECT -170.500 -176.750 -170.240 -176.490 ;
        RECT -169.620 -176.750 -169.360 -176.490 ;
        RECT -165.540 -177.110 -165.280 -176.850 ;
        RECT -164.660 -177.110 -164.400 -176.850 ;
        RECT -160.580 -176.750 -160.320 -176.490 ;
        RECT -159.700 -176.750 -159.440 -176.490 ;
        RECT -155.620 -177.110 -155.360 -176.850 ;
        RECT -154.740 -177.110 -154.480 -176.850 ;
        RECT -150.660 -176.750 -150.400 -176.490 ;
        RECT -149.780 -176.750 -149.520 -176.490 ;
        RECT -145.700 -177.110 -145.440 -176.850 ;
        RECT -144.820 -177.110 -144.560 -176.850 ;
        RECT -140.740 -176.750 -140.480 -176.490 ;
        RECT -139.860 -176.750 -139.600 -176.490 ;
        RECT -135.780 -177.110 -135.520 -176.850 ;
        RECT -134.900 -177.110 -134.640 -176.850 ;
        RECT -130.820 -176.750 -130.560 -176.490 ;
        RECT -129.940 -176.750 -129.680 -176.490 ;
        RECT -125.860 -177.110 -125.600 -176.850 ;
        RECT -124.980 -177.110 -124.720 -176.850 ;
        RECT -120.900 -176.750 -120.640 -176.490 ;
        RECT -120.020 -176.750 -119.760 -176.490 ;
        RECT -115.940 -177.110 -115.680 -176.850 ;
        RECT -115.060 -177.110 -114.800 -176.850 ;
        RECT -110.980 -176.750 -110.720 -176.490 ;
        RECT -110.100 -176.750 -109.840 -176.490 ;
        RECT -106.020 -177.110 -105.760 -176.850 ;
        RECT -105.140 -177.110 -104.880 -176.850 ;
        RECT -101.060 -176.750 -100.800 -176.490 ;
        RECT -100.180 -176.750 -99.920 -176.490 ;
        RECT -96.100 -177.110 -95.840 -176.850 ;
        RECT -95.220 -177.110 -94.960 -176.850 ;
        RECT -91.140 -176.750 -90.880 -176.490 ;
        RECT -90.260 -176.750 -90.000 -176.490 ;
        RECT -86.180 -177.110 -85.920 -176.850 ;
        RECT -85.300 -177.110 -85.040 -176.850 ;
        RECT -81.220 -176.750 -80.960 -176.490 ;
        RECT -80.340 -176.750 -80.080 -176.490 ;
        RECT -76.260 -177.110 -76.000 -176.850 ;
        RECT -75.380 -177.110 -75.120 -176.850 ;
        RECT -71.300 -176.750 -71.040 -176.490 ;
        RECT -70.420 -176.750 -70.160 -176.490 ;
        RECT -66.340 -177.110 -66.080 -176.850 ;
        RECT -65.460 -177.110 -65.200 -176.850 ;
        RECT -61.380 -176.750 -61.120 -176.490 ;
        RECT -60.500 -176.750 -60.240 -176.490 ;
        RECT -56.420 -177.110 -56.160 -176.850 ;
        RECT -55.540 -177.110 -55.280 -176.850 ;
        RECT -51.460 -176.750 -51.200 -176.490 ;
        RECT -50.580 -176.750 -50.320 -176.490 ;
        RECT -46.500 -177.110 -46.240 -176.850 ;
        RECT -45.620 -177.110 -45.360 -176.850 ;
        RECT -41.540 -176.750 -41.280 -176.490 ;
        RECT -40.660 -176.750 -40.400 -176.490 ;
        RECT -36.580 -177.110 -36.320 -176.850 ;
        RECT -35.700 -177.110 -35.440 -176.850 ;
        RECT -31.620 -176.750 -31.360 -176.490 ;
        RECT -30.740 -176.750 -30.480 -176.490 ;
        RECT -26.660 -177.110 -26.400 -176.850 ;
        RECT -25.780 -177.110 -25.520 -176.850 ;
        RECT -21.700 -176.750 -21.440 -176.490 ;
        RECT -20.820 -176.750 -20.560 -176.490 ;
        RECT -16.740 -177.110 -16.480 -176.850 ;
        RECT -15.860 -177.110 -15.600 -176.850 ;
        RECT -11.780 -176.750 -11.520 -176.490 ;
        RECT -10.900 -176.750 -10.640 -176.490 ;
        RECT -6.820 -177.110 -6.560 -176.850 ;
        RECT -5.940 -177.110 -5.680 -176.850 ;
        RECT -1.860 -176.750 -1.600 -176.490 ;
        RECT -0.980 -176.750 -0.720 -176.490 ;
        RECT 3.100 -177.110 3.360 -176.850 ;
        RECT 3.980 -177.110 4.240 -176.850 ;
        RECT 8.060 -176.750 8.320 -176.490 ;
        RECT 8.940 -176.750 9.200 -176.490 ;
        RECT 13.020 -177.110 13.280 -176.850 ;
        RECT 13.900 -177.110 14.160 -176.850 ;
        RECT 17.980 -176.750 18.240 -176.490 ;
        RECT 18.860 -176.750 19.120 -176.490 ;
        RECT 22.940 -177.110 23.200 -176.850 ;
        RECT 23.820 -177.110 24.080 -176.850 ;
        RECT 27.900 -176.750 28.160 -176.490 ;
      LAYER met2 ;
        RECT 37.260 96.660 37.720 96.680 ;
        RECT 39.160 96.660 39.950 96.740 ;
        RECT 37.260 95.310 39.950 96.660 ;
        RECT -291.010 92.040 -290.550 92.350 ;
        RECT -288.820 92.040 -288.680 92.440 ;
        RECT -283.860 92.040 -283.720 92.440 ;
        RECT -281.990 92.040 -280.630 92.350 ;
        RECT -278.900 92.040 -278.760 92.440 ;
        RECT -273.940 92.040 -273.800 92.440 ;
        RECT -272.070 92.040 -270.710 92.350 ;
        RECT -268.980 92.040 -268.840 92.440 ;
        RECT -264.020 92.040 -263.880 92.440 ;
        RECT -262.150 92.040 -260.790 92.350 ;
        RECT -259.060 92.040 -258.920 92.440 ;
        RECT -254.100 92.040 -253.960 92.440 ;
        RECT -252.230 92.040 -250.870 92.350 ;
        RECT -249.140 92.040 -249.000 92.440 ;
        RECT -244.180 92.040 -244.040 92.440 ;
        RECT -242.310 92.040 -240.950 92.350 ;
        RECT -239.220 92.040 -239.080 92.440 ;
        RECT -234.260 92.040 -234.120 92.440 ;
        RECT -232.390 92.040 -231.030 92.350 ;
        RECT -229.300 92.040 -229.160 92.440 ;
        RECT -224.340 92.040 -224.200 92.440 ;
        RECT -222.470 92.040 -221.110 92.350 ;
        RECT -219.380 92.040 -219.240 92.440 ;
        RECT -214.420 92.040 -214.280 92.440 ;
        RECT -212.550 92.040 -211.190 92.350 ;
        RECT -209.460 92.040 -209.320 92.440 ;
        RECT -204.500 92.040 -204.360 92.440 ;
        RECT -202.630 92.040 -201.270 92.350 ;
        RECT -199.540 92.040 -199.400 92.440 ;
        RECT -194.580 92.040 -194.440 92.440 ;
        RECT -192.710 92.040 -191.350 92.350 ;
        RECT -189.620 92.040 -189.480 92.440 ;
        RECT -184.660 92.040 -184.520 92.440 ;
        RECT -182.790 92.040 -181.430 92.350 ;
        RECT -179.700 92.040 -179.560 92.440 ;
        RECT -174.740 92.040 -174.600 92.440 ;
        RECT -172.870 92.040 -171.510 92.350 ;
        RECT -169.780 92.040 -169.640 92.440 ;
        RECT -164.820 92.040 -164.680 92.440 ;
        RECT -162.950 92.040 -161.590 92.350 ;
        RECT -159.860 92.040 -159.720 92.440 ;
        RECT -154.900 92.040 -154.760 92.440 ;
        RECT -153.030 92.040 -151.670 92.350 ;
        RECT -149.940 92.040 -149.800 92.440 ;
        RECT -144.980 92.040 -144.840 92.440 ;
        RECT -143.110 92.040 -141.750 92.350 ;
        RECT -140.020 92.040 -139.880 92.440 ;
        RECT -135.060 92.040 -134.920 92.440 ;
        RECT -133.190 92.040 -131.830 92.350 ;
        RECT -130.100 92.040 -129.960 92.440 ;
        RECT -125.140 92.040 -125.000 92.440 ;
        RECT -123.270 92.040 -121.910 92.350 ;
        RECT -120.180 92.040 -120.040 92.440 ;
        RECT -115.220 92.040 -115.080 92.440 ;
        RECT -113.350 92.040 -111.990 92.350 ;
        RECT -110.260 92.040 -110.120 92.440 ;
        RECT -105.300 92.040 -105.160 92.440 ;
        RECT -103.430 92.040 -102.070 92.350 ;
        RECT -100.340 92.040 -100.200 92.440 ;
        RECT -95.380 92.040 -95.240 92.440 ;
        RECT -93.510 92.040 -92.150 92.350 ;
        RECT -90.420 92.040 -90.280 92.440 ;
        RECT -85.460 92.040 -85.320 92.440 ;
        RECT -83.590 92.040 -82.230 92.350 ;
        RECT -80.500 92.040 -80.360 92.440 ;
        RECT -75.540 92.040 -75.400 92.440 ;
        RECT -73.670 92.040 -72.310 92.350 ;
        RECT -70.580 92.040 -70.440 92.440 ;
        RECT -65.620 92.040 -65.480 92.440 ;
        RECT -63.750 92.040 -62.390 92.350 ;
        RECT -60.660 92.040 -60.520 92.440 ;
        RECT -55.700 92.040 -55.560 92.440 ;
        RECT -53.830 92.040 -52.470 92.350 ;
        RECT -50.740 92.040 -50.600 92.440 ;
        RECT -45.780 92.040 -45.640 92.440 ;
        RECT -43.910 92.040 -42.550 92.350 ;
        RECT -40.820 92.040 -40.680 92.440 ;
        RECT -35.860 92.040 -35.720 92.440 ;
        RECT -33.990 92.040 -32.630 92.350 ;
        RECT -30.900 92.040 -30.760 92.440 ;
        RECT -25.940 92.040 -25.800 92.440 ;
        RECT -24.070 92.040 -22.710 92.350 ;
        RECT -20.980 92.040 -20.840 92.440 ;
        RECT -16.020 92.040 -15.880 92.440 ;
        RECT -14.150 92.040 -12.790 92.350 ;
        RECT -11.060 92.040 -10.920 92.440 ;
        RECT -6.100 92.040 -5.960 92.440 ;
        RECT -4.230 92.040 -2.870 92.350 ;
        RECT -1.140 92.040 -1.000 92.440 ;
        RECT 3.820 92.040 3.960 92.440 ;
        RECT 5.690 92.040 7.050 92.350 ;
        RECT 8.780 92.040 8.920 92.440 ;
        RECT 13.740 92.040 13.880 92.440 ;
        RECT 15.610 92.040 16.970 92.350 ;
        RECT 18.700 92.040 18.840 92.440 ;
        RECT 23.660 92.040 23.800 92.440 ;
        RECT 37.260 92.370 37.720 95.310 ;
        RECT 32.950 92.360 37.720 92.370 ;
        RECT 25.530 92.040 37.720 92.360 ;
        RECT -291.010 91.910 37.720 92.040 ;
        RECT -291.010 91.900 34.270 91.910 ;
        RECT -288.820 91.500 -288.680 91.900 ;
        RECT -286.950 91.590 -285.590 91.900 ;
        RECT -283.860 91.500 -283.720 91.900 ;
        RECT -278.900 91.500 -278.760 91.900 ;
        RECT -277.030 91.590 -275.670 91.900 ;
        RECT -273.940 91.500 -273.800 91.900 ;
        RECT -268.980 91.500 -268.840 91.900 ;
        RECT -267.110 91.590 -265.750 91.900 ;
        RECT -264.020 91.500 -263.880 91.900 ;
        RECT -259.060 91.500 -258.920 91.900 ;
        RECT -257.190 91.590 -255.830 91.900 ;
        RECT -254.100 91.500 -253.960 91.900 ;
        RECT -249.140 91.500 -249.000 91.900 ;
        RECT -247.270 91.590 -245.910 91.900 ;
        RECT -244.180 91.500 -244.040 91.900 ;
        RECT -239.220 91.500 -239.080 91.900 ;
        RECT -237.350 91.590 -235.990 91.900 ;
        RECT -234.260 91.500 -234.120 91.900 ;
        RECT -229.300 91.500 -229.160 91.900 ;
        RECT -227.430 91.590 -226.070 91.900 ;
        RECT -224.340 91.500 -224.200 91.900 ;
        RECT -219.380 91.500 -219.240 91.900 ;
        RECT -217.510 91.590 -216.150 91.900 ;
        RECT -214.420 91.500 -214.280 91.900 ;
        RECT -209.460 91.500 -209.320 91.900 ;
        RECT -207.590 91.590 -206.230 91.900 ;
        RECT -204.500 91.500 -204.360 91.900 ;
        RECT -199.540 91.500 -199.400 91.900 ;
        RECT -197.670 91.590 -196.310 91.900 ;
        RECT -194.580 91.500 -194.440 91.900 ;
        RECT -189.620 91.500 -189.480 91.900 ;
        RECT -187.750 91.590 -186.390 91.900 ;
        RECT -184.660 91.500 -184.520 91.900 ;
        RECT -179.700 91.500 -179.560 91.900 ;
        RECT -177.830 91.590 -176.470 91.900 ;
        RECT -174.740 91.500 -174.600 91.900 ;
        RECT -169.780 91.500 -169.640 91.900 ;
        RECT -167.910 91.590 -166.550 91.900 ;
        RECT -164.820 91.500 -164.680 91.900 ;
        RECT -159.860 91.500 -159.720 91.900 ;
        RECT -157.990 91.590 -156.630 91.900 ;
        RECT -154.900 91.500 -154.760 91.900 ;
        RECT -149.940 91.500 -149.800 91.900 ;
        RECT -148.070 91.590 -146.710 91.900 ;
        RECT -144.980 91.500 -144.840 91.900 ;
        RECT -140.020 91.500 -139.880 91.900 ;
        RECT -138.150 91.590 -136.790 91.900 ;
        RECT -135.060 91.500 -134.920 91.900 ;
        RECT -130.100 91.500 -129.960 91.900 ;
        RECT -128.230 91.590 -126.870 91.900 ;
        RECT -125.140 91.500 -125.000 91.900 ;
        RECT -120.180 91.500 -120.040 91.900 ;
        RECT -118.310 91.590 -116.950 91.900 ;
        RECT -115.220 91.500 -115.080 91.900 ;
        RECT -110.260 91.500 -110.120 91.900 ;
        RECT -108.390 91.590 -107.030 91.900 ;
        RECT -105.300 91.500 -105.160 91.900 ;
        RECT -100.340 91.500 -100.200 91.900 ;
        RECT -98.470 91.590 -97.110 91.900 ;
        RECT -95.380 91.500 -95.240 91.900 ;
        RECT -90.420 91.500 -90.280 91.900 ;
        RECT -88.550 91.590 -87.190 91.900 ;
        RECT -85.460 91.500 -85.320 91.900 ;
        RECT -80.500 91.500 -80.360 91.900 ;
        RECT -78.630 91.590 -77.270 91.900 ;
        RECT -75.540 91.500 -75.400 91.900 ;
        RECT -70.580 91.500 -70.440 91.900 ;
        RECT -68.710 91.590 -67.350 91.900 ;
        RECT -65.620 91.500 -65.480 91.900 ;
        RECT -60.660 91.500 -60.520 91.900 ;
        RECT -58.790 91.590 -57.430 91.900 ;
        RECT -55.700 91.500 -55.560 91.900 ;
        RECT -50.740 91.500 -50.600 91.900 ;
        RECT -48.870 91.590 -47.510 91.900 ;
        RECT -45.780 91.500 -45.640 91.900 ;
        RECT -40.820 91.500 -40.680 91.900 ;
        RECT -38.950 91.590 -37.590 91.900 ;
        RECT -35.860 91.500 -35.720 91.900 ;
        RECT -30.900 91.500 -30.760 91.900 ;
        RECT -29.030 91.590 -27.670 91.900 ;
        RECT -25.940 91.500 -25.800 91.900 ;
        RECT -20.980 91.500 -20.840 91.900 ;
        RECT -19.110 91.590 -17.750 91.900 ;
        RECT -16.020 91.500 -15.880 91.900 ;
        RECT -11.060 91.500 -10.920 91.900 ;
        RECT -9.190 91.590 -7.830 91.900 ;
        RECT -6.100 91.500 -5.960 91.900 ;
        RECT -1.140 91.500 -1.000 91.900 ;
        RECT 0.730 91.590 2.090 91.900 ;
        RECT 3.820 91.500 3.960 91.900 ;
        RECT 8.780 91.500 8.920 91.900 ;
        RECT 10.650 91.590 12.010 91.900 ;
        RECT 13.740 91.500 13.880 91.900 ;
        RECT 18.700 91.500 18.840 91.900 ;
        RECT 20.570 91.590 21.930 91.900 ;
        RECT 23.660 91.500 23.800 91.900 ;
        RECT 39.160 83.840 39.950 95.310 ;
        RECT 39.160 9.780 39.860 83.840 ;
        RECT 37.600 8.970 39.860 9.780 ;
        RECT 37.510 8.080 39.860 8.970 ;
        RECT -290.760 4.330 -290.300 4.640 ;
        RECT -288.570 4.330 -288.430 4.730 ;
        RECT -283.610 4.330 -283.470 4.730 ;
        RECT -281.740 4.330 -280.380 4.640 ;
        RECT -278.650 4.330 -278.510 4.730 ;
        RECT -273.690 4.330 -273.550 4.730 ;
        RECT -271.820 4.330 -270.460 4.640 ;
        RECT -268.730 4.330 -268.590 4.730 ;
        RECT -263.770 4.330 -263.630 4.730 ;
        RECT -261.900 4.330 -260.540 4.640 ;
        RECT -258.810 4.330 -258.670 4.730 ;
        RECT -253.850 4.330 -253.710 4.730 ;
        RECT -251.980 4.330 -250.620 4.640 ;
        RECT -248.890 4.330 -248.750 4.730 ;
        RECT -243.930 4.330 -243.790 4.730 ;
        RECT -242.060 4.330 -240.700 4.640 ;
        RECT -238.970 4.330 -238.830 4.730 ;
        RECT -234.010 4.330 -233.870 4.730 ;
        RECT -232.140 4.330 -230.780 4.640 ;
        RECT -229.050 4.330 -228.910 4.730 ;
        RECT -224.090 4.330 -223.950 4.730 ;
        RECT -222.220 4.330 -220.860 4.640 ;
        RECT -219.130 4.330 -218.990 4.730 ;
        RECT -214.170 4.330 -214.030 4.730 ;
        RECT -212.300 4.330 -210.940 4.640 ;
        RECT -209.210 4.330 -209.070 4.730 ;
        RECT -204.250 4.330 -204.110 4.730 ;
        RECT -202.380 4.330 -201.020 4.640 ;
        RECT -199.290 4.330 -199.150 4.730 ;
        RECT -194.330 4.330 -194.190 4.730 ;
        RECT -192.460 4.330 -191.100 4.640 ;
        RECT -189.370 4.330 -189.230 4.730 ;
        RECT -184.410 4.330 -184.270 4.730 ;
        RECT -182.540 4.330 -181.180 4.640 ;
        RECT -179.450 4.330 -179.310 4.730 ;
        RECT -174.490 4.330 -174.350 4.730 ;
        RECT -172.620 4.330 -171.260 4.640 ;
        RECT -169.530 4.330 -169.390 4.730 ;
        RECT -164.570 4.330 -164.430 4.730 ;
        RECT -162.700 4.330 -161.340 4.640 ;
        RECT -159.610 4.330 -159.470 4.730 ;
        RECT -154.650 4.330 -154.510 4.730 ;
        RECT -152.780 4.330 -151.420 4.640 ;
        RECT -149.690 4.330 -149.550 4.730 ;
        RECT -144.730 4.330 -144.590 4.730 ;
        RECT -142.860 4.330 -141.500 4.640 ;
        RECT -139.770 4.330 -139.630 4.730 ;
        RECT -134.810 4.330 -134.670 4.730 ;
        RECT -132.940 4.330 -131.580 4.640 ;
        RECT -129.850 4.330 -129.710 4.730 ;
        RECT -124.890 4.330 -124.750 4.730 ;
        RECT -123.020 4.330 -121.660 4.640 ;
        RECT -119.930 4.330 -119.790 4.730 ;
        RECT -114.970 4.330 -114.830 4.730 ;
        RECT -113.100 4.330 -111.740 4.640 ;
        RECT -110.010 4.330 -109.870 4.730 ;
        RECT -105.050 4.330 -104.910 4.730 ;
        RECT -103.180 4.330 -101.820 4.640 ;
        RECT -100.090 4.330 -99.950 4.730 ;
        RECT -95.130 4.330 -94.990 4.730 ;
        RECT -93.260 4.330 -91.900 4.640 ;
        RECT -90.170 4.330 -90.030 4.730 ;
        RECT -85.210 4.330 -85.070 4.730 ;
        RECT -83.340 4.330 -81.980 4.640 ;
        RECT -80.250 4.330 -80.110 4.730 ;
        RECT -75.290 4.330 -75.150 4.730 ;
        RECT -73.420 4.330 -72.060 4.640 ;
        RECT -70.330 4.330 -70.190 4.730 ;
        RECT -65.370 4.330 -65.230 4.730 ;
        RECT -63.500 4.330 -62.140 4.640 ;
        RECT -60.410 4.330 -60.270 4.730 ;
        RECT -55.450 4.330 -55.310 4.730 ;
        RECT -53.580 4.330 -52.220 4.640 ;
        RECT -50.490 4.330 -50.350 4.730 ;
        RECT -45.530 4.330 -45.390 4.730 ;
        RECT -43.660 4.330 -42.300 4.640 ;
        RECT -40.570 4.330 -40.430 4.730 ;
        RECT -35.610 4.330 -35.470 4.730 ;
        RECT -33.740 4.330 -32.380 4.640 ;
        RECT -30.650 4.330 -30.510 4.730 ;
        RECT -25.690 4.330 -25.550 4.730 ;
        RECT -23.820 4.330 -22.460 4.640 ;
        RECT -20.730 4.330 -20.590 4.730 ;
        RECT -15.770 4.330 -15.630 4.730 ;
        RECT -13.900 4.330 -12.540 4.640 ;
        RECT -10.810 4.330 -10.670 4.730 ;
        RECT -5.850 4.330 -5.710 4.730 ;
        RECT -3.980 4.330 -2.620 4.640 ;
        RECT -0.890 4.330 -0.750 4.730 ;
        RECT 4.070 4.330 4.210 4.730 ;
        RECT 5.940 4.330 7.300 4.640 ;
        RECT 9.030 4.330 9.170 4.730 ;
        RECT 13.990 4.330 14.130 4.730 ;
        RECT 15.860 4.330 17.220 4.640 ;
        RECT 18.950 4.330 19.090 4.730 ;
        RECT 23.910 4.330 24.050 4.730 ;
        RECT 37.510 4.660 37.970 8.080 ;
        RECT 33.200 4.650 37.970 4.660 ;
        RECT 25.780 4.330 37.970 4.650 ;
        RECT -290.760 4.200 37.970 4.330 ;
        RECT -290.760 4.190 34.520 4.200 ;
        RECT -288.570 3.790 -288.430 4.190 ;
        RECT -286.700 3.880 -285.340 4.190 ;
        RECT -283.610 3.790 -283.470 4.190 ;
        RECT -278.650 3.790 -278.510 4.190 ;
        RECT -276.780 3.880 -275.420 4.190 ;
        RECT -273.690 3.790 -273.550 4.190 ;
        RECT -268.730 3.790 -268.590 4.190 ;
        RECT -266.860 3.880 -265.500 4.190 ;
        RECT -263.770 3.790 -263.630 4.190 ;
        RECT -258.810 3.790 -258.670 4.190 ;
        RECT -256.940 3.880 -255.580 4.190 ;
        RECT -253.850 3.790 -253.710 4.190 ;
        RECT -248.890 3.790 -248.750 4.190 ;
        RECT -247.020 3.880 -245.660 4.190 ;
        RECT -243.930 3.790 -243.790 4.190 ;
        RECT -238.970 3.790 -238.830 4.190 ;
        RECT -237.100 3.880 -235.740 4.190 ;
        RECT -234.010 3.790 -233.870 4.190 ;
        RECT -229.050 3.790 -228.910 4.190 ;
        RECT -227.180 3.880 -225.820 4.190 ;
        RECT -224.090 3.790 -223.950 4.190 ;
        RECT -219.130 3.790 -218.990 4.190 ;
        RECT -217.260 3.880 -215.900 4.190 ;
        RECT -214.170 3.790 -214.030 4.190 ;
        RECT -209.210 3.790 -209.070 4.190 ;
        RECT -207.340 3.880 -205.980 4.190 ;
        RECT -204.250 3.790 -204.110 4.190 ;
        RECT -199.290 3.790 -199.150 4.190 ;
        RECT -197.420 3.880 -196.060 4.190 ;
        RECT -194.330 3.790 -194.190 4.190 ;
        RECT -189.370 3.790 -189.230 4.190 ;
        RECT -187.500 3.880 -186.140 4.190 ;
        RECT -184.410 3.790 -184.270 4.190 ;
        RECT -179.450 3.790 -179.310 4.190 ;
        RECT -177.580 3.880 -176.220 4.190 ;
        RECT -174.490 3.790 -174.350 4.190 ;
        RECT -169.530 3.790 -169.390 4.190 ;
        RECT -167.660 3.880 -166.300 4.190 ;
        RECT -164.570 3.790 -164.430 4.190 ;
        RECT -159.610 3.790 -159.470 4.190 ;
        RECT -157.740 3.880 -156.380 4.190 ;
        RECT -154.650 3.790 -154.510 4.190 ;
        RECT -149.690 3.790 -149.550 4.190 ;
        RECT -147.820 3.880 -146.460 4.190 ;
        RECT -144.730 3.790 -144.590 4.190 ;
        RECT -139.770 3.790 -139.630 4.190 ;
        RECT -137.900 3.880 -136.540 4.190 ;
        RECT -134.810 3.790 -134.670 4.190 ;
        RECT -129.850 3.790 -129.710 4.190 ;
        RECT -127.980 3.880 -126.620 4.190 ;
        RECT -124.890 3.790 -124.750 4.190 ;
        RECT -119.930 3.790 -119.790 4.190 ;
        RECT -118.060 3.880 -116.700 4.190 ;
        RECT -114.970 3.790 -114.830 4.190 ;
        RECT -110.010 3.790 -109.870 4.190 ;
        RECT -108.140 3.880 -106.780 4.190 ;
        RECT -105.050 3.790 -104.910 4.190 ;
        RECT -100.090 3.790 -99.950 4.190 ;
        RECT -98.220 3.880 -96.860 4.190 ;
        RECT -95.130 3.790 -94.990 4.190 ;
        RECT -90.170 3.790 -90.030 4.190 ;
        RECT -88.300 3.880 -86.940 4.190 ;
        RECT -85.210 3.790 -85.070 4.190 ;
        RECT -80.250 3.790 -80.110 4.190 ;
        RECT -78.380 3.880 -77.020 4.190 ;
        RECT -75.290 3.790 -75.150 4.190 ;
        RECT -70.330 3.790 -70.190 4.190 ;
        RECT -68.460 3.880 -67.100 4.190 ;
        RECT -65.370 3.790 -65.230 4.190 ;
        RECT -60.410 3.790 -60.270 4.190 ;
        RECT -58.540 3.880 -57.180 4.190 ;
        RECT -55.450 3.790 -55.310 4.190 ;
        RECT -50.490 3.790 -50.350 4.190 ;
        RECT -48.620 3.880 -47.260 4.190 ;
        RECT -45.530 3.790 -45.390 4.190 ;
        RECT -40.570 3.790 -40.430 4.190 ;
        RECT -38.700 3.880 -37.340 4.190 ;
        RECT -35.610 3.790 -35.470 4.190 ;
        RECT -30.650 3.790 -30.510 4.190 ;
        RECT -28.780 3.880 -27.420 4.190 ;
        RECT -25.690 3.790 -25.550 4.190 ;
        RECT -20.730 3.790 -20.590 4.190 ;
        RECT -18.860 3.880 -17.500 4.190 ;
        RECT -15.770 3.790 -15.630 4.190 ;
        RECT -10.810 3.790 -10.670 4.190 ;
        RECT -8.940 3.880 -7.580 4.190 ;
        RECT -5.850 3.790 -5.710 4.190 ;
        RECT -0.890 3.790 -0.750 4.190 ;
        RECT 0.980 3.880 2.340 4.190 ;
        RECT 4.070 3.790 4.210 4.190 ;
        RECT 9.030 3.790 9.170 4.190 ;
        RECT 10.900 3.880 12.260 4.190 ;
        RECT 13.990 3.790 14.130 4.190 ;
        RECT 18.950 3.790 19.090 4.190 ;
        RECT 20.820 3.880 22.180 4.190 ;
        RECT 23.910 3.790 24.050 4.190 ;
        RECT 39.160 2.190 39.860 8.080 ;
        RECT 39.160 -3.260 39.960 2.190 ;
        RECT 39.260 -84.280 39.960 -3.260 ;
        RECT 39.260 -87.390 40.110 -84.280 ;
        RECT -289.000 -89.020 -288.540 -88.710 ;
        RECT -286.810 -89.020 -286.670 -88.620 ;
        RECT -281.850 -89.020 -281.710 -88.620 ;
        RECT -279.980 -89.020 -278.620 -88.710 ;
        RECT -276.890 -89.020 -276.750 -88.620 ;
        RECT -271.930 -89.020 -271.790 -88.620 ;
        RECT -270.060 -89.020 -268.700 -88.710 ;
        RECT -266.970 -89.020 -266.830 -88.620 ;
        RECT -262.010 -89.020 -261.870 -88.620 ;
        RECT -260.140 -89.020 -258.780 -88.710 ;
        RECT -257.050 -89.020 -256.910 -88.620 ;
        RECT -252.090 -89.020 -251.950 -88.620 ;
        RECT -250.220 -89.020 -248.860 -88.710 ;
        RECT -247.130 -89.020 -246.990 -88.620 ;
        RECT -242.170 -89.020 -242.030 -88.620 ;
        RECT -240.300 -89.020 -238.940 -88.710 ;
        RECT -237.210 -89.020 -237.070 -88.620 ;
        RECT -232.250 -89.020 -232.110 -88.620 ;
        RECT -230.380 -89.020 -229.020 -88.710 ;
        RECT -227.290 -89.020 -227.150 -88.620 ;
        RECT -222.330 -89.020 -222.190 -88.620 ;
        RECT -220.460 -89.020 -219.100 -88.710 ;
        RECT -217.370 -89.020 -217.230 -88.620 ;
        RECT -212.410 -89.020 -212.270 -88.620 ;
        RECT -210.540 -89.020 -209.180 -88.710 ;
        RECT -207.450 -89.020 -207.310 -88.620 ;
        RECT -202.490 -89.020 -202.350 -88.620 ;
        RECT -200.620 -89.020 -199.260 -88.710 ;
        RECT -197.530 -89.020 -197.390 -88.620 ;
        RECT -192.570 -89.020 -192.430 -88.620 ;
        RECT -190.700 -89.020 -189.340 -88.710 ;
        RECT -187.610 -89.020 -187.470 -88.620 ;
        RECT -182.650 -89.020 -182.510 -88.620 ;
        RECT -180.780 -89.020 -179.420 -88.710 ;
        RECT -177.690 -89.020 -177.550 -88.620 ;
        RECT -172.730 -89.020 -172.590 -88.620 ;
        RECT -170.860 -89.020 -169.500 -88.710 ;
        RECT -167.770 -89.020 -167.630 -88.620 ;
        RECT -162.810 -89.020 -162.670 -88.620 ;
        RECT -160.940 -89.020 -159.580 -88.710 ;
        RECT -157.850 -89.020 -157.710 -88.620 ;
        RECT -152.890 -89.020 -152.750 -88.620 ;
        RECT -151.020 -89.020 -149.660 -88.710 ;
        RECT -147.930 -89.020 -147.790 -88.620 ;
        RECT -142.970 -89.020 -142.830 -88.620 ;
        RECT -141.100 -89.020 -139.740 -88.710 ;
        RECT -138.010 -89.020 -137.870 -88.620 ;
        RECT -133.050 -89.020 -132.910 -88.620 ;
        RECT -131.180 -89.020 -129.820 -88.710 ;
        RECT -128.090 -89.020 -127.950 -88.620 ;
        RECT -123.130 -89.020 -122.990 -88.620 ;
        RECT -121.260 -89.020 -119.900 -88.710 ;
        RECT -118.170 -89.020 -118.030 -88.620 ;
        RECT -113.210 -89.020 -113.070 -88.620 ;
        RECT -111.340 -89.020 -109.980 -88.710 ;
        RECT -108.250 -89.020 -108.110 -88.620 ;
        RECT -103.290 -89.020 -103.150 -88.620 ;
        RECT -101.420 -89.020 -100.060 -88.710 ;
        RECT -98.330 -89.020 -98.190 -88.620 ;
        RECT -93.370 -89.020 -93.230 -88.620 ;
        RECT -91.500 -89.020 -90.140 -88.710 ;
        RECT -88.410 -89.020 -88.270 -88.620 ;
        RECT -83.450 -89.020 -83.310 -88.620 ;
        RECT -81.580 -89.020 -80.220 -88.710 ;
        RECT -78.490 -89.020 -78.350 -88.620 ;
        RECT -73.530 -89.020 -73.390 -88.620 ;
        RECT -71.660 -89.020 -70.300 -88.710 ;
        RECT -68.570 -89.020 -68.430 -88.620 ;
        RECT -63.610 -89.020 -63.470 -88.620 ;
        RECT -61.740 -89.020 -60.380 -88.710 ;
        RECT -58.650 -89.020 -58.510 -88.620 ;
        RECT -53.690 -89.020 -53.550 -88.620 ;
        RECT -51.820 -89.020 -50.460 -88.710 ;
        RECT -48.730 -89.020 -48.590 -88.620 ;
        RECT -43.770 -89.020 -43.630 -88.620 ;
        RECT -41.900 -89.020 -40.540 -88.710 ;
        RECT -38.810 -89.020 -38.670 -88.620 ;
        RECT -33.850 -89.020 -33.710 -88.620 ;
        RECT -31.980 -89.020 -30.620 -88.710 ;
        RECT -28.890 -89.020 -28.750 -88.620 ;
        RECT -23.930 -89.020 -23.790 -88.620 ;
        RECT -22.060 -89.020 -20.700 -88.710 ;
        RECT -18.970 -89.020 -18.830 -88.620 ;
        RECT -14.010 -89.020 -13.870 -88.620 ;
        RECT -12.140 -89.020 -10.780 -88.710 ;
        RECT -9.050 -89.020 -8.910 -88.620 ;
        RECT -4.090 -89.020 -3.950 -88.620 ;
        RECT -2.220 -89.020 -0.860 -88.710 ;
        RECT 0.870 -89.020 1.010 -88.620 ;
        RECT 5.830 -89.020 5.970 -88.620 ;
        RECT 7.700 -89.020 9.060 -88.710 ;
        RECT 10.790 -89.020 10.930 -88.620 ;
        RECT 15.750 -89.020 15.890 -88.620 ;
        RECT 17.620 -89.020 18.980 -88.710 ;
        RECT 20.710 -89.020 20.850 -88.620 ;
        RECT 25.670 -89.020 25.810 -88.620 ;
        RECT 39.270 -88.690 40.110 -87.390 ;
        RECT 34.960 -88.700 40.110 -88.690 ;
        RECT 27.540 -89.020 40.110 -88.700 ;
        RECT -289.000 -89.150 40.110 -89.020 ;
        RECT -289.000 -89.160 36.280 -89.150 ;
        RECT -286.810 -89.560 -286.670 -89.160 ;
        RECT -284.940 -89.470 -283.580 -89.160 ;
        RECT -281.850 -89.560 -281.710 -89.160 ;
        RECT -276.890 -89.560 -276.750 -89.160 ;
        RECT -275.020 -89.470 -273.660 -89.160 ;
        RECT -271.930 -89.560 -271.790 -89.160 ;
        RECT -266.970 -89.560 -266.830 -89.160 ;
        RECT -265.100 -89.470 -263.740 -89.160 ;
        RECT -262.010 -89.560 -261.870 -89.160 ;
        RECT -257.050 -89.560 -256.910 -89.160 ;
        RECT -255.180 -89.470 -253.820 -89.160 ;
        RECT -252.090 -89.560 -251.950 -89.160 ;
        RECT -247.130 -89.560 -246.990 -89.160 ;
        RECT -245.260 -89.470 -243.900 -89.160 ;
        RECT -242.170 -89.560 -242.030 -89.160 ;
        RECT -237.210 -89.560 -237.070 -89.160 ;
        RECT -235.340 -89.470 -233.980 -89.160 ;
        RECT -232.250 -89.560 -232.110 -89.160 ;
        RECT -227.290 -89.560 -227.150 -89.160 ;
        RECT -225.420 -89.470 -224.060 -89.160 ;
        RECT -222.330 -89.560 -222.190 -89.160 ;
        RECT -217.370 -89.560 -217.230 -89.160 ;
        RECT -215.500 -89.470 -214.140 -89.160 ;
        RECT -212.410 -89.560 -212.270 -89.160 ;
        RECT -207.450 -89.560 -207.310 -89.160 ;
        RECT -205.580 -89.470 -204.220 -89.160 ;
        RECT -202.490 -89.560 -202.350 -89.160 ;
        RECT -197.530 -89.560 -197.390 -89.160 ;
        RECT -195.660 -89.470 -194.300 -89.160 ;
        RECT -192.570 -89.560 -192.430 -89.160 ;
        RECT -187.610 -89.560 -187.470 -89.160 ;
        RECT -185.740 -89.470 -184.380 -89.160 ;
        RECT -182.650 -89.560 -182.510 -89.160 ;
        RECT -177.690 -89.560 -177.550 -89.160 ;
        RECT -175.820 -89.470 -174.460 -89.160 ;
        RECT -172.730 -89.560 -172.590 -89.160 ;
        RECT -167.770 -89.560 -167.630 -89.160 ;
        RECT -165.900 -89.470 -164.540 -89.160 ;
        RECT -162.810 -89.560 -162.670 -89.160 ;
        RECT -157.850 -89.560 -157.710 -89.160 ;
        RECT -155.980 -89.470 -154.620 -89.160 ;
        RECT -152.890 -89.560 -152.750 -89.160 ;
        RECT -147.930 -89.560 -147.790 -89.160 ;
        RECT -146.060 -89.470 -144.700 -89.160 ;
        RECT -142.970 -89.560 -142.830 -89.160 ;
        RECT -138.010 -89.560 -137.870 -89.160 ;
        RECT -136.140 -89.470 -134.780 -89.160 ;
        RECT -133.050 -89.560 -132.910 -89.160 ;
        RECT -128.090 -89.560 -127.950 -89.160 ;
        RECT -126.220 -89.470 -124.860 -89.160 ;
        RECT -123.130 -89.560 -122.990 -89.160 ;
        RECT -118.170 -89.560 -118.030 -89.160 ;
        RECT -116.300 -89.470 -114.940 -89.160 ;
        RECT -113.210 -89.560 -113.070 -89.160 ;
        RECT -108.250 -89.560 -108.110 -89.160 ;
        RECT -106.380 -89.470 -105.020 -89.160 ;
        RECT -103.290 -89.560 -103.150 -89.160 ;
        RECT -98.330 -89.560 -98.190 -89.160 ;
        RECT -96.460 -89.470 -95.100 -89.160 ;
        RECT -93.370 -89.560 -93.230 -89.160 ;
        RECT -88.410 -89.560 -88.270 -89.160 ;
        RECT -86.540 -89.470 -85.180 -89.160 ;
        RECT -83.450 -89.560 -83.310 -89.160 ;
        RECT -78.490 -89.560 -78.350 -89.160 ;
        RECT -76.620 -89.470 -75.260 -89.160 ;
        RECT -73.530 -89.560 -73.390 -89.160 ;
        RECT -68.570 -89.560 -68.430 -89.160 ;
        RECT -66.700 -89.470 -65.340 -89.160 ;
        RECT -63.610 -89.560 -63.470 -89.160 ;
        RECT -58.650 -89.560 -58.510 -89.160 ;
        RECT -56.780 -89.470 -55.420 -89.160 ;
        RECT -53.690 -89.560 -53.550 -89.160 ;
        RECT -48.730 -89.560 -48.590 -89.160 ;
        RECT -46.860 -89.470 -45.500 -89.160 ;
        RECT -43.770 -89.560 -43.630 -89.160 ;
        RECT -38.810 -89.560 -38.670 -89.160 ;
        RECT -36.940 -89.470 -35.580 -89.160 ;
        RECT -33.850 -89.560 -33.710 -89.160 ;
        RECT -28.890 -89.560 -28.750 -89.160 ;
        RECT -27.020 -89.470 -25.660 -89.160 ;
        RECT -23.930 -89.560 -23.790 -89.160 ;
        RECT -18.970 -89.560 -18.830 -89.160 ;
        RECT -17.100 -89.470 -15.740 -89.160 ;
        RECT -14.010 -89.560 -13.870 -89.160 ;
        RECT -9.050 -89.560 -8.910 -89.160 ;
        RECT -7.180 -89.470 -5.820 -89.160 ;
        RECT -4.090 -89.560 -3.950 -89.160 ;
        RECT 0.870 -89.560 1.010 -89.160 ;
        RECT 2.740 -89.470 4.100 -89.160 ;
        RECT 5.830 -89.560 5.970 -89.160 ;
        RECT 10.790 -89.560 10.930 -89.160 ;
        RECT 12.660 -89.470 14.020 -89.160 ;
        RECT 15.750 -89.560 15.890 -89.160 ;
        RECT 20.710 -89.560 20.850 -89.160 ;
        RECT 22.580 -89.470 23.940 -89.160 ;
        RECT 25.670 -89.560 25.810 -89.160 ;
        RECT 39.410 -173.860 40.110 -89.150 ;
        RECT -288.750 -176.730 -288.290 -176.420 ;
        RECT -286.560 -176.730 -286.420 -176.330 ;
        RECT -281.600 -176.730 -281.460 -176.330 ;
        RECT -279.730 -176.730 -278.370 -176.420 ;
        RECT -276.640 -176.730 -276.500 -176.330 ;
        RECT -271.680 -176.730 -271.540 -176.330 ;
        RECT -269.810 -176.730 -268.450 -176.420 ;
        RECT -266.720 -176.730 -266.580 -176.330 ;
        RECT -261.760 -176.730 -261.620 -176.330 ;
        RECT -259.890 -176.730 -258.530 -176.420 ;
        RECT -256.800 -176.730 -256.660 -176.330 ;
        RECT -251.840 -176.730 -251.700 -176.330 ;
        RECT -249.970 -176.730 -248.610 -176.420 ;
        RECT -246.880 -176.730 -246.740 -176.330 ;
        RECT -241.920 -176.730 -241.780 -176.330 ;
        RECT -240.050 -176.730 -238.690 -176.420 ;
        RECT -236.960 -176.730 -236.820 -176.330 ;
        RECT -232.000 -176.730 -231.860 -176.330 ;
        RECT -230.130 -176.730 -228.770 -176.420 ;
        RECT -227.040 -176.730 -226.900 -176.330 ;
        RECT -222.080 -176.730 -221.940 -176.330 ;
        RECT -220.210 -176.730 -218.850 -176.420 ;
        RECT -217.120 -176.730 -216.980 -176.330 ;
        RECT -212.160 -176.730 -212.020 -176.330 ;
        RECT -210.290 -176.730 -208.930 -176.420 ;
        RECT -207.200 -176.730 -207.060 -176.330 ;
        RECT -202.240 -176.730 -202.100 -176.330 ;
        RECT -200.370 -176.730 -199.010 -176.420 ;
        RECT -197.280 -176.730 -197.140 -176.330 ;
        RECT -192.320 -176.730 -192.180 -176.330 ;
        RECT -190.450 -176.730 -189.090 -176.420 ;
        RECT -187.360 -176.730 -187.220 -176.330 ;
        RECT -182.400 -176.730 -182.260 -176.330 ;
        RECT -180.530 -176.730 -179.170 -176.420 ;
        RECT -177.440 -176.730 -177.300 -176.330 ;
        RECT -172.480 -176.730 -172.340 -176.330 ;
        RECT -170.610 -176.730 -169.250 -176.420 ;
        RECT -167.520 -176.730 -167.380 -176.330 ;
        RECT -162.560 -176.730 -162.420 -176.330 ;
        RECT -160.690 -176.730 -159.330 -176.420 ;
        RECT -157.600 -176.730 -157.460 -176.330 ;
        RECT -152.640 -176.730 -152.500 -176.330 ;
        RECT -150.770 -176.730 -149.410 -176.420 ;
        RECT -147.680 -176.730 -147.540 -176.330 ;
        RECT -142.720 -176.730 -142.580 -176.330 ;
        RECT -140.850 -176.730 -139.490 -176.420 ;
        RECT -137.760 -176.730 -137.620 -176.330 ;
        RECT -132.800 -176.730 -132.660 -176.330 ;
        RECT -130.930 -176.730 -129.570 -176.420 ;
        RECT -127.840 -176.730 -127.700 -176.330 ;
        RECT -122.880 -176.730 -122.740 -176.330 ;
        RECT -121.010 -176.730 -119.650 -176.420 ;
        RECT -117.920 -176.730 -117.780 -176.330 ;
        RECT -112.960 -176.730 -112.820 -176.330 ;
        RECT -111.090 -176.730 -109.730 -176.420 ;
        RECT -108.000 -176.730 -107.860 -176.330 ;
        RECT -103.040 -176.730 -102.900 -176.330 ;
        RECT -101.170 -176.730 -99.810 -176.420 ;
        RECT -98.080 -176.730 -97.940 -176.330 ;
        RECT -93.120 -176.730 -92.980 -176.330 ;
        RECT -91.250 -176.730 -89.890 -176.420 ;
        RECT -88.160 -176.730 -88.020 -176.330 ;
        RECT -83.200 -176.730 -83.060 -176.330 ;
        RECT -81.330 -176.730 -79.970 -176.420 ;
        RECT -78.240 -176.730 -78.100 -176.330 ;
        RECT -73.280 -176.730 -73.140 -176.330 ;
        RECT -71.410 -176.730 -70.050 -176.420 ;
        RECT -68.320 -176.730 -68.180 -176.330 ;
        RECT -63.360 -176.730 -63.220 -176.330 ;
        RECT -61.490 -176.730 -60.130 -176.420 ;
        RECT -58.400 -176.730 -58.260 -176.330 ;
        RECT -53.440 -176.730 -53.300 -176.330 ;
        RECT -51.570 -176.730 -50.210 -176.420 ;
        RECT -48.480 -176.730 -48.340 -176.330 ;
        RECT -43.520 -176.730 -43.380 -176.330 ;
        RECT -41.650 -176.730 -40.290 -176.420 ;
        RECT -38.560 -176.730 -38.420 -176.330 ;
        RECT -33.600 -176.730 -33.460 -176.330 ;
        RECT -31.730 -176.730 -30.370 -176.420 ;
        RECT -28.640 -176.730 -28.500 -176.330 ;
        RECT -23.680 -176.730 -23.540 -176.330 ;
        RECT -21.810 -176.730 -20.450 -176.420 ;
        RECT -18.720 -176.730 -18.580 -176.330 ;
        RECT -13.760 -176.730 -13.620 -176.330 ;
        RECT -11.890 -176.730 -10.530 -176.420 ;
        RECT -8.800 -176.730 -8.660 -176.330 ;
        RECT -3.840 -176.730 -3.700 -176.330 ;
        RECT -1.970 -176.730 -0.610 -176.420 ;
        RECT 1.120 -176.730 1.260 -176.330 ;
        RECT 6.080 -176.730 6.220 -176.330 ;
        RECT 7.950 -176.730 9.310 -176.420 ;
        RECT 11.040 -176.730 11.180 -176.330 ;
        RECT 16.000 -176.730 16.140 -176.330 ;
        RECT 17.870 -176.730 19.230 -176.420 ;
        RECT 20.960 -176.730 21.100 -176.330 ;
        RECT 25.920 -176.730 26.060 -176.330 ;
        RECT 39.520 -176.400 39.980 -173.860 ;
        RECT 35.210 -176.410 39.980 -176.400 ;
        RECT 27.790 -176.730 39.980 -176.410 ;
        RECT -288.750 -176.860 39.980 -176.730 ;
        RECT -288.750 -176.870 36.530 -176.860 ;
        RECT -286.560 -177.270 -286.420 -176.870 ;
        RECT -284.690 -177.180 -283.330 -176.870 ;
        RECT -281.600 -177.270 -281.460 -176.870 ;
        RECT -276.640 -177.270 -276.500 -176.870 ;
        RECT -274.770 -177.180 -273.410 -176.870 ;
        RECT -271.680 -177.270 -271.540 -176.870 ;
        RECT -266.720 -177.270 -266.580 -176.870 ;
        RECT -264.850 -177.180 -263.490 -176.870 ;
        RECT -261.760 -177.270 -261.620 -176.870 ;
        RECT -256.800 -177.270 -256.660 -176.870 ;
        RECT -254.930 -177.180 -253.570 -176.870 ;
        RECT -251.840 -177.270 -251.700 -176.870 ;
        RECT -246.880 -177.270 -246.740 -176.870 ;
        RECT -245.010 -177.180 -243.650 -176.870 ;
        RECT -241.920 -177.270 -241.780 -176.870 ;
        RECT -236.960 -177.270 -236.820 -176.870 ;
        RECT -235.090 -177.180 -233.730 -176.870 ;
        RECT -232.000 -177.270 -231.860 -176.870 ;
        RECT -227.040 -177.270 -226.900 -176.870 ;
        RECT -225.170 -177.180 -223.810 -176.870 ;
        RECT -222.080 -177.270 -221.940 -176.870 ;
        RECT -217.120 -177.270 -216.980 -176.870 ;
        RECT -215.250 -177.180 -213.890 -176.870 ;
        RECT -212.160 -177.270 -212.020 -176.870 ;
        RECT -207.200 -177.270 -207.060 -176.870 ;
        RECT -205.330 -177.180 -203.970 -176.870 ;
        RECT -202.240 -177.270 -202.100 -176.870 ;
        RECT -197.280 -177.270 -197.140 -176.870 ;
        RECT -195.410 -177.180 -194.050 -176.870 ;
        RECT -192.320 -177.270 -192.180 -176.870 ;
        RECT -187.360 -177.270 -187.220 -176.870 ;
        RECT -185.490 -177.180 -184.130 -176.870 ;
        RECT -182.400 -177.270 -182.260 -176.870 ;
        RECT -177.440 -177.270 -177.300 -176.870 ;
        RECT -175.570 -177.180 -174.210 -176.870 ;
        RECT -172.480 -177.270 -172.340 -176.870 ;
        RECT -167.520 -177.270 -167.380 -176.870 ;
        RECT -165.650 -177.180 -164.290 -176.870 ;
        RECT -162.560 -177.270 -162.420 -176.870 ;
        RECT -157.600 -177.270 -157.460 -176.870 ;
        RECT -155.730 -177.180 -154.370 -176.870 ;
        RECT -152.640 -177.270 -152.500 -176.870 ;
        RECT -147.680 -177.270 -147.540 -176.870 ;
        RECT -145.810 -177.180 -144.450 -176.870 ;
        RECT -142.720 -177.270 -142.580 -176.870 ;
        RECT -137.760 -177.270 -137.620 -176.870 ;
        RECT -135.890 -177.180 -134.530 -176.870 ;
        RECT -132.800 -177.270 -132.660 -176.870 ;
        RECT -127.840 -177.270 -127.700 -176.870 ;
        RECT -125.970 -177.180 -124.610 -176.870 ;
        RECT -122.880 -177.270 -122.740 -176.870 ;
        RECT -117.920 -177.270 -117.780 -176.870 ;
        RECT -116.050 -177.180 -114.690 -176.870 ;
        RECT -112.960 -177.270 -112.820 -176.870 ;
        RECT -108.000 -177.270 -107.860 -176.870 ;
        RECT -106.130 -177.180 -104.770 -176.870 ;
        RECT -103.040 -177.270 -102.900 -176.870 ;
        RECT -98.080 -177.270 -97.940 -176.870 ;
        RECT -96.210 -177.180 -94.850 -176.870 ;
        RECT -93.120 -177.270 -92.980 -176.870 ;
        RECT -88.160 -177.270 -88.020 -176.870 ;
        RECT -86.290 -177.180 -84.930 -176.870 ;
        RECT -83.200 -177.270 -83.060 -176.870 ;
        RECT -78.240 -177.270 -78.100 -176.870 ;
        RECT -76.370 -177.180 -75.010 -176.870 ;
        RECT -73.280 -177.270 -73.140 -176.870 ;
        RECT -68.320 -177.270 -68.180 -176.870 ;
        RECT -66.450 -177.180 -65.090 -176.870 ;
        RECT -63.360 -177.270 -63.220 -176.870 ;
        RECT -58.400 -177.270 -58.260 -176.870 ;
        RECT -56.530 -177.180 -55.170 -176.870 ;
        RECT -53.440 -177.270 -53.300 -176.870 ;
        RECT -48.480 -177.270 -48.340 -176.870 ;
        RECT -46.610 -177.180 -45.250 -176.870 ;
        RECT -43.520 -177.270 -43.380 -176.870 ;
        RECT -38.560 -177.270 -38.420 -176.870 ;
        RECT -36.690 -177.180 -35.330 -176.870 ;
        RECT -33.600 -177.270 -33.460 -176.870 ;
        RECT -28.640 -177.270 -28.500 -176.870 ;
        RECT -26.770 -177.180 -25.410 -176.870 ;
        RECT -23.680 -177.270 -23.540 -176.870 ;
        RECT -18.720 -177.270 -18.580 -176.870 ;
        RECT -16.850 -177.180 -15.490 -176.870 ;
        RECT -13.760 -177.270 -13.620 -176.870 ;
        RECT -8.800 -177.270 -8.660 -176.870 ;
        RECT -6.930 -177.180 -5.570 -176.870 ;
        RECT -3.840 -177.270 -3.700 -176.870 ;
        RECT 1.120 -177.270 1.260 -176.870 ;
        RECT 2.990 -177.180 4.350 -176.870 ;
        RECT 6.080 -177.270 6.220 -176.870 ;
        RECT 11.040 -177.270 11.180 -176.870 ;
        RECT 12.910 -177.180 14.270 -176.870 ;
        RECT 16.000 -177.270 16.140 -176.870 ;
        RECT 20.960 -177.270 21.100 -176.870 ;
        RECT 22.830 -177.180 24.190 -176.870 ;
        RECT 25.920 -177.270 26.060 -176.870 ;
    END
  END i_srclk
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -286.485 93.835 -286.055 94.620 ;
        RECT -276.565 93.835 -276.135 94.620 ;
        RECT -266.645 93.835 -266.215 94.620 ;
        RECT -256.725 93.835 -256.295 94.620 ;
        RECT -246.805 93.835 -246.375 94.620 ;
        RECT -236.885 93.835 -236.455 94.620 ;
        RECT -226.965 93.835 -226.535 94.620 ;
        RECT -217.045 93.835 -216.615 94.620 ;
        RECT -207.125 93.835 -206.695 94.620 ;
        RECT -197.205 93.835 -196.775 94.620 ;
        RECT -187.285 93.835 -186.855 94.620 ;
        RECT -177.365 93.835 -176.935 94.620 ;
        RECT -167.445 93.835 -167.015 94.620 ;
        RECT -157.525 93.835 -157.095 94.620 ;
        RECT -147.605 93.835 -147.175 94.620 ;
        RECT -137.685 93.835 -137.255 94.620 ;
        RECT -127.765 93.835 -127.335 94.620 ;
        RECT -117.845 93.835 -117.415 94.620 ;
        RECT -107.925 93.835 -107.495 94.620 ;
        RECT -98.005 93.835 -97.575 94.620 ;
        RECT -88.085 93.835 -87.655 94.620 ;
        RECT -78.165 93.835 -77.735 94.620 ;
        RECT -68.245 93.835 -67.815 94.620 ;
        RECT -58.325 93.835 -57.895 94.620 ;
        RECT -48.405 93.835 -47.975 94.620 ;
        RECT -38.485 93.835 -38.055 94.620 ;
        RECT -28.565 93.835 -28.135 94.620 ;
        RECT -18.645 93.835 -18.215 94.620 ;
        RECT -8.725 93.835 -8.295 94.620 ;
        RECT 1.195 93.835 1.625 94.620 ;
        RECT 11.115 93.835 11.545 94.620 ;
        RECT 21.035 93.835 21.465 94.620 ;
        RECT -282.915 92.315 -279.705 93.225 ;
        RECT -272.995 92.315 -269.785 93.225 ;
        RECT -263.075 92.315 -259.865 93.225 ;
        RECT -253.155 92.315 -249.945 93.225 ;
        RECT -243.235 92.315 -240.025 93.225 ;
        RECT -233.315 92.315 -230.105 93.225 ;
        RECT -223.395 92.315 -220.185 93.225 ;
        RECT -213.475 92.315 -210.265 93.225 ;
        RECT -203.555 92.315 -200.345 93.225 ;
        RECT -193.635 92.315 -190.425 93.225 ;
        RECT -183.715 92.315 -180.505 93.225 ;
        RECT -173.795 92.315 -170.585 93.225 ;
        RECT -163.875 92.315 -160.665 93.225 ;
        RECT -153.955 92.315 -150.745 93.225 ;
        RECT -144.035 92.315 -140.825 93.225 ;
        RECT -134.115 92.315 -130.905 93.225 ;
        RECT -124.195 92.315 -120.985 93.225 ;
        RECT -114.275 92.315 -111.065 93.225 ;
        RECT -104.355 92.315 -101.145 93.225 ;
        RECT -94.435 92.315 -91.225 93.225 ;
        RECT -84.515 92.315 -81.305 93.225 ;
        RECT -74.595 92.315 -71.385 93.225 ;
        RECT -64.675 92.315 -61.465 93.225 ;
        RECT -54.755 92.315 -51.545 93.225 ;
        RECT -44.835 92.315 -41.625 93.225 ;
        RECT -34.915 92.315 -31.705 93.225 ;
        RECT -24.995 92.315 -21.785 93.225 ;
        RECT -15.075 92.315 -11.865 93.225 ;
        RECT -5.155 92.315 -1.945 93.225 ;
        RECT 4.765 92.315 7.975 93.225 ;
        RECT 14.685 92.315 17.895 93.225 ;
        RECT -287.875 90.715 -284.665 91.625 ;
        RECT -277.955 90.715 -274.745 91.625 ;
        RECT -268.035 90.715 -264.825 91.625 ;
        RECT -258.115 90.715 -254.905 91.625 ;
        RECT -248.195 90.715 -244.985 91.625 ;
        RECT -238.275 90.715 -235.065 91.625 ;
        RECT -228.355 90.715 -225.145 91.625 ;
        RECT -218.435 90.715 -215.225 91.625 ;
        RECT -208.515 90.715 -205.305 91.625 ;
        RECT -198.595 90.715 -195.385 91.625 ;
        RECT -188.675 90.715 -185.465 91.625 ;
        RECT -178.755 90.715 -175.545 91.625 ;
        RECT -168.835 90.715 -165.625 91.625 ;
        RECT -158.915 90.715 -155.705 91.625 ;
        RECT -148.995 90.715 -145.785 91.625 ;
        RECT -139.075 90.715 -135.865 91.625 ;
        RECT -129.155 90.715 -125.945 91.625 ;
        RECT -119.235 90.715 -116.025 91.625 ;
        RECT -109.315 90.715 -106.105 91.625 ;
        RECT -99.395 90.715 -96.185 91.625 ;
        RECT -89.475 90.715 -86.265 91.625 ;
        RECT -79.555 90.715 -76.345 91.625 ;
        RECT -69.635 90.715 -66.425 91.625 ;
        RECT -59.715 90.715 -56.505 91.625 ;
        RECT -49.795 90.715 -46.585 91.625 ;
        RECT -39.875 90.715 -36.665 91.625 ;
        RECT -29.955 90.715 -26.745 91.625 ;
        RECT -20.035 90.715 -16.825 91.625 ;
        RECT -10.115 90.715 -6.905 91.625 ;
        RECT -0.195 90.715 3.015 91.625 ;
        RECT 9.725 90.715 12.935 91.625 ;
        RECT 19.645 90.715 22.855 91.625 ;
        RECT -281.525 89.410 -281.095 90.195 ;
        RECT -271.605 89.410 -271.175 90.195 ;
        RECT -261.685 89.410 -261.255 90.195 ;
        RECT -251.765 89.410 -251.335 90.195 ;
        RECT -241.845 89.410 -241.415 90.195 ;
        RECT -231.925 89.410 -231.495 90.195 ;
        RECT -222.005 89.410 -221.575 90.195 ;
        RECT -212.085 89.410 -211.655 90.195 ;
        RECT -202.165 89.410 -201.735 90.195 ;
        RECT -192.245 89.410 -191.815 90.195 ;
        RECT -182.325 89.410 -181.895 90.195 ;
        RECT -172.405 89.410 -171.975 90.195 ;
        RECT -162.485 89.410 -162.055 90.195 ;
        RECT -152.565 89.410 -152.135 90.195 ;
        RECT -142.645 89.410 -142.215 90.195 ;
        RECT -132.725 89.410 -132.295 90.195 ;
        RECT -122.805 89.410 -122.375 90.195 ;
        RECT -112.885 89.410 -112.455 90.195 ;
        RECT -102.965 89.410 -102.535 90.195 ;
        RECT -93.045 89.410 -92.615 90.195 ;
        RECT -83.125 89.410 -82.695 90.195 ;
        RECT -73.205 89.410 -72.775 90.195 ;
        RECT -63.285 89.410 -62.855 90.195 ;
        RECT -53.365 89.410 -52.935 90.195 ;
        RECT -43.445 89.410 -43.015 90.195 ;
        RECT -33.525 89.410 -33.095 90.195 ;
        RECT -23.605 89.410 -23.175 90.195 ;
        RECT -13.685 89.410 -13.255 90.195 ;
        RECT -3.765 89.410 -3.335 90.195 ;
        RECT 6.155 89.410 6.585 90.195 ;
        RECT 16.075 89.410 16.505 90.195 ;
        RECT -286.235 6.125 -285.805 6.910 ;
        RECT -276.315 6.125 -275.885 6.910 ;
        RECT -266.395 6.125 -265.965 6.910 ;
        RECT -256.475 6.125 -256.045 6.910 ;
        RECT -246.555 6.125 -246.125 6.910 ;
        RECT -236.635 6.125 -236.205 6.910 ;
        RECT -226.715 6.125 -226.285 6.910 ;
        RECT -216.795 6.125 -216.365 6.910 ;
        RECT -206.875 6.125 -206.445 6.910 ;
        RECT -196.955 6.125 -196.525 6.910 ;
        RECT -187.035 6.125 -186.605 6.910 ;
        RECT -177.115 6.125 -176.685 6.910 ;
        RECT -167.195 6.125 -166.765 6.910 ;
        RECT -157.275 6.125 -156.845 6.910 ;
        RECT -147.355 6.125 -146.925 6.910 ;
        RECT -137.435 6.125 -137.005 6.910 ;
        RECT -127.515 6.125 -127.085 6.910 ;
        RECT -117.595 6.125 -117.165 6.910 ;
        RECT -107.675 6.125 -107.245 6.910 ;
        RECT -97.755 6.125 -97.325 6.910 ;
        RECT -87.835 6.125 -87.405 6.910 ;
        RECT -77.915 6.125 -77.485 6.910 ;
        RECT -67.995 6.125 -67.565 6.910 ;
        RECT -58.075 6.125 -57.645 6.910 ;
        RECT -48.155 6.125 -47.725 6.910 ;
        RECT -38.235 6.125 -37.805 6.910 ;
        RECT -28.315 6.125 -27.885 6.910 ;
        RECT -18.395 6.125 -17.965 6.910 ;
        RECT -8.475 6.125 -8.045 6.910 ;
        RECT 1.445 6.125 1.875 6.910 ;
        RECT 11.365 6.125 11.795 6.910 ;
        RECT 21.285 6.125 21.715 6.910 ;
        RECT -282.665 4.605 -279.455 5.515 ;
        RECT -272.745 4.605 -269.535 5.515 ;
        RECT -262.825 4.605 -259.615 5.515 ;
        RECT -252.905 4.605 -249.695 5.515 ;
        RECT -242.985 4.605 -239.775 5.515 ;
        RECT -233.065 4.605 -229.855 5.515 ;
        RECT -223.145 4.605 -219.935 5.515 ;
        RECT -213.225 4.605 -210.015 5.515 ;
        RECT -203.305 4.605 -200.095 5.515 ;
        RECT -193.385 4.605 -190.175 5.515 ;
        RECT -183.465 4.605 -180.255 5.515 ;
        RECT -173.545 4.605 -170.335 5.515 ;
        RECT -163.625 4.605 -160.415 5.515 ;
        RECT -153.705 4.605 -150.495 5.515 ;
        RECT -143.785 4.605 -140.575 5.515 ;
        RECT -133.865 4.605 -130.655 5.515 ;
        RECT -123.945 4.605 -120.735 5.515 ;
        RECT -114.025 4.605 -110.815 5.515 ;
        RECT -104.105 4.605 -100.895 5.515 ;
        RECT -94.185 4.605 -90.975 5.515 ;
        RECT -84.265 4.605 -81.055 5.515 ;
        RECT -74.345 4.605 -71.135 5.515 ;
        RECT -64.425 4.605 -61.215 5.515 ;
        RECT -54.505 4.605 -51.295 5.515 ;
        RECT -44.585 4.605 -41.375 5.515 ;
        RECT -34.665 4.605 -31.455 5.515 ;
        RECT -24.745 4.605 -21.535 5.515 ;
        RECT -14.825 4.605 -11.615 5.515 ;
        RECT -4.905 4.605 -1.695 5.515 ;
        RECT 5.015 4.605 8.225 5.515 ;
        RECT 14.935 4.605 18.145 5.515 ;
        RECT -287.625 3.005 -284.415 3.915 ;
        RECT -277.705 3.005 -274.495 3.915 ;
        RECT -267.785 3.005 -264.575 3.915 ;
        RECT -257.865 3.005 -254.655 3.915 ;
        RECT -247.945 3.005 -244.735 3.915 ;
        RECT -238.025 3.005 -234.815 3.915 ;
        RECT -228.105 3.005 -224.895 3.915 ;
        RECT -218.185 3.005 -214.975 3.915 ;
        RECT -208.265 3.005 -205.055 3.915 ;
        RECT -198.345 3.005 -195.135 3.915 ;
        RECT -188.425 3.005 -185.215 3.915 ;
        RECT -178.505 3.005 -175.295 3.915 ;
        RECT -168.585 3.005 -165.375 3.915 ;
        RECT -158.665 3.005 -155.455 3.915 ;
        RECT -148.745 3.005 -145.535 3.915 ;
        RECT -138.825 3.005 -135.615 3.915 ;
        RECT -128.905 3.005 -125.695 3.915 ;
        RECT -118.985 3.005 -115.775 3.915 ;
        RECT -109.065 3.005 -105.855 3.915 ;
        RECT -99.145 3.005 -95.935 3.915 ;
        RECT -89.225 3.005 -86.015 3.915 ;
        RECT -79.305 3.005 -76.095 3.915 ;
        RECT -69.385 3.005 -66.175 3.915 ;
        RECT -59.465 3.005 -56.255 3.915 ;
        RECT -49.545 3.005 -46.335 3.915 ;
        RECT -39.625 3.005 -36.415 3.915 ;
        RECT -29.705 3.005 -26.495 3.915 ;
        RECT -19.785 3.005 -16.575 3.915 ;
        RECT -9.865 3.005 -6.655 3.915 ;
        RECT 0.055 3.005 3.265 3.915 ;
        RECT 9.975 3.005 13.185 3.915 ;
        RECT 19.895 3.005 23.105 3.915 ;
        RECT -281.275 1.700 -280.845 2.485 ;
        RECT -271.355 1.700 -270.925 2.485 ;
        RECT -261.435 1.700 -261.005 2.485 ;
        RECT -251.515 1.700 -251.085 2.485 ;
        RECT -241.595 1.700 -241.165 2.485 ;
        RECT -231.675 1.700 -231.245 2.485 ;
        RECT -221.755 1.700 -221.325 2.485 ;
        RECT -211.835 1.700 -211.405 2.485 ;
        RECT -201.915 1.700 -201.485 2.485 ;
        RECT -191.995 1.700 -191.565 2.485 ;
        RECT -182.075 1.700 -181.645 2.485 ;
        RECT -172.155 1.700 -171.725 2.485 ;
        RECT -162.235 1.700 -161.805 2.485 ;
        RECT -152.315 1.700 -151.885 2.485 ;
        RECT -142.395 1.700 -141.965 2.485 ;
        RECT -132.475 1.700 -132.045 2.485 ;
        RECT -122.555 1.700 -122.125 2.485 ;
        RECT -112.635 1.700 -112.205 2.485 ;
        RECT -102.715 1.700 -102.285 2.485 ;
        RECT -92.795 1.700 -92.365 2.485 ;
        RECT -82.875 1.700 -82.445 2.485 ;
        RECT -72.955 1.700 -72.525 2.485 ;
        RECT -63.035 1.700 -62.605 2.485 ;
        RECT -53.115 1.700 -52.685 2.485 ;
        RECT -43.195 1.700 -42.765 2.485 ;
        RECT -33.275 1.700 -32.845 2.485 ;
        RECT -23.355 1.700 -22.925 2.485 ;
        RECT -13.435 1.700 -13.005 2.485 ;
        RECT -3.515 1.700 -3.085 2.485 ;
        RECT 6.405 1.700 6.835 2.485 ;
        RECT 16.325 1.700 16.755 2.485 ;
        RECT -284.475 -87.225 -284.045 -86.440 ;
        RECT -274.555 -87.225 -274.125 -86.440 ;
        RECT -264.635 -87.225 -264.205 -86.440 ;
        RECT -254.715 -87.225 -254.285 -86.440 ;
        RECT -244.795 -87.225 -244.365 -86.440 ;
        RECT -234.875 -87.225 -234.445 -86.440 ;
        RECT -224.955 -87.225 -224.525 -86.440 ;
        RECT -215.035 -87.225 -214.605 -86.440 ;
        RECT -205.115 -87.225 -204.685 -86.440 ;
        RECT -195.195 -87.225 -194.765 -86.440 ;
        RECT -185.275 -87.225 -184.845 -86.440 ;
        RECT -175.355 -87.225 -174.925 -86.440 ;
        RECT -165.435 -87.225 -165.005 -86.440 ;
        RECT -155.515 -87.225 -155.085 -86.440 ;
        RECT -145.595 -87.225 -145.165 -86.440 ;
        RECT -135.675 -87.225 -135.245 -86.440 ;
        RECT -125.755 -87.225 -125.325 -86.440 ;
        RECT -115.835 -87.225 -115.405 -86.440 ;
        RECT -105.915 -87.225 -105.485 -86.440 ;
        RECT -95.995 -87.225 -95.565 -86.440 ;
        RECT -86.075 -87.225 -85.645 -86.440 ;
        RECT -76.155 -87.225 -75.725 -86.440 ;
        RECT -66.235 -87.225 -65.805 -86.440 ;
        RECT -56.315 -87.225 -55.885 -86.440 ;
        RECT -46.395 -87.225 -45.965 -86.440 ;
        RECT -36.475 -87.225 -36.045 -86.440 ;
        RECT -26.555 -87.225 -26.125 -86.440 ;
        RECT -16.635 -87.225 -16.205 -86.440 ;
        RECT -6.715 -87.225 -6.285 -86.440 ;
        RECT 3.205 -87.225 3.635 -86.440 ;
        RECT 13.125 -87.225 13.555 -86.440 ;
        RECT 23.045 -87.225 23.475 -86.440 ;
        RECT -280.905 -88.745 -277.695 -87.835 ;
        RECT -270.985 -88.745 -267.775 -87.835 ;
        RECT -261.065 -88.745 -257.855 -87.835 ;
        RECT -251.145 -88.745 -247.935 -87.835 ;
        RECT -241.225 -88.745 -238.015 -87.835 ;
        RECT -231.305 -88.745 -228.095 -87.835 ;
        RECT -221.385 -88.745 -218.175 -87.835 ;
        RECT -211.465 -88.745 -208.255 -87.835 ;
        RECT -201.545 -88.745 -198.335 -87.835 ;
        RECT -191.625 -88.745 -188.415 -87.835 ;
        RECT -181.705 -88.745 -178.495 -87.835 ;
        RECT -171.785 -88.745 -168.575 -87.835 ;
        RECT -161.865 -88.745 -158.655 -87.835 ;
        RECT -151.945 -88.745 -148.735 -87.835 ;
        RECT -142.025 -88.745 -138.815 -87.835 ;
        RECT -132.105 -88.745 -128.895 -87.835 ;
        RECT -122.185 -88.745 -118.975 -87.835 ;
        RECT -112.265 -88.745 -109.055 -87.835 ;
        RECT -102.345 -88.745 -99.135 -87.835 ;
        RECT -92.425 -88.745 -89.215 -87.835 ;
        RECT -82.505 -88.745 -79.295 -87.835 ;
        RECT -72.585 -88.745 -69.375 -87.835 ;
        RECT -62.665 -88.745 -59.455 -87.835 ;
        RECT -52.745 -88.745 -49.535 -87.835 ;
        RECT -42.825 -88.745 -39.615 -87.835 ;
        RECT -32.905 -88.745 -29.695 -87.835 ;
        RECT -22.985 -88.745 -19.775 -87.835 ;
        RECT -13.065 -88.745 -9.855 -87.835 ;
        RECT -3.145 -88.745 0.065 -87.835 ;
        RECT 6.775 -88.745 9.985 -87.835 ;
        RECT 16.695 -88.745 19.905 -87.835 ;
        RECT -285.865 -90.345 -282.655 -89.435 ;
        RECT -275.945 -90.345 -272.735 -89.435 ;
        RECT -266.025 -90.345 -262.815 -89.435 ;
        RECT -256.105 -90.345 -252.895 -89.435 ;
        RECT -246.185 -90.345 -242.975 -89.435 ;
        RECT -236.265 -90.345 -233.055 -89.435 ;
        RECT -226.345 -90.345 -223.135 -89.435 ;
        RECT -216.425 -90.345 -213.215 -89.435 ;
        RECT -206.505 -90.345 -203.295 -89.435 ;
        RECT -196.585 -90.345 -193.375 -89.435 ;
        RECT -186.665 -90.345 -183.455 -89.435 ;
        RECT -176.745 -90.345 -173.535 -89.435 ;
        RECT -166.825 -90.345 -163.615 -89.435 ;
        RECT -156.905 -90.345 -153.695 -89.435 ;
        RECT -146.985 -90.345 -143.775 -89.435 ;
        RECT -137.065 -90.345 -133.855 -89.435 ;
        RECT -127.145 -90.345 -123.935 -89.435 ;
        RECT -117.225 -90.345 -114.015 -89.435 ;
        RECT -107.305 -90.345 -104.095 -89.435 ;
        RECT -97.385 -90.345 -94.175 -89.435 ;
        RECT -87.465 -90.345 -84.255 -89.435 ;
        RECT -77.545 -90.345 -74.335 -89.435 ;
        RECT -67.625 -90.345 -64.415 -89.435 ;
        RECT -57.705 -90.345 -54.495 -89.435 ;
        RECT -47.785 -90.345 -44.575 -89.435 ;
        RECT -37.865 -90.345 -34.655 -89.435 ;
        RECT -27.945 -90.345 -24.735 -89.435 ;
        RECT -18.025 -90.345 -14.815 -89.435 ;
        RECT -8.105 -90.345 -4.895 -89.435 ;
        RECT 1.815 -90.345 5.025 -89.435 ;
        RECT 11.735 -90.345 14.945 -89.435 ;
        RECT 21.655 -90.345 24.865 -89.435 ;
        RECT -279.515 -91.650 -279.085 -90.865 ;
        RECT -269.595 -91.650 -269.165 -90.865 ;
        RECT -259.675 -91.650 -259.245 -90.865 ;
        RECT -249.755 -91.650 -249.325 -90.865 ;
        RECT -239.835 -91.650 -239.405 -90.865 ;
        RECT -229.915 -91.650 -229.485 -90.865 ;
        RECT -219.995 -91.650 -219.565 -90.865 ;
        RECT -210.075 -91.650 -209.645 -90.865 ;
        RECT -200.155 -91.650 -199.725 -90.865 ;
        RECT -190.235 -91.650 -189.805 -90.865 ;
        RECT -180.315 -91.650 -179.885 -90.865 ;
        RECT -170.395 -91.650 -169.965 -90.865 ;
        RECT -160.475 -91.650 -160.045 -90.865 ;
        RECT -150.555 -91.650 -150.125 -90.865 ;
        RECT -140.635 -91.650 -140.205 -90.865 ;
        RECT -130.715 -91.650 -130.285 -90.865 ;
        RECT -120.795 -91.650 -120.365 -90.865 ;
        RECT -110.875 -91.650 -110.445 -90.865 ;
        RECT -100.955 -91.650 -100.525 -90.865 ;
        RECT -91.035 -91.650 -90.605 -90.865 ;
        RECT -81.115 -91.650 -80.685 -90.865 ;
        RECT -71.195 -91.650 -70.765 -90.865 ;
        RECT -61.275 -91.650 -60.845 -90.865 ;
        RECT -51.355 -91.650 -50.925 -90.865 ;
        RECT -41.435 -91.650 -41.005 -90.865 ;
        RECT -31.515 -91.650 -31.085 -90.865 ;
        RECT -21.595 -91.650 -21.165 -90.865 ;
        RECT -11.675 -91.650 -11.245 -90.865 ;
        RECT -1.755 -91.650 -1.325 -90.865 ;
        RECT 8.165 -91.650 8.595 -90.865 ;
        RECT 18.085 -91.650 18.515 -90.865 ;
        RECT -284.225 -174.935 -283.795 -174.150 ;
        RECT -274.305 -174.935 -273.875 -174.150 ;
        RECT -264.385 -174.935 -263.955 -174.150 ;
        RECT -254.465 -174.935 -254.035 -174.150 ;
        RECT -244.545 -174.935 -244.115 -174.150 ;
        RECT -234.625 -174.935 -234.195 -174.150 ;
        RECT -224.705 -174.935 -224.275 -174.150 ;
        RECT -214.785 -174.935 -214.355 -174.150 ;
        RECT -204.865 -174.935 -204.435 -174.150 ;
        RECT -194.945 -174.935 -194.515 -174.150 ;
        RECT -185.025 -174.935 -184.595 -174.150 ;
        RECT -175.105 -174.935 -174.675 -174.150 ;
        RECT -165.185 -174.935 -164.755 -174.150 ;
        RECT -155.265 -174.935 -154.835 -174.150 ;
        RECT -145.345 -174.935 -144.915 -174.150 ;
        RECT -135.425 -174.935 -134.995 -174.150 ;
        RECT -125.505 -174.935 -125.075 -174.150 ;
        RECT -115.585 -174.935 -115.155 -174.150 ;
        RECT -105.665 -174.935 -105.235 -174.150 ;
        RECT -95.745 -174.935 -95.315 -174.150 ;
        RECT -85.825 -174.935 -85.395 -174.150 ;
        RECT -75.905 -174.935 -75.475 -174.150 ;
        RECT -65.985 -174.935 -65.555 -174.150 ;
        RECT -56.065 -174.935 -55.635 -174.150 ;
        RECT -46.145 -174.935 -45.715 -174.150 ;
        RECT -36.225 -174.935 -35.795 -174.150 ;
        RECT -26.305 -174.935 -25.875 -174.150 ;
        RECT -16.385 -174.935 -15.955 -174.150 ;
        RECT -6.465 -174.935 -6.035 -174.150 ;
        RECT 3.455 -174.935 3.885 -174.150 ;
        RECT 13.375 -174.935 13.805 -174.150 ;
        RECT 23.295 -174.935 23.725 -174.150 ;
        RECT -280.655 -176.455 -277.445 -175.545 ;
        RECT -270.735 -176.455 -267.525 -175.545 ;
        RECT -260.815 -176.455 -257.605 -175.545 ;
        RECT -250.895 -176.455 -247.685 -175.545 ;
        RECT -240.975 -176.455 -237.765 -175.545 ;
        RECT -231.055 -176.455 -227.845 -175.545 ;
        RECT -221.135 -176.455 -217.925 -175.545 ;
        RECT -211.215 -176.455 -208.005 -175.545 ;
        RECT -201.295 -176.455 -198.085 -175.545 ;
        RECT -191.375 -176.455 -188.165 -175.545 ;
        RECT -181.455 -176.455 -178.245 -175.545 ;
        RECT -171.535 -176.455 -168.325 -175.545 ;
        RECT -161.615 -176.455 -158.405 -175.545 ;
        RECT -151.695 -176.455 -148.485 -175.545 ;
        RECT -141.775 -176.455 -138.565 -175.545 ;
        RECT -131.855 -176.455 -128.645 -175.545 ;
        RECT -121.935 -176.455 -118.725 -175.545 ;
        RECT -112.015 -176.455 -108.805 -175.545 ;
        RECT -102.095 -176.455 -98.885 -175.545 ;
        RECT -92.175 -176.455 -88.965 -175.545 ;
        RECT -82.255 -176.455 -79.045 -175.545 ;
        RECT -72.335 -176.455 -69.125 -175.545 ;
        RECT -62.415 -176.455 -59.205 -175.545 ;
        RECT -52.495 -176.455 -49.285 -175.545 ;
        RECT -42.575 -176.455 -39.365 -175.545 ;
        RECT -32.655 -176.455 -29.445 -175.545 ;
        RECT -22.735 -176.455 -19.525 -175.545 ;
        RECT -12.815 -176.455 -9.605 -175.545 ;
        RECT -2.895 -176.455 0.315 -175.545 ;
        RECT 7.025 -176.455 10.235 -175.545 ;
        RECT 16.945 -176.455 20.155 -175.545 ;
        RECT -285.615 -178.055 -282.405 -177.145 ;
        RECT -275.695 -178.055 -272.485 -177.145 ;
        RECT -265.775 -178.055 -262.565 -177.145 ;
        RECT -255.855 -178.055 -252.645 -177.145 ;
        RECT -245.935 -178.055 -242.725 -177.145 ;
        RECT -236.015 -178.055 -232.805 -177.145 ;
        RECT -226.095 -178.055 -222.885 -177.145 ;
        RECT -216.175 -178.055 -212.965 -177.145 ;
        RECT -206.255 -178.055 -203.045 -177.145 ;
        RECT -196.335 -178.055 -193.125 -177.145 ;
        RECT -186.415 -178.055 -183.205 -177.145 ;
        RECT -176.495 -178.055 -173.285 -177.145 ;
        RECT -166.575 -178.055 -163.365 -177.145 ;
        RECT -156.655 -178.055 -153.445 -177.145 ;
        RECT -146.735 -178.055 -143.525 -177.145 ;
        RECT -136.815 -178.055 -133.605 -177.145 ;
        RECT -126.895 -178.055 -123.685 -177.145 ;
        RECT -116.975 -178.055 -113.765 -177.145 ;
        RECT -107.055 -178.055 -103.845 -177.145 ;
        RECT -97.135 -178.055 -93.925 -177.145 ;
        RECT -87.215 -178.055 -84.005 -177.145 ;
        RECT -77.295 -178.055 -74.085 -177.145 ;
        RECT -67.375 -178.055 -64.165 -177.145 ;
        RECT -57.455 -178.055 -54.245 -177.145 ;
        RECT -47.535 -178.055 -44.325 -177.145 ;
        RECT -37.615 -178.055 -34.405 -177.145 ;
        RECT -27.695 -178.055 -24.485 -177.145 ;
        RECT -17.775 -178.055 -14.565 -177.145 ;
        RECT -7.855 -178.055 -4.645 -177.145 ;
        RECT 2.065 -178.055 5.275 -177.145 ;
        RECT 11.985 -178.055 15.195 -177.145 ;
        RECT 21.905 -178.055 25.115 -177.145 ;
        RECT -279.265 -179.360 -278.835 -178.575 ;
        RECT -269.345 -179.360 -268.915 -178.575 ;
        RECT -259.425 -179.360 -258.995 -178.575 ;
        RECT -249.505 -179.360 -249.075 -178.575 ;
        RECT -239.585 -179.360 -239.155 -178.575 ;
        RECT -229.665 -179.360 -229.235 -178.575 ;
        RECT -219.745 -179.360 -219.315 -178.575 ;
        RECT -209.825 -179.360 -209.395 -178.575 ;
        RECT -199.905 -179.360 -199.475 -178.575 ;
        RECT -189.985 -179.360 -189.555 -178.575 ;
        RECT -180.065 -179.360 -179.635 -178.575 ;
        RECT -170.145 -179.360 -169.715 -178.575 ;
        RECT -160.225 -179.360 -159.795 -178.575 ;
        RECT -150.305 -179.360 -149.875 -178.575 ;
        RECT -140.385 -179.360 -139.955 -178.575 ;
        RECT -130.465 -179.360 -130.035 -178.575 ;
        RECT -120.545 -179.360 -120.115 -178.575 ;
        RECT -110.625 -179.360 -110.195 -178.575 ;
        RECT -100.705 -179.360 -100.275 -178.575 ;
        RECT -90.785 -179.360 -90.355 -178.575 ;
        RECT -80.865 -179.360 -80.435 -178.575 ;
        RECT -70.945 -179.360 -70.515 -178.575 ;
        RECT -61.025 -179.360 -60.595 -178.575 ;
        RECT -51.105 -179.360 -50.675 -178.575 ;
        RECT -41.185 -179.360 -40.755 -178.575 ;
        RECT -31.265 -179.360 -30.835 -178.575 ;
        RECT -21.345 -179.360 -20.915 -178.575 ;
        RECT -11.425 -179.360 -10.995 -178.575 ;
        RECT -1.505 -179.360 -1.075 -178.575 ;
        RECT 8.415 -179.360 8.845 -178.575 ;
        RECT 18.335 -179.360 18.765 -178.575 ;
      LAYER li1 ;
        RECT -288.125 94.615 -287.955 95.140 ;
        RECT -286.500 94.725 -286.040 94.895 ;
        RECT -288.505 94.285 -287.955 94.615 ;
        RECT -288.125 93.760 -287.955 94.285 ;
        RECT -286.415 94.000 -286.125 94.725 ;
        RECT -284.585 94.615 -284.415 95.140 ;
        RECT -278.205 94.615 -278.035 95.140 ;
        RECT -276.580 94.725 -276.120 94.895 ;
        RECT -284.585 94.285 -284.035 94.615 ;
        RECT -278.585 94.285 -278.035 94.615 ;
        RECT -284.585 93.760 -284.415 94.285 ;
        RECT -278.205 93.760 -278.035 94.285 ;
        RECT -276.495 94.000 -276.205 94.725 ;
        RECT -274.665 94.615 -274.495 95.140 ;
        RECT -268.285 94.615 -268.115 95.140 ;
        RECT -266.660 94.725 -266.200 94.895 ;
        RECT -274.665 94.285 -274.115 94.615 ;
        RECT -268.665 94.285 -268.115 94.615 ;
        RECT -274.665 93.760 -274.495 94.285 ;
        RECT -268.285 93.760 -268.115 94.285 ;
        RECT -266.575 94.000 -266.285 94.725 ;
        RECT -264.745 94.615 -264.575 95.140 ;
        RECT -258.365 94.615 -258.195 95.140 ;
        RECT -256.740 94.725 -256.280 94.895 ;
        RECT -264.745 94.285 -264.195 94.615 ;
        RECT -258.745 94.285 -258.195 94.615 ;
        RECT -264.745 93.760 -264.575 94.285 ;
        RECT -258.365 93.760 -258.195 94.285 ;
        RECT -256.655 94.000 -256.365 94.725 ;
        RECT -254.825 94.615 -254.655 95.140 ;
        RECT -248.445 94.615 -248.275 95.140 ;
        RECT -246.820 94.725 -246.360 94.895 ;
        RECT -254.825 94.285 -254.275 94.615 ;
        RECT -248.825 94.285 -248.275 94.615 ;
        RECT -254.825 93.760 -254.655 94.285 ;
        RECT -248.445 93.760 -248.275 94.285 ;
        RECT -246.735 94.000 -246.445 94.725 ;
        RECT -244.905 94.615 -244.735 95.140 ;
        RECT -238.525 94.615 -238.355 95.140 ;
        RECT -236.900 94.725 -236.440 94.895 ;
        RECT -244.905 94.285 -244.355 94.615 ;
        RECT -238.905 94.285 -238.355 94.615 ;
        RECT -244.905 93.760 -244.735 94.285 ;
        RECT -238.525 93.760 -238.355 94.285 ;
        RECT -236.815 94.000 -236.525 94.725 ;
        RECT -234.985 94.615 -234.815 95.140 ;
        RECT -228.605 94.615 -228.435 95.140 ;
        RECT -226.980 94.725 -226.520 94.895 ;
        RECT -234.985 94.285 -234.435 94.615 ;
        RECT -228.985 94.285 -228.435 94.615 ;
        RECT -234.985 93.760 -234.815 94.285 ;
        RECT -228.605 93.760 -228.435 94.285 ;
        RECT -226.895 94.000 -226.605 94.725 ;
        RECT -225.065 94.615 -224.895 95.140 ;
        RECT -218.685 94.615 -218.515 95.140 ;
        RECT -217.060 94.725 -216.600 94.895 ;
        RECT -225.065 94.285 -224.515 94.615 ;
        RECT -219.065 94.285 -218.515 94.615 ;
        RECT -225.065 93.760 -224.895 94.285 ;
        RECT -218.685 93.760 -218.515 94.285 ;
        RECT -216.975 94.000 -216.685 94.725 ;
        RECT -215.145 94.615 -214.975 95.140 ;
        RECT -208.765 94.615 -208.595 95.140 ;
        RECT -207.140 94.725 -206.680 94.895 ;
        RECT -215.145 94.285 -214.595 94.615 ;
        RECT -209.145 94.285 -208.595 94.615 ;
        RECT -215.145 93.760 -214.975 94.285 ;
        RECT -208.765 93.760 -208.595 94.285 ;
        RECT -207.055 94.000 -206.765 94.725 ;
        RECT -205.225 94.615 -205.055 95.140 ;
        RECT -198.845 94.615 -198.675 95.140 ;
        RECT -197.220 94.725 -196.760 94.895 ;
        RECT -205.225 94.285 -204.675 94.615 ;
        RECT -199.225 94.285 -198.675 94.615 ;
        RECT -205.225 93.760 -205.055 94.285 ;
        RECT -198.845 93.760 -198.675 94.285 ;
        RECT -197.135 94.000 -196.845 94.725 ;
        RECT -195.305 94.615 -195.135 95.140 ;
        RECT -188.925 94.615 -188.755 95.140 ;
        RECT -187.300 94.725 -186.840 94.895 ;
        RECT -195.305 94.285 -194.755 94.615 ;
        RECT -189.305 94.285 -188.755 94.615 ;
        RECT -195.305 93.760 -195.135 94.285 ;
        RECT -188.925 93.760 -188.755 94.285 ;
        RECT -187.215 94.000 -186.925 94.725 ;
        RECT -185.385 94.615 -185.215 95.140 ;
        RECT -179.005 94.615 -178.835 95.140 ;
        RECT -177.380 94.725 -176.920 94.895 ;
        RECT -185.385 94.285 -184.835 94.615 ;
        RECT -179.385 94.285 -178.835 94.615 ;
        RECT -185.385 93.760 -185.215 94.285 ;
        RECT -179.005 93.760 -178.835 94.285 ;
        RECT -177.295 94.000 -177.005 94.725 ;
        RECT -175.465 94.615 -175.295 95.140 ;
        RECT -169.085 94.615 -168.915 95.140 ;
        RECT -167.460 94.725 -167.000 94.895 ;
        RECT -175.465 94.285 -174.915 94.615 ;
        RECT -169.465 94.285 -168.915 94.615 ;
        RECT -175.465 93.760 -175.295 94.285 ;
        RECT -169.085 93.760 -168.915 94.285 ;
        RECT -167.375 94.000 -167.085 94.725 ;
        RECT -165.545 94.615 -165.375 95.140 ;
        RECT -159.165 94.615 -158.995 95.140 ;
        RECT -157.540 94.725 -157.080 94.895 ;
        RECT -165.545 94.285 -164.995 94.615 ;
        RECT -159.545 94.285 -158.995 94.615 ;
        RECT -165.545 93.760 -165.375 94.285 ;
        RECT -159.165 93.760 -158.995 94.285 ;
        RECT -157.455 94.000 -157.165 94.725 ;
        RECT -155.625 94.615 -155.455 95.140 ;
        RECT -149.245 94.615 -149.075 95.140 ;
        RECT -147.620 94.725 -147.160 94.895 ;
        RECT -155.625 94.285 -155.075 94.615 ;
        RECT -149.625 94.285 -149.075 94.615 ;
        RECT -155.625 93.760 -155.455 94.285 ;
        RECT -149.245 93.760 -149.075 94.285 ;
        RECT -147.535 94.000 -147.245 94.725 ;
        RECT -145.705 94.615 -145.535 95.140 ;
        RECT -139.325 94.615 -139.155 95.140 ;
        RECT -137.700 94.725 -137.240 94.895 ;
        RECT -145.705 94.285 -145.155 94.615 ;
        RECT -139.705 94.285 -139.155 94.615 ;
        RECT -145.705 93.760 -145.535 94.285 ;
        RECT -139.325 93.760 -139.155 94.285 ;
        RECT -137.615 94.000 -137.325 94.725 ;
        RECT -135.785 94.615 -135.615 95.140 ;
        RECT -129.405 94.615 -129.235 95.140 ;
        RECT -127.780 94.725 -127.320 94.895 ;
        RECT -135.785 94.285 -135.235 94.615 ;
        RECT -129.785 94.285 -129.235 94.615 ;
        RECT -135.785 93.760 -135.615 94.285 ;
        RECT -129.405 93.760 -129.235 94.285 ;
        RECT -127.695 94.000 -127.405 94.725 ;
        RECT -125.865 94.615 -125.695 95.140 ;
        RECT -119.485 94.615 -119.315 95.140 ;
        RECT -117.860 94.725 -117.400 94.895 ;
        RECT -125.865 94.285 -125.315 94.615 ;
        RECT -119.865 94.285 -119.315 94.615 ;
        RECT -125.865 93.760 -125.695 94.285 ;
        RECT -119.485 93.760 -119.315 94.285 ;
        RECT -117.775 94.000 -117.485 94.725 ;
        RECT -115.945 94.615 -115.775 95.140 ;
        RECT -109.565 94.615 -109.395 95.140 ;
        RECT -107.940 94.725 -107.480 94.895 ;
        RECT -115.945 94.285 -115.395 94.615 ;
        RECT -109.945 94.285 -109.395 94.615 ;
        RECT -115.945 93.760 -115.775 94.285 ;
        RECT -109.565 93.760 -109.395 94.285 ;
        RECT -107.855 94.000 -107.565 94.725 ;
        RECT -106.025 94.615 -105.855 95.140 ;
        RECT -99.645 94.615 -99.475 95.140 ;
        RECT -98.020 94.725 -97.560 94.895 ;
        RECT -106.025 94.285 -105.475 94.615 ;
        RECT -100.025 94.285 -99.475 94.615 ;
        RECT -106.025 93.760 -105.855 94.285 ;
        RECT -99.645 93.760 -99.475 94.285 ;
        RECT -97.935 94.000 -97.645 94.725 ;
        RECT -96.105 94.615 -95.935 95.140 ;
        RECT -89.725 94.615 -89.555 95.140 ;
        RECT -88.100 94.725 -87.640 94.895 ;
        RECT -96.105 94.285 -95.555 94.615 ;
        RECT -90.105 94.285 -89.555 94.615 ;
        RECT -96.105 93.760 -95.935 94.285 ;
        RECT -89.725 93.760 -89.555 94.285 ;
        RECT -88.015 94.000 -87.725 94.725 ;
        RECT -86.185 94.615 -86.015 95.140 ;
        RECT -79.805 94.615 -79.635 95.140 ;
        RECT -78.180 94.725 -77.720 94.895 ;
        RECT -86.185 94.285 -85.635 94.615 ;
        RECT -80.185 94.285 -79.635 94.615 ;
        RECT -86.185 93.760 -86.015 94.285 ;
        RECT -79.805 93.760 -79.635 94.285 ;
        RECT -78.095 94.000 -77.805 94.725 ;
        RECT -76.265 94.615 -76.095 95.140 ;
        RECT -69.885 94.615 -69.715 95.140 ;
        RECT -68.260 94.725 -67.800 94.895 ;
        RECT -76.265 94.285 -75.715 94.615 ;
        RECT -70.265 94.285 -69.715 94.615 ;
        RECT -76.265 93.760 -76.095 94.285 ;
        RECT -69.885 93.760 -69.715 94.285 ;
        RECT -68.175 94.000 -67.885 94.725 ;
        RECT -66.345 94.615 -66.175 95.140 ;
        RECT -59.965 94.615 -59.795 95.140 ;
        RECT -58.340 94.725 -57.880 94.895 ;
        RECT -66.345 94.285 -65.795 94.615 ;
        RECT -60.345 94.285 -59.795 94.615 ;
        RECT -66.345 93.760 -66.175 94.285 ;
        RECT -59.965 93.760 -59.795 94.285 ;
        RECT -58.255 94.000 -57.965 94.725 ;
        RECT -56.425 94.615 -56.255 95.140 ;
        RECT -50.045 94.615 -49.875 95.140 ;
        RECT -48.420 94.725 -47.960 94.895 ;
        RECT -56.425 94.285 -55.875 94.615 ;
        RECT -50.425 94.285 -49.875 94.615 ;
        RECT -56.425 93.760 -56.255 94.285 ;
        RECT -50.045 93.760 -49.875 94.285 ;
        RECT -48.335 94.000 -48.045 94.725 ;
        RECT -46.505 94.615 -46.335 95.140 ;
        RECT -40.125 94.615 -39.955 95.140 ;
        RECT -38.500 94.725 -38.040 94.895 ;
        RECT -46.505 94.285 -45.955 94.615 ;
        RECT -40.505 94.285 -39.955 94.615 ;
        RECT -46.505 93.760 -46.335 94.285 ;
        RECT -40.125 93.760 -39.955 94.285 ;
        RECT -38.415 94.000 -38.125 94.725 ;
        RECT -36.585 94.615 -36.415 95.140 ;
        RECT -30.205 94.615 -30.035 95.140 ;
        RECT -28.580 94.725 -28.120 94.895 ;
        RECT -36.585 94.285 -36.035 94.615 ;
        RECT -30.585 94.285 -30.035 94.615 ;
        RECT -36.585 93.760 -36.415 94.285 ;
        RECT -30.205 93.760 -30.035 94.285 ;
        RECT -28.495 94.000 -28.205 94.725 ;
        RECT -26.665 94.615 -26.495 95.140 ;
        RECT -20.285 94.615 -20.115 95.140 ;
        RECT -18.660 94.725 -18.200 94.895 ;
        RECT -26.665 94.285 -26.115 94.615 ;
        RECT -20.665 94.285 -20.115 94.615 ;
        RECT -26.665 93.760 -26.495 94.285 ;
        RECT -20.285 93.760 -20.115 94.285 ;
        RECT -18.575 94.000 -18.285 94.725 ;
        RECT -16.745 94.615 -16.575 95.140 ;
        RECT -10.365 94.615 -10.195 95.140 ;
        RECT -8.740 94.725 -8.280 94.895 ;
        RECT -16.745 94.285 -16.195 94.615 ;
        RECT -10.745 94.285 -10.195 94.615 ;
        RECT -16.745 93.760 -16.575 94.285 ;
        RECT -10.365 93.760 -10.195 94.285 ;
        RECT -8.655 94.000 -8.365 94.725 ;
        RECT -6.825 94.615 -6.655 95.140 ;
        RECT -0.445 94.615 -0.275 95.140 ;
        RECT 1.180 94.725 1.640 94.895 ;
        RECT -6.825 94.285 -6.275 94.615 ;
        RECT -0.825 94.285 -0.275 94.615 ;
        RECT -6.825 93.760 -6.655 94.285 ;
        RECT -0.445 93.760 -0.275 94.285 ;
        RECT 1.265 94.000 1.555 94.725 ;
        RECT 3.095 94.615 3.265 95.140 ;
        RECT 9.475 94.615 9.645 95.140 ;
        RECT 11.100 94.725 11.560 94.895 ;
        RECT 3.095 94.285 3.645 94.615 ;
        RECT 9.095 94.285 9.645 94.615 ;
        RECT 3.095 93.760 3.265 94.285 ;
        RECT 9.475 93.760 9.645 94.285 ;
        RECT 11.185 94.000 11.475 94.725 ;
        RECT 13.015 94.615 13.185 95.140 ;
        RECT 19.395 94.615 19.565 95.140 ;
        RECT 21.020 94.725 21.480 94.895 ;
        RECT 13.015 94.285 13.565 94.615 ;
        RECT 19.015 94.285 19.565 94.615 ;
        RECT 13.015 93.760 13.185 94.285 ;
        RECT 19.395 93.760 19.565 94.285 ;
        RECT 21.105 94.000 21.395 94.725 ;
        RECT 22.935 94.615 23.105 95.140 ;
        RECT 22.935 94.285 23.485 94.615 ;
        RECT 22.935 93.760 23.105 94.285 ;
        RECT -282.920 93.245 -279.700 93.415 ;
        RECT -273.000 93.245 -269.780 93.415 ;
        RECT -263.080 93.245 -259.860 93.415 ;
        RECT -253.160 93.245 -249.940 93.415 ;
        RECT -243.240 93.245 -240.020 93.415 ;
        RECT -233.320 93.245 -230.100 93.415 ;
        RECT -223.400 93.245 -220.180 93.415 ;
        RECT -213.480 93.245 -210.260 93.415 ;
        RECT -203.560 93.245 -200.340 93.415 ;
        RECT -193.640 93.245 -190.420 93.415 ;
        RECT -183.720 93.245 -180.500 93.415 ;
        RECT -173.800 93.245 -170.580 93.415 ;
        RECT -163.880 93.245 -160.660 93.415 ;
        RECT -153.960 93.245 -150.740 93.415 ;
        RECT -144.040 93.245 -140.820 93.415 ;
        RECT -134.120 93.245 -130.900 93.415 ;
        RECT -124.200 93.245 -120.980 93.415 ;
        RECT -114.280 93.245 -111.060 93.415 ;
        RECT -104.360 93.245 -101.140 93.415 ;
        RECT -94.440 93.245 -91.220 93.415 ;
        RECT -84.520 93.245 -81.300 93.415 ;
        RECT -74.600 93.245 -71.380 93.415 ;
        RECT -64.680 93.245 -61.460 93.415 ;
        RECT -54.760 93.245 -51.540 93.415 ;
        RECT -44.840 93.245 -41.620 93.415 ;
        RECT -34.920 93.245 -31.700 93.415 ;
        RECT -25.000 93.245 -21.780 93.415 ;
        RECT -15.080 93.245 -11.860 93.415 ;
        RECT -5.160 93.245 -1.940 93.415 ;
        RECT 4.760 93.245 7.980 93.415 ;
        RECT 14.680 93.245 17.900 93.415 ;
        RECT -281.935 92.445 -281.625 93.245 ;
        RECT -281.455 92.520 -281.165 93.245 ;
        RECT -280.995 92.445 -280.685 93.245 ;
        RECT -272.015 92.445 -271.705 93.245 ;
        RECT -271.535 92.520 -271.245 93.245 ;
        RECT -271.075 92.445 -270.765 93.245 ;
        RECT -262.095 92.445 -261.785 93.245 ;
        RECT -261.615 92.520 -261.325 93.245 ;
        RECT -261.155 92.445 -260.845 93.245 ;
        RECT -252.175 92.445 -251.865 93.245 ;
        RECT -251.695 92.520 -251.405 93.245 ;
        RECT -251.235 92.445 -250.925 93.245 ;
        RECT -242.255 92.445 -241.945 93.245 ;
        RECT -241.775 92.520 -241.485 93.245 ;
        RECT -241.315 92.445 -241.005 93.245 ;
        RECT -232.335 92.445 -232.025 93.245 ;
        RECT -231.855 92.520 -231.565 93.245 ;
        RECT -231.395 92.445 -231.085 93.245 ;
        RECT -222.415 92.445 -222.105 93.245 ;
        RECT -221.935 92.520 -221.645 93.245 ;
        RECT -221.475 92.445 -221.165 93.245 ;
        RECT -212.495 92.445 -212.185 93.245 ;
        RECT -212.015 92.520 -211.725 93.245 ;
        RECT -211.555 92.445 -211.245 93.245 ;
        RECT -202.575 92.445 -202.265 93.245 ;
        RECT -202.095 92.520 -201.805 93.245 ;
        RECT -201.635 92.445 -201.325 93.245 ;
        RECT -192.655 92.445 -192.345 93.245 ;
        RECT -192.175 92.520 -191.885 93.245 ;
        RECT -191.715 92.445 -191.405 93.245 ;
        RECT -182.735 92.445 -182.425 93.245 ;
        RECT -182.255 92.520 -181.965 93.245 ;
        RECT -181.795 92.445 -181.485 93.245 ;
        RECT -172.815 92.445 -172.505 93.245 ;
        RECT -172.335 92.520 -172.045 93.245 ;
        RECT -171.875 92.445 -171.565 93.245 ;
        RECT -162.895 92.445 -162.585 93.245 ;
        RECT -162.415 92.520 -162.125 93.245 ;
        RECT -161.955 92.445 -161.645 93.245 ;
        RECT -152.975 92.445 -152.665 93.245 ;
        RECT -152.495 92.520 -152.205 93.245 ;
        RECT -152.035 92.445 -151.725 93.245 ;
        RECT -143.055 92.445 -142.745 93.245 ;
        RECT -142.575 92.520 -142.285 93.245 ;
        RECT -142.115 92.445 -141.805 93.245 ;
        RECT -133.135 92.445 -132.825 93.245 ;
        RECT -132.655 92.520 -132.365 93.245 ;
        RECT -132.195 92.445 -131.885 93.245 ;
        RECT -123.215 92.445 -122.905 93.245 ;
        RECT -122.735 92.520 -122.445 93.245 ;
        RECT -122.275 92.445 -121.965 93.245 ;
        RECT -113.295 92.445 -112.985 93.245 ;
        RECT -112.815 92.520 -112.525 93.245 ;
        RECT -112.355 92.445 -112.045 93.245 ;
        RECT -103.375 92.445 -103.065 93.245 ;
        RECT -102.895 92.520 -102.605 93.245 ;
        RECT -102.435 92.445 -102.125 93.245 ;
        RECT -93.455 92.445 -93.145 93.245 ;
        RECT -92.975 92.520 -92.685 93.245 ;
        RECT -92.515 92.445 -92.205 93.245 ;
        RECT -83.535 92.445 -83.225 93.245 ;
        RECT -83.055 92.520 -82.765 93.245 ;
        RECT -82.595 92.445 -82.285 93.245 ;
        RECT -73.615 92.445 -73.305 93.245 ;
        RECT -73.135 92.520 -72.845 93.245 ;
        RECT -72.675 92.445 -72.365 93.245 ;
        RECT -63.695 92.445 -63.385 93.245 ;
        RECT -63.215 92.520 -62.925 93.245 ;
        RECT -62.755 92.445 -62.445 93.245 ;
        RECT -53.775 92.445 -53.465 93.245 ;
        RECT -53.295 92.520 -53.005 93.245 ;
        RECT -52.835 92.445 -52.525 93.245 ;
        RECT -43.855 92.445 -43.545 93.245 ;
        RECT -43.375 92.520 -43.085 93.245 ;
        RECT -42.915 92.445 -42.605 93.245 ;
        RECT -33.935 92.445 -33.625 93.245 ;
        RECT -33.455 92.520 -33.165 93.245 ;
        RECT -32.995 92.445 -32.685 93.245 ;
        RECT -24.015 92.445 -23.705 93.245 ;
        RECT -23.535 92.520 -23.245 93.245 ;
        RECT -23.075 92.445 -22.765 93.245 ;
        RECT -14.095 92.445 -13.785 93.245 ;
        RECT -13.615 92.520 -13.325 93.245 ;
        RECT -13.155 92.445 -12.845 93.245 ;
        RECT -4.175 92.445 -3.865 93.245 ;
        RECT -3.695 92.520 -3.405 93.245 ;
        RECT -3.235 92.445 -2.925 93.245 ;
        RECT 5.745 92.445 6.055 93.245 ;
        RECT 6.225 92.520 6.515 93.245 ;
        RECT 6.685 92.445 6.995 93.245 ;
        RECT 15.665 92.445 15.975 93.245 ;
        RECT 16.145 92.520 16.435 93.245 ;
        RECT 16.605 92.445 16.915 93.245 ;
        RECT -286.895 90.695 -286.585 91.495 ;
        RECT -286.415 90.695 -286.125 91.420 ;
        RECT -285.955 90.695 -285.645 91.495 ;
        RECT -276.975 90.695 -276.665 91.495 ;
        RECT -276.495 90.695 -276.205 91.420 ;
        RECT -276.035 90.695 -275.725 91.495 ;
        RECT -267.055 90.695 -266.745 91.495 ;
        RECT -266.575 90.695 -266.285 91.420 ;
        RECT -266.115 90.695 -265.805 91.495 ;
        RECT -257.135 90.695 -256.825 91.495 ;
        RECT -256.655 90.695 -256.365 91.420 ;
        RECT -256.195 90.695 -255.885 91.495 ;
        RECT -247.215 90.695 -246.905 91.495 ;
        RECT -246.735 90.695 -246.445 91.420 ;
        RECT -246.275 90.695 -245.965 91.495 ;
        RECT -237.295 90.695 -236.985 91.495 ;
        RECT -236.815 90.695 -236.525 91.420 ;
        RECT -236.355 90.695 -236.045 91.495 ;
        RECT -227.375 90.695 -227.065 91.495 ;
        RECT -226.895 90.695 -226.605 91.420 ;
        RECT -226.435 90.695 -226.125 91.495 ;
        RECT -217.455 90.695 -217.145 91.495 ;
        RECT -216.975 90.695 -216.685 91.420 ;
        RECT -216.515 90.695 -216.205 91.495 ;
        RECT -207.535 90.695 -207.225 91.495 ;
        RECT -207.055 90.695 -206.765 91.420 ;
        RECT -206.595 90.695 -206.285 91.495 ;
        RECT -197.615 90.695 -197.305 91.495 ;
        RECT -197.135 90.695 -196.845 91.420 ;
        RECT -196.675 90.695 -196.365 91.495 ;
        RECT -187.695 90.695 -187.385 91.495 ;
        RECT -187.215 90.695 -186.925 91.420 ;
        RECT -186.755 90.695 -186.445 91.495 ;
        RECT -177.775 90.695 -177.465 91.495 ;
        RECT -177.295 90.695 -177.005 91.420 ;
        RECT -176.835 90.695 -176.525 91.495 ;
        RECT -167.855 90.695 -167.545 91.495 ;
        RECT -167.375 90.695 -167.085 91.420 ;
        RECT -166.915 90.695 -166.605 91.495 ;
        RECT -157.935 90.695 -157.625 91.495 ;
        RECT -157.455 90.695 -157.165 91.420 ;
        RECT -156.995 90.695 -156.685 91.495 ;
        RECT -148.015 90.695 -147.705 91.495 ;
        RECT -147.535 90.695 -147.245 91.420 ;
        RECT -147.075 90.695 -146.765 91.495 ;
        RECT -138.095 90.695 -137.785 91.495 ;
        RECT -137.615 90.695 -137.325 91.420 ;
        RECT -137.155 90.695 -136.845 91.495 ;
        RECT -128.175 90.695 -127.865 91.495 ;
        RECT -127.695 90.695 -127.405 91.420 ;
        RECT -127.235 90.695 -126.925 91.495 ;
        RECT -118.255 90.695 -117.945 91.495 ;
        RECT -117.775 90.695 -117.485 91.420 ;
        RECT -117.315 90.695 -117.005 91.495 ;
        RECT -108.335 90.695 -108.025 91.495 ;
        RECT -107.855 90.695 -107.565 91.420 ;
        RECT -107.395 90.695 -107.085 91.495 ;
        RECT -98.415 90.695 -98.105 91.495 ;
        RECT -97.935 90.695 -97.645 91.420 ;
        RECT -97.475 90.695 -97.165 91.495 ;
        RECT -88.495 90.695 -88.185 91.495 ;
        RECT -88.015 90.695 -87.725 91.420 ;
        RECT -87.555 90.695 -87.245 91.495 ;
        RECT -78.575 90.695 -78.265 91.495 ;
        RECT -78.095 90.695 -77.805 91.420 ;
        RECT -77.635 90.695 -77.325 91.495 ;
        RECT -68.655 90.695 -68.345 91.495 ;
        RECT -68.175 90.695 -67.885 91.420 ;
        RECT -67.715 90.695 -67.405 91.495 ;
        RECT -58.735 90.695 -58.425 91.495 ;
        RECT -58.255 90.695 -57.965 91.420 ;
        RECT -57.795 90.695 -57.485 91.495 ;
        RECT -48.815 90.695 -48.505 91.495 ;
        RECT -48.335 90.695 -48.045 91.420 ;
        RECT -47.875 90.695 -47.565 91.495 ;
        RECT -38.895 90.695 -38.585 91.495 ;
        RECT -38.415 90.695 -38.125 91.420 ;
        RECT -37.955 90.695 -37.645 91.495 ;
        RECT -28.975 90.695 -28.665 91.495 ;
        RECT -28.495 90.695 -28.205 91.420 ;
        RECT -28.035 90.695 -27.725 91.495 ;
        RECT -19.055 90.695 -18.745 91.495 ;
        RECT -18.575 90.695 -18.285 91.420 ;
        RECT -18.115 90.695 -17.805 91.495 ;
        RECT -9.135 90.695 -8.825 91.495 ;
        RECT -8.655 90.695 -8.365 91.420 ;
        RECT -8.195 90.695 -7.885 91.495 ;
        RECT 0.785 90.695 1.095 91.495 ;
        RECT 1.265 90.695 1.555 91.420 ;
        RECT 1.725 90.695 2.035 91.495 ;
        RECT 10.705 90.695 11.015 91.495 ;
        RECT 11.185 90.695 11.475 91.420 ;
        RECT 11.645 90.695 11.955 91.495 ;
        RECT 20.625 90.695 20.935 91.495 ;
        RECT 21.105 90.695 21.395 91.420 ;
        RECT 21.565 90.695 21.875 91.495 ;
        RECT -287.880 90.525 -284.660 90.695 ;
        RECT -277.960 90.525 -274.740 90.695 ;
        RECT -268.040 90.525 -264.820 90.695 ;
        RECT -258.120 90.525 -254.900 90.695 ;
        RECT -248.200 90.525 -244.980 90.695 ;
        RECT -238.280 90.525 -235.060 90.695 ;
        RECT -228.360 90.525 -225.140 90.695 ;
        RECT -218.440 90.525 -215.220 90.695 ;
        RECT -208.520 90.525 -205.300 90.695 ;
        RECT -198.600 90.525 -195.380 90.695 ;
        RECT -188.680 90.525 -185.460 90.695 ;
        RECT -178.760 90.525 -175.540 90.695 ;
        RECT -168.840 90.525 -165.620 90.695 ;
        RECT -158.920 90.525 -155.700 90.695 ;
        RECT -149.000 90.525 -145.780 90.695 ;
        RECT -139.080 90.525 -135.860 90.695 ;
        RECT -129.160 90.525 -125.940 90.695 ;
        RECT -119.240 90.525 -116.020 90.695 ;
        RECT -109.320 90.525 -106.100 90.695 ;
        RECT -99.400 90.525 -96.180 90.695 ;
        RECT -89.480 90.525 -86.260 90.695 ;
        RECT -79.560 90.525 -76.340 90.695 ;
        RECT -69.640 90.525 -66.420 90.695 ;
        RECT -59.720 90.525 -56.500 90.695 ;
        RECT -49.800 90.525 -46.580 90.695 ;
        RECT -39.880 90.525 -36.660 90.695 ;
        RECT -29.960 90.525 -26.740 90.695 ;
        RECT -20.040 90.525 -16.820 90.695 ;
        RECT -10.120 90.525 -6.900 90.695 ;
        RECT -0.200 90.525 3.020 90.695 ;
        RECT 9.720 90.525 12.940 90.695 ;
        RECT 19.640 90.525 22.860 90.695 ;
        RECT -283.165 89.655 -282.995 90.180 ;
        RECT -283.545 89.325 -282.995 89.655 ;
        RECT -283.165 88.800 -282.995 89.325 ;
        RECT -281.455 89.305 -281.165 90.030 ;
        RECT -279.625 89.655 -279.455 90.180 ;
        RECT -273.245 89.655 -273.075 90.180 ;
        RECT -279.625 89.325 -279.075 89.655 ;
        RECT -273.625 89.325 -273.075 89.655 ;
        RECT -281.540 89.135 -281.080 89.305 ;
        RECT -279.625 88.800 -279.455 89.325 ;
        RECT -273.245 88.800 -273.075 89.325 ;
        RECT -271.535 89.305 -271.245 90.030 ;
        RECT -269.705 89.655 -269.535 90.180 ;
        RECT -263.325 89.655 -263.155 90.180 ;
        RECT -269.705 89.325 -269.155 89.655 ;
        RECT -263.705 89.325 -263.155 89.655 ;
        RECT -271.620 89.135 -271.160 89.305 ;
        RECT -269.705 88.800 -269.535 89.325 ;
        RECT -263.325 88.800 -263.155 89.325 ;
        RECT -261.615 89.305 -261.325 90.030 ;
        RECT -259.785 89.655 -259.615 90.180 ;
        RECT -253.405 89.655 -253.235 90.180 ;
        RECT -259.785 89.325 -259.235 89.655 ;
        RECT -253.785 89.325 -253.235 89.655 ;
        RECT -261.700 89.135 -261.240 89.305 ;
        RECT -259.785 88.800 -259.615 89.325 ;
        RECT -253.405 88.800 -253.235 89.325 ;
        RECT -251.695 89.305 -251.405 90.030 ;
        RECT -249.865 89.655 -249.695 90.180 ;
        RECT -243.485 89.655 -243.315 90.180 ;
        RECT -249.865 89.325 -249.315 89.655 ;
        RECT -243.865 89.325 -243.315 89.655 ;
        RECT -251.780 89.135 -251.320 89.305 ;
        RECT -249.865 88.800 -249.695 89.325 ;
        RECT -243.485 88.800 -243.315 89.325 ;
        RECT -241.775 89.305 -241.485 90.030 ;
        RECT -239.945 89.655 -239.775 90.180 ;
        RECT -233.565 89.655 -233.395 90.180 ;
        RECT -239.945 89.325 -239.395 89.655 ;
        RECT -233.945 89.325 -233.395 89.655 ;
        RECT -241.860 89.135 -241.400 89.305 ;
        RECT -239.945 88.800 -239.775 89.325 ;
        RECT -233.565 88.800 -233.395 89.325 ;
        RECT -231.855 89.305 -231.565 90.030 ;
        RECT -230.025 89.655 -229.855 90.180 ;
        RECT -223.645 89.655 -223.475 90.180 ;
        RECT -230.025 89.325 -229.475 89.655 ;
        RECT -224.025 89.325 -223.475 89.655 ;
        RECT -231.940 89.135 -231.480 89.305 ;
        RECT -230.025 88.800 -229.855 89.325 ;
        RECT -223.645 88.800 -223.475 89.325 ;
        RECT -221.935 89.305 -221.645 90.030 ;
        RECT -220.105 89.655 -219.935 90.180 ;
        RECT -213.725 89.655 -213.555 90.180 ;
        RECT -220.105 89.325 -219.555 89.655 ;
        RECT -214.105 89.325 -213.555 89.655 ;
        RECT -222.020 89.135 -221.560 89.305 ;
        RECT -220.105 88.800 -219.935 89.325 ;
        RECT -213.725 88.800 -213.555 89.325 ;
        RECT -212.015 89.305 -211.725 90.030 ;
        RECT -210.185 89.655 -210.015 90.180 ;
        RECT -203.805 89.655 -203.635 90.180 ;
        RECT -210.185 89.325 -209.635 89.655 ;
        RECT -204.185 89.325 -203.635 89.655 ;
        RECT -212.100 89.135 -211.640 89.305 ;
        RECT -210.185 88.800 -210.015 89.325 ;
        RECT -203.805 88.800 -203.635 89.325 ;
        RECT -202.095 89.305 -201.805 90.030 ;
        RECT -200.265 89.655 -200.095 90.180 ;
        RECT -193.885 89.655 -193.715 90.180 ;
        RECT -200.265 89.325 -199.715 89.655 ;
        RECT -194.265 89.325 -193.715 89.655 ;
        RECT -202.180 89.135 -201.720 89.305 ;
        RECT -200.265 88.800 -200.095 89.325 ;
        RECT -193.885 88.800 -193.715 89.325 ;
        RECT -192.175 89.305 -191.885 90.030 ;
        RECT -190.345 89.655 -190.175 90.180 ;
        RECT -183.965 89.655 -183.795 90.180 ;
        RECT -190.345 89.325 -189.795 89.655 ;
        RECT -184.345 89.325 -183.795 89.655 ;
        RECT -192.260 89.135 -191.800 89.305 ;
        RECT -190.345 88.800 -190.175 89.325 ;
        RECT -183.965 88.800 -183.795 89.325 ;
        RECT -182.255 89.305 -181.965 90.030 ;
        RECT -180.425 89.655 -180.255 90.180 ;
        RECT -174.045 89.655 -173.875 90.180 ;
        RECT -180.425 89.325 -179.875 89.655 ;
        RECT -174.425 89.325 -173.875 89.655 ;
        RECT -182.340 89.135 -181.880 89.305 ;
        RECT -180.425 88.800 -180.255 89.325 ;
        RECT -174.045 88.800 -173.875 89.325 ;
        RECT -172.335 89.305 -172.045 90.030 ;
        RECT -170.505 89.655 -170.335 90.180 ;
        RECT -164.125 89.655 -163.955 90.180 ;
        RECT -170.505 89.325 -169.955 89.655 ;
        RECT -164.505 89.325 -163.955 89.655 ;
        RECT -172.420 89.135 -171.960 89.305 ;
        RECT -170.505 88.800 -170.335 89.325 ;
        RECT -164.125 88.800 -163.955 89.325 ;
        RECT -162.415 89.305 -162.125 90.030 ;
        RECT -160.585 89.655 -160.415 90.180 ;
        RECT -154.205 89.655 -154.035 90.180 ;
        RECT -160.585 89.325 -160.035 89.655 ;
        RECT -154.585 89.325 -154.035 89.655 ;
        RECT -162.500 89.135 -162.040 89.305 ;
        RECT -160.585 88.800 -160.415 89.325 ;
        RECT -154.205 88.800 -154.035 89.325 ;
        RECT -152.495 89.305 -152.205 90.030 ;
        RECT -150.665 89.655 -150.495 90.180 ;
        RECT -144.285 89.655 -144.115 90.180 ;
        RECT -150.665 89.325 -150.115 89.655 ;
        RECT -144.665 89.325 -144.115 89.655 ;
        RECT -152.580 89.135 -152.120 89.305 ;
        RECT -150.665 88.800 -150.495 89.325 ;
        RECT -144.285 88.800 -144.115 89.325 ;
        RECT -142.575 89.305 -142.285 90.030 ;
        RECT -140.745 89.655 -140.575 90.180 ;
        RECT -134.365 89.655 -134.195 90.180 ;
        RECT -140.745 89.325 -140.195 89.655 ;
        RECT -134.745 89.325 -134.195 89.655 ;
        RECT -142.660 89.135 -142.200 89.305 ;
        RECT -140.745 88.800 -140.575 89.325 ;
        RECT -134.365 88.800 -134.195 89.325 ;
        RECT -132.655 89.305 -132.365 90.030 ;
        RECT -130.825 89.655 -130.655 90.180 ;
        RECT -124.445 89.655 -124.275 90.180 ;
        RECT -130.825 89.325 -130.275 89.655 ;
        RECT -124.825 89.325 -124.275 89.655 ;
        RECT -132.740 89.135 -132.280 89.305 ;
        RECT -130.825 88.800 -130.655 89.325 ;
        RECT -124.445 88.800 -124.275 89.325 ;
        RECT -122.735 89.305 -122.445 90.030 ;
        RECT -120.905 89.655 -120.735 90.180 ;
        RECT -114.525 89.655 -114.355 90.180 ;
        RECT -120.905 89.325 -120.355 89.655 ;
        RECT -114.905 89.325 -114.355 89.655 ;
        RECT -122.820 89.135 -122.360 89.305 ;
        RECT -120.905 88.800 -120.735 89.325 ;
        RECT -114.525 88.800 -114.355 89.325 ;
        RECT -112.815 89.305 -112.525 90.030 ;
        RECT -110.985 89.655 -110.815 90.180 ;
        RECT -104.605 89.655 -104.435 90.180 ;
        RECT -110.985 89.325 -110.435 89.655 ;
        RECT -104.985 89.325 -104.435 89.655 ;
        RECT -112.900 89.135 -112.440 89.305 ;
        RECT -110.985 88.800 -110.815 89.325 ;
        RECT -104.605 88.800 -104.435 89.325 ;
        RECT -102.895 89.305 -102.605 90.030 ;
        RECT -101.065 89.655 -100.895 90.180 ;
        RECT -94.685 89.655 -94.515 90.180 ;
        RECT -101.065 89.325 -100.515 89.655 ;
        RECT -95.065 89.325 -94.515 89.655 ;
        RECT -102.980 89.135 -102.520 89.305 ;
        RECT -101.065 88.800 -100.895 89.325 ;
        RECT -94.685 88.800 -94.515 89.325 ;
        RECT -92.975 89.305 -92.685 90.030 ;
        RECT -91.145 89.655 -90.975 90.180 ;
        RECT -84.765 89.655 -84.595 90.180 ;
        RECT -91.145 89.325 -90.595 89.655 ;
        RECT -85.145 89.325 -84.595 89.655 ;
        RECT -93.060 89.135 -92.600 89.305 ;
        RECT -91.145 88.800 -90.975 89.325 ;
        RECT -84.765 88.800 -84.595 89.325 ;
        RECT -83.055 89.305 -82.765 90.030 ;
        RECT -81.225 89.655 -81.055 90.180 ;
        RECT -74.845 89.655 -74.675 90.180 ;
        RECT -81.225 89.325 -80.675 89.655 ;
        RECT -75.225 89.325 -74.675 89.655 ;
        RECT -83.140 89.135 -82.680 89.305 ;
        RECT -81.225 88.800 -81.055 89.325 ;
        RECT -74.845 88.800 -74.675 89.325 ;
        RECT -73.135 89.305 -72.845 90.030 ;
        RECT -71.305 89.655 -71.135 90.180 ;
        RECT -64.925 89.655 -64.755 90.180 ;
        RECT -71.305 89.325 -70.755 89.655 ;
        RECT -65.305 89.325 -64.755 89.655 ;
        RECT -73.220 89.135 -72.760 89.305 ;
        RECT -71.305 88.800 -71.135 89.325 ;
        RECT -64.925 88.800 -64.755 89.325 ;
        RECT -63.215 89.305 -62.925 90.030 ;
        RECT -61.385 89.655 -61.215 90.180 ;
        RECT -55.005 89.655 -54.835 90.180 ;
        RECT -61.385 89.325 -60.835 89.655 ;
        RECT -55.385 89.325 -54.835 89.655 ;
        RECT -63.300 89.135 -62.840 89.305 ;
        RECT -61.385 88.800 -61.215 89.325 ;
        RECT -55.005 88.800 -54.835 89.325 ;
        RECT -53.295 89.305 -53.005 90.030 ;
        RECT -51.465 89.655 -51.295 90.180 ;
        RECT -45.085 89.655 -44.915 90.180 ;
        RECT -51.465 89.325 -50.915 89.655 ;
        RECT -45.465 89.325 -44.915 89.655 ;
        RECT -53.380 89.135 -52.920 89.305 ;
        RECT -51.465 88.800 -51.295 89.325 ;
        RECT -45.085 88.800 -44.915 89.325 ;
        RECT -43.375 89.305 -43.085 90.030 ;
        RECT -41.545 89.655 -41.375 90.180 ;
        RECT -35.165 89.655 -34.995 90.180 ;
        RECT -41.545 89.325 -40.995 89.655 ;
        RECT -35.545 89.325 -34.995 89.655 ;
        RECT -43.460 89.135 -43.000 89.305 ;
        RECT -41.545 88.800 -41.375 89.325 ;
        RECT -35.165 88.800 -34.995 89.325 ;
        RECT -33.455 89.305 -33.165 90.030 ;
        RECT -31.625 89.655 -31.455 90.180 ;
        RECT -25.245 89.655 -25.075 90.180 ;
        RECT -31.625 89.325 -31.075 89.655 ;
        RECT -25.625 89.325 -25.075 89.655 ;
        RECT -33.540 89.135 -33.080 89.305 ;
        RECT -31.625 88.800 -31.455 89.325 ;
        RECT -25.245 88.800 -25.075 89.325 ;
        RECT -23.535 89.305 -23.245 90.030 ;
        RECT -21.705 89.655 -21.535 90.180 ;
        RECT -15.325 89.655 -15.155 90.180 ;
        RECT -21.705 89.325 -21.155 89.655 ;
        RECT -15.705 89.325 -15.155 89.655 ;
        RECT -23.620 89.135 -23.160 89.305 ;
        RECT -21.705 88.800 -21.535 89.325 ;
        RECT -15.325 88.800 -15.155 89.325 ;
        RECT -13.615 89.305 -13.325 90.030 ;
        RECT -11.785 89.655 -11.615 90.180 ;
        RECT -5.405 89.655 -5.235 90.180 ;
        RECT -11.785 89.325 -11.235 89.655 ;
        RECT -5.785 89.325 -5.235 89.655 ;
        RECT -13.700 89.135 -13.240 89.305 ;
        RECT -11.785 88.800 -11.615 89.325 ;
        RECT -5.405 88.800 -5.235 89.325 ;
        RECT -3.695 89.305 -3.405 90.030 ;
        RECT -1.865 89.655 -1.695 90.180 ;
        RECT 4.515 89.655 4.685 90.180 ;
        RECT -1.865 89.325 -1.315 89.655 ;
        RECT 4.135 89.325 4.685 89.655 ;
        RECT -3.780 89.135 -3.320 89.305 ;
        RECT -1.865 88.800 -1.695 89.325 ;
        RECT 4.515 88.800 4.685 89.325 ;
        RECT 6.225 89.305 6.515 90.030 ;
        RECT 8.055 89.655 8.225 90.180 ;
        RECT 14.435 89.655 14.605 90.180 ;
        RECT 8.055 89.325 8.605 89.655 ;
        RECT 14.055 89.325 14.605 89.655 ;
        RECT 6.140 89.135 6.600 89.305 ;
        RECT 8.055 88.800 8.225 89.325 ;
        RECT 14.435 88.800 14.605 89.325 ;
        RECT 16.145 89.305 16.435 90.030 ;
        RECT 17.975 89.655 18.145 90.180 ;
        RECT 17.975 89.325 18.525 89.655 ;
        RECT 16.060 89.135 16.520 89.305 ;
        RECT 17.975 88.800 18.145 89.325 ;
        RECT -287.875 6.905 -287.705 7.430 ;
        RECT -286.250 7.015 -285.790 7.185 ;
        RECT -288.255 6.575 -287.705 6.905 ;
        RECT -287.875 6.050 -287.705 6.575 ;
        RECT -286.165 6.290 -285.875 7.015 ;
        RECT -284.335 6.905 -284.165 7.430 ;
        RECT -277.955 6.905 -277.785 7.430 ;
        RECT -276.330 7.015 -275.870 7.185 ;
        RECT -284.335 6.575 -283.785 6.905 ;
        RECT -278.335 6.575 -277.785 6.905 ;
        RECT -284.335 6.050 -284.165 6.575 ;
        RECT -277.955 6.050 -277.785 6.575 ;
        RECT -276.245 6.290 -275.955 7.015 ;
        RECT -274.415 6.905 -274.245 7.430 ;
        RECT -268.035 6.905 -267.865 7.430 ;
        RECT -266.410 7.015 -265.950 7.185 ;
        RECT -274.415 6.575 -273.865 6.905 ;
        RECT -268.415 6.575 -267.865 6.905 ;
        RECT -274.415 6.050 -274.245 6.575 ;
        RECT -268.035 6.050 -267.865 6.575 ;
        RECT -266.325 6.290 -266.035 7.015 ;
        RECT -264.495 6.905 -264.325 7.430 ;
        RECT -258.115 6.905 -257.945 7.430 ;
        RECT -256.490 7.015 -256.030 7.185 ;
        RECT -264.495 6.575 -263.945 6.905 ;
        RECT -258.495 6.575 -257.945 6.905 ;
        RECT -264.495 6.050 -264.325 6.575 ;
        RECT -258.115 6.050 -257.945 6.575 ;
        RECT -256.405 6.290 -256.115 7.015 ;
        RECT -254.575 6.905 -254.405 7.430 ;
        RECT -248.195 6.905 -248.025 7.430 ;
        RECT -246.570 7.015 -246.110 7.185 ;
        RECT -254.575 6.575 -254.025 6.905 ;
        RECT -248.575 6.575 -248.025 6.905 ;
        RECT -254.575 6.050 -254.405 6.575 ;
        RECT -248.195 6.050 -248.025 6.575 ;
        RECT -246.485 6.290 -246.195 7.015 ;
        RECT -244.655 6.905 -244.485 7.430 ;
        RECT -238.275 6.905 -238.105 7.430 ;
        RECT -236.650 7.015 -236.190 7.185 ;
        RECT -244.655 6.575 -244.105 6.905 ;
        RECT -238.655 6.575 -238.105 6.905 ;
        RECT -244.655 6.050 -244.485 6.575 ;
        RECT -238.275 6.050 -238.105 6.575 ;
        RECT -236.565 6.290 -236.275 7.015 ;
        RECT -234.735 6.905 -234.565 7.430 ;
        RECT -228.355 6.905 -228.185 7.430 ;
        RECT -226.730 7.015 -226.270 7.185 ;
        RECT -234.735 6.575 -234.185 6.905 ;
        RECT -228.735 6.575 -228.185 6.905 ;
        RECT -234.735 6.050 -234.565 6.575 ;
        RECT -228.355 6.050 -228.185 6.575 ;
        RECT -226.645 6.290 -226.355 7.015 ;
        RECT -224.815 6.905 -224.645 7.430 ;
        RECT -218.435 6.905 -218.265 7.430 ;
        RECT -216.810 7.015 -216.350 7.185 ;
        RECT -224.815 6.575 -224.265 6.905 ;
        RECT -218.815 6.575 -218.265 6.905 ;
        RECT -224.815 6.050 -224.645 6.575 ;
        RECT -218.435 6.050 -218.265 6.575 ;
        RECT -216.725 6.290 -216.435 7.015 ;
        RECT -214.895 6.905 -214.725 7.430 ;
        RECT -208.515 6.905 -208.345 7.430 ;
        RECT -206.890 7.015 -206.430 7.185 ;
        RECT -214.895 6.575 -214.345 6.905 ;
        RECT -208.895 6.575 -208.345 6.905 ;
        RECT -214.895 6.050 -214.725 6.575 ;
        RECT -208.515 6.050 -208.345 6.575 ;
        RECT -206.805 6.290 -206.515 7.015 ;
        RECT -204.975 6.905 -204.805 7.430 ;
        RECT -198.595 6.905 -198.425 7.430 ;
        RECT -196.970 7.015 -196.510 7.185 ;
        RECT -204.975 6.575 -204.425 6.905 ;
        RECT -198.975 6.575 -198.425 6.905 ;
        RECT -204.975 6.050 -204.805 6.575 ;
        RECT -198.595 6.050 -198.425 6.575 ;
        RECT -196.885 6.290 -196.595 7.015 ;
        RECT -195.055 6.905 -194.885 7.430 ;
        RECT -188.675 6.905 -188.505 7.430 ;
        RECT -187.050 7.015 -186.590 7.185 ;
        RECT -195.055 6.575 -194.505 6.905 ;
        RECT -189.055 6.575 -188.505 6.905 ;
        RECT -195.055 6.050 -194.885 6.575 ;
        RECT -188.675 6.050 -188.505 6.575 ;
        RECT -186.965 6.290 -186.675 7.015 ;
        RECT -185.135 6.905 -184.965 7.430 ;
        RECT -178.755 6.905 -178.585 7.430 ;
        RECT -177.130 7.015 -176.670 7.185 ;
        RECT -185.135 6.575 -184.585 6.905 ;
        RECT -179.135 6.575 -178.585 6.905 ;
        RECT -185.135 6.050 -184.965 6.575 ;
        RECT -178.755 6.050 -178.585 6.575 ;
        RECT -177.045 6.290 -176.755 7.015 ;
        RECT -175.215 6.905 -175.045 7.430 ;
        RECT -168.835 6.905 -168.665 7.430 ;
        RECT -167.210 7.015 -166.750 7.185 ;
        RECT -175.215 6.575 -174.665 6.905 ;
        RECT -169.215 6.575 -168.665 6.905 ;
        RECT -175.215 6.050 -175.045 6.575 ;
        RECT -168.835 6.050 -168.665 6.575 ;
        RECT -167.125 6.290 -166.835 7.015 ;
        RECT -165.295 6.905 -165.125 7.430 ;
        RECT -158.915 6.905 -158.745 7.430 ;
        RECT -157.290 7.015 -156.830 7.185 ;
        RECT -165.295 6.575 -164.745 6.905 ;
        RECT -159.295 6.575 -158.745 6.905 ;
        RECT -165.295 6.050 -165.125 6.575 ;
        RECT -158.915 6.050 -158.745 6.575 ;
        RECT -157.205 6.290 -156.915 7.015 ;
        RECT -155.375 6.905 -155.205 7.430 ;
        RECT -148.995 6.905 -148.825 7.430 ;
        RECT -147.370 7.015 -146.910 7.185 ;
        RECT -155.375 6.575 -154.825 6.905 ;
        RECT -149.375 6.575 -148.825 6.905 ;
        RECT -155.375 6.050 -155.205 6.575 ;
        RECT -148.995 6.050 -148.825 6.575 ;
        RECT -147.285 6.290 -146.995 7.015 ;
        RECT -145.455 6.905 -145.285 7.430 ;
        RECT -139.075 6.905 -138.905 7.430 ;
        RECT -137.450 7.015 -136.990 7.185 ;
        RECT -145.455 6.575 -144.905 6.905 ;
        RECT -139.455 6.575 -138.905 6.905 ;
        RECT -145.455 6.050 -145.285 6.575 ;
        RECT -139.075 6.050 -138.905 6.575 ;
        RECT -137.365 6.290 -137.075 7.015 ;
        RECT -135.535 6.905 -135.365 7.430 ;
        RECT -129.155 6.905 -128.985 7.430 ;
        RECT -127.530 7.015 -127.070 7.185 ;
        RECT -135.535 6.575 -134.985 6.905 ;
        RECT -129.535 6.575 -128.985 6.905 ;
        RECT -135.535 6.050 -135.365 6.575 ;
        RECT -129.155 6.050 -128.985 6.575 ;
        RECT -127.445 6.290 -127.155 7.015 ;
        RECT -125.615 6.905 -125.445 7.430 ;
        RECT -119.235 6.905 -119.065 7.430 ;
        RECT -117.610 7.015 -117.150 7.185 ;
        RECT -125.615 6.575 -125.065 6.905 ;
        RECT -119.615 6.575 -119.065 6.905 ;
        RECT -125.615 6.050 -125.445 6.575 ;
        RECT -119.235 6.050 -119.065 6.575 ;
        RECT -117.525 6.290 -117.235 7.015 ;
        RECT -115.695 6.905 -115.525 7.430 ;
        RECT -109.315 6.905 -109.145 7.430 ;
        RECT -107.690 7.015 -107.230 7.185 ;
        RECT -115.695 6.575 -115.145 6.905 ;
        RECT -109.695 6.575 -109.145 6.905 ;
        RECT -115.695 6.050 -115.525 6.575 ;
        RECT -109.315 6.050 -109.145 6.575 ;
        RECT -107.605 6.290 -107.315 7.015 ;
        RECT -105.775 6.905 -105.605 7.430 ;
        RECT -99.395 6.905 -99.225 7.430 ;
        RECT -97.770 7.015 -97.310 7.185 ;
        RECT -105.775 6.575 -105.225 6.905 ;
        RECT -99.775 6.575 -99.225 6.905 ;
        RECT -105.775 6.050 -105.605 6.575 ;
        RECT -99.395 6.050 -99.225 6.575 ;
        RECT -97.685 6.290 -97.395 7.015 ;
        RECT -95.855 6.905 -95.685 7.430 ;
        RECT -89.475 6.905 -89.305 7.430 ;
        RECT -87.850 7.015 -87.390 7.185 ;
        RECT -95.855 6.575 -95.305 6.905 ;
        RECT -89.855 6.575 -89.305 6.905 ;
        RECT -95.855 6.050 -95.685 6.575 ;
        RECT -89.475 6.050 -89.305 6.575 ;
        RECT -87.765 6.290 -87.475 7.015 ;
        RECT -85.935 6.905 -85.765 7.430 ;
        RECT -79.555 6.905 -79.385 7.430 ;
        RECT -77.930 7.015 -77.470 7.185 ;
        RECT -85.935 6.575 -85.385 6.905 ;
        RECT -79.935 6.575 -79.385 6.905 ;
        RECT -85.935 6.050 -85.765 6.575 ;
        RECT -79.555 6.050 -79.385 6.575 ;
        RECT -77.845 6.290 -77.555 7.015 ;
        RECT -76.015 6.905 -75.845 7.430 ;
        RECT -69.635 6.905 -69.465 7.430 ;
        RECT -68.010 7.015 -67.550 7.185 ;
        RECT -76.015 6.575 -75.465 6.905 ;
        RECT -70.015 6.575 -69.465 6.905 ;
        RECT -76.015 6.050 -75.845 6.575 ;
        RECT -69.635 6.050 -69.465 6.575 ;
        RECT -67.925 6.290 -67.635 7.015 ;
        RECT -66.095 6.905 -65.925 7.430 ;
        RECT -59.715 6.905 -59.545 7.430 ;
        RECT -58.090 7.015 -57.630 7.185 ;
        RECT -66.095 6.575 -65.545 6.905 ;
        RECT -60.095 6.575 -59.545 6.905 ;
        RECT -66.095 6.050 -65.925 6.575 ;
        RECT -59.715 6.050 -59.545 6.575 ;
        RECT -58.005 6.290 -57.715 7.015 ;
        RECT -56.175 6.905 -56.005 7.430 ;
        RECT -49.795 6.905 -49.625 7.430 ;
        RECT -48.170 7.015 -47.710 7.185 ;
        RECT -56.175 6.575 -55.625 6.905 ;
        RECT -50.175 6.575 -49.625 6.905 ;
        RECT -56.175 6.050 -56.005 6.575 ;
        RECT -49.795 6.050 -49.625 6.575 ;
        RECT -48.085 6.290 -47.795 7.015 ;
        RECT -46.255 6.905 -46.085 7.430 ;
        RECT -39.875 6.905 -39.705 7.430 ;
        RECT -38.250 7.015 -37.790 7.185 ;
        RECT -46.255 6.575 -45.705 6.905 ;
        RECT -40.255 6.575 -39.705 6.905 ;
        RECT -46.255 6.050 -46.085 6.575 ;
        RECT -39.875 6.050 -39.705 6.575 ;
        RECT -38.165 6.290 -37.875 7.015 ;
        RECT -36.335 6.905 -36.165 7.430 ;
        RECT -29.955 6.905 -29.785 7.430 ;
        RECT -28.330 7.015 -27.870 7.185 ;
        RECT -36.335 6.575 -35.785 6.905 ;
        RECT -30.335 6.575 -29.785 6.905 ;
        RECT -36.335 6.050 -36.165 6.575 ;
        RECT -29.955 6.050 -29.785 6.575 ;
        RECT -28.245 6.290 -27.955 7.015 ;
        RECT -26.415 6.905 -26.245 7.430 ;
        RECT -20.035 6.905 -19.865 7.430 ;
        RECT -18.410 7.015 -17.950 7.185 ;
        RECT -26.415 6.575 -25.865 6.905 ;
        RECT -20.415 6.575 -19.865 6.905 ;
        RECT -26.415 6.050 -26.245 6.575 ;
        RECT -20.035 6.050 -19.865 6.575 ;
        RECT -18.325 6.290 -18.035 7.015 ;
        RECT -16.495 6.905 -16.325 7.430 ;
        RECT -10.115 6.905 -9.945 7.430 ;
        RECT -8.490 7.015 -8.030 7.185 ;
        RECT -16.495 6.575 -15.945 6.905 ;
        RECT -10.495 6.575 -9.945 6.905 ;
        RECT -16.495 6.050 -16.325 6.575 ;
        RECT -10.115 6.050 -9.945 6.575 ;
        RECT -8.405 6.290 -8.115 7.015 ;
        RECT -6.575 6.905 -6.405 7.430 ;
        RECT -0.195 6.905 -0.025 7.430 ;
        RECT 1.430 7.015 1.890 7.185 ;
        RECT -6.575 6.575 -6.025 6.905 ;
        RECT -0.575 6.575 -0.025 6.905 ;
        RECT -6.575 6.050 -6.405 6.575 ;
        RECT -0.195 6.050 -0.025 6.575 ;
        RECT 1.515 6.290 1.805 7.015 ;
        RECT 3.345 6.905 3.515 7.430 ;
        RECT 9.725 6.905 9.895 7.430 ;
        RECT 11.350 7.015 11.810 7.185 ;
        RECT 3.345 6.575 3.895 6.905 ;
        RECT 9.345 6.575 9.895 6.905 ;
        RECT 3.345 6.050 3.515 6.575 ;
        RECT 9.725 6.050 9.895 6.575 ;
        RECT 11.435 6.290 11.725 7.015 ;
        RECT 13.265 6.905 13.435 7.430 ;
        RECT 19.645 6.905 19.815 7.430 ;
        RECT 21.270 7.015 21.730 7.185 ;
        RECT 13.265 6.575 13.815 6.905 ;
        RECT 19.265 6.575 19.815 6.905 ;
        RECT 13.265 6.050 13.435 6.575 ;
        RECT 19.645 6.050 19.815 6.575 ;
        RECT 21.355 6.290 21.645 7.015 ;
        RECT 23.185 6.905 23.355 7.430 ;
        RECT 23.185 6.575 23.735 6.905 ;
        RECT 23.185 6.050 23.355 6.575 ;
        RECT -282.670 5.535 -279.450 5.705 ;
        RECT -272.750 5.535 -269.530 5.705 ;
        RECT -262.830 5.535 -259.610 5.705 ;
        RECT -252.910 5.535 -249.690 5.705 ;
        RECT -242.990 5.535 -239.770 5.705 ;
        RECT -233.070 5.535 -229.850 5.705 ;
        RECT -223.150 5.535 -219.930 5.705 ;
        RECT -213.230 5.535 -210.010 5.705 ;
        RECT -203.310 5.535 -200.090 5.705 ;
        RECT -193.390 5.535 -190.170 5.705 ;
        RECT -183.470 5.535 -180.250 5.705 ;
        RECT -173.550 5.535 -170.330 5.705 ;
        RECT -163.630 5.535 -160.410 5.705 ;
        RECT -153.710 5.535 -150.490 5.705 ;
        RECT -143.790 5.535 -140.570 5.705 ;
        RECT -133.870 5.535 -130.650 5.705 ;
        RECT -123.950 5.535 -120.730 5.705 ;
        RECT -114.030 5.535 -110.810 5.705 ;
        RECT -104.110 5.535 -100.890 5.705 ;
        RECT -94.190 5.535 -90.970 5.705 ;
        RECT -84.270 5.535 -81.050 5.705 ;
        RECT -74.350 5.535 -71.130 5.705 ;
        RECT -64.430 5.535 -61.210 5.705 ;
        RECT -54.510 5.535 -51.290 5.705 ;
        RECT -44.590 5.535 -41.370 5.705 ;
        RECT -34.670 5.535 -31.450 5.705 ;
        RECT -24.750 5.535 -21.530 5.705 ;
        RECT -14.830 5.535 -11.610 5.705 ;
        RECT -4.910 5.535 -1.690 5.705 ;
        RECT 5.010 5.535 8.230 5.705 ;
        RECT 14.930 5.535 18.150 5.705 ;
        RECT -281.685 4.735 -281.375 5.535 ;
        RECT -281.205 4.810 -280.915 5.535 ;
        RECT -280.745 4.735 -280.435 5.535 ;
        RECT -271.765 4.735 -271.455 5.535 ;
        RECT -271.285 4.810 -270.995 5.535 ;
        RECT -270.825 4.735 -270.515 5.535 ;
        RECT -261.845 4.735 -261.535 5.535 ;
        RECT -261.365 4.810 -261.075 5.535 ;
        RECT -260.905 4.735 -260.595 5.535 ;
        RECT -251.925 4.735 -251.615 5.535 ;
        RECT -251.445 4.810 -251.155 5.535 ;
        RECT -250.985 4.735 -250.675 5.535 ;
        RECT -242.005 4.735 -241.695 5.535 ;
        RECT -241.525 4.810 -241.235 5.535 ;
        RECT -241.065 4.735 -240.755 5.535 ;
        RECT -232.085 4.735 -231.775 5.535 ;
        RECT -231.605 4.810 -231.315 5.535 ;
        RECT -231.145 4.735 -230.835 5.535 ;
        RECT -222.165 4.735 -221.855 5.535 ;
        RECT -221.685 4.810 -221.395 5.535 ;
        RECT -221.225 4.735 -220.915 5.535 ;
        RECT -212.245 4.735 -211.935 5.535 ;
        RECT -211.765 4.810 -211.475 5.535 ;
        RECT -211.305 4.735 -210.995 5.535 ;
        RECT -202.325 4.735 -202.015 5.535 ;
        RECT -201.845 4.810 -201.555 5.535 ;
        RECT -201.385 4.735 -201.075 5.535 ;
        RECT -192.405 4.735 -192.095 5.535 ;
        RECT -191.925 4.810 -191.635 5.535 ;
        RECT -191.465 4.735 -191.155 5.535 ;
        RECT -182.485 4.735 -182.175 5.535 ;
        RECT -182.005 4.810 -181.715 5.535 ;
        RECT -181.545 4.735 -181.235 5.535 ;
        RECT -172.565 4.735 -172.255 5.535 ;
        RECT -172.085 4.810 -171.795 5.535 ;
        RECT -171.625 4.735 -171.315 5.535 ;
        RECT -162.645 4.735 -162.335 5.535 ;
        RECT -162.165 4.810 -161.875 5.535 ;
        RECT -161.705 4.735 -161.395 5.535 ;
        RECT -152.725 4.735 -152.415 5.535 ;
        RECT -152.245 4.810 -151.955 5.535 ;
        RECT -151.785 4.735 -151.475 5.535 ;
        RECT -142.805 4.735 -142.495 5.535 ;
        RECT -142.325 4.810 -142.035 5.535 ;
        RECT -141.865 4.735 -141.555 5.535 ;
        RECT -132.885 4.735 -132.575 5.535 ;
        RECT -132.405 4.810 -132.115 5.535 ;
        RECT -131.945 4.735 -131.635 5.535 ;
        RECT -122.965 4.735 -122.655 5.535 ;
        RECT -122.485 4.810 -122.195 5.535 ;
        RECT -122.025 4.735 -121.715 5.535 ;
        RECT -113.045 4.735 -112.735 5.535 ;
        RECT -112.565 4.810 -112.275 5.535 ;
        RECT -112.105 4.735 -111.795 5.535 ;
        RECT -103.125 4.735 -102.815 5.535 ;
        RECT -102.645 4.810 -102.355 5.535 ;
        RECT -102.185 4.735 -101.875 5.535 ;
        RECT -93.205 4.735 -92.895 5.535 ;
        RECT -92.725 4.810 -92.435 5.535 ;
        RECT -92.265 4.735 -91.955 5.535 ;
        RECT -83.285 4.735 -82.975 5.535 ;
        RECT -82.805 4.810 -82.515 5.535 ;
        RECT -82.345 4.735 -82.035 5.535 ;
        RECT -73.365 4.735 -73.055 5.535 ;
        RECT -72.885 4.810 -72.595 5.535 ;
        RECT -72.425 4.735 -72.115 5.535 ;
        RECT -63.445 4.735 -63.135 5.535 ;
        RECT -62.965 4.810 -62.675 5.535 ;
        RECT -62.505 4.735 -62.195 5.535 ;
        RECT -53.525 4.735 -53.215 5.535 ;
        RECT -53.045 4.810 -52.755 5.535 ;
        RECT -52.585 4.735 -52.275 5.535 ;
        RECT -43.605 4.735 -43.295 5.535 ;
        RECT -43.125 4.810 -42.835 5.535 ;
        RECT -42.665 4.735 -42.355 5.535 ;
        RECT -33.685 4.735 -33.375 5.535 ;
        RECT -33.205 4.810 -32.915 5.535 ;
        RECT -32.745 4.735 -32.435 5.535 ;
        RECT -23.765 4.735 -23.455 5.535 ;
        RECT -23.285 4.810 -22.995 5.535 ;
        RECT -22.825 4.735 -22.515 5.535 ;
        RECT -13.845 4.735 -13.535 5.535 ;
        RECT -13.365 4.810 -13.075 5.535 ;
        RECT -12.905 4.735 -12.595 5.535 ;
        RECT -3.925 4.735 -3.615 5.535 ;
        RECT -3.445 4.810 -3.155 5.535 ;
        RECT -2.985 4.735 -2.675 5.535 ;
        RECT 5.995 4.735 6.305 5.535 ;
        RECT 6.475 4.810 6.765 5.535 ;
        RECT 6.935 4.735 7.245 5.535 ;
        RECT 15.915 4.735 16.225 5.535 ;
        RECT 16.395 4.810 16.685 5.535 ;
        RECT 16.855 4.735 17.165 5.535 ;
        RECT -286.645 2.985 -286.335 3.785 ;
        RECT -286.165 2.985 -285.875 3.710 ;
        RECT -285.705 2.985 -285.395 3.785 ;
        RECT -276.725 2.985 -276.415 3.785 ;
        RECT -276.245 2.985 -275.955 3.710 ;
        RECT -275.785 2.985 -275.475 3.785 ;
        RECT -266.805 2.985 -266.495 3.785 ;
        RECT -266.325 2.985 -266.035 3.710 ;
        RECT -265.865 2.985 -265.555 3.785 ;
        RECT -256.885 2.985 -256.575 3.785 ;
        RECT -256.405 2.985 -256.115 3.710 ;
        RECT -255.945 2.985 -255.635 3.785 ;
        RECT -246.965 2.985 -246.655 3.785 ;
        RECT -246.485 2.985 -246.195 3.710 ;
        RECT -246.025 2.985 -245.715 3.785 ;
        RECT -237.045 2.985 -236.735 3.785 ;
        RECT -236.565 2.985 -236.275 3.710 ;
        RECT -236.105 2.985 -235.795 3.785 ;
        RECT -227.125 2.985 -226.815 3.785 ;
        RECT -226.645 2.985 -226.355 3.710 ;
        RECT -226.185 2.985 -225.875 3.785 ;
        RECT -217.205 2.985 -216.895 3.785 ;
        RECT -216.725 2.985 -216.435 3.710 ;
        RECT -216.265 2.985 -215.955 3.785 ;
        RECT -207.285 2.985 -206.975 3.785 ;
        RECT -206.805 2.985 -206.515 3.710 ;
        RECT -206.345 2.985 -206.035 3.785 ;
        RECT -197.365 2.985 -197.055 3.785 ;
        RECT -196.885 2.985 -196.595 3.710 ;
        RECT -196.425 2.985 -196.115 3.785 ;
        RECT -187.445 2.985 -187.135 3.785 ;
        RECT -186.965 2.985 -186.675 3.710 ;
        RECT -186.505 2.985 -186.195 3.785 ;
        RECT -177.525 2.985 -177.215 3.785 ;
        RECT -177.045 2.985 -176.755 3.710 ;
        RECT -176.585 2.985 -176.275 3.785 ;
        RECT -167.605 2.985 -167.295 3.785 ;
        RECT -167.125 2.985 -166.835 3.710 ;
        RECT -166.665 2.985 -166.355 3.785 ;
        RECT -157.685 2.985 -157.375 3.785 ;
        RECT -157.205 2.985 -156.915 3.710 ;
        RECT -156.745 2.985 -156.435 3.785 ;
        RECT -147.765 2.985 -147.455 3.785 ;
        RECT -147.285 2.985 -146.995 3.710 ;
        RECT -146.825 2.985 -146.515 3.785 ;
        RECT -137.845 2.985 -137.535 3.785 ;
        RECT -137.365 2.985 -137.075 3.710 ;
        RECT -136.905 2.985 -136.595 3.785 ;
        RECT -127.925 2.985 -127.615 3.785 ;
        RECT -127.445 2.985 -127.155 3.710 ;
        RECT -126.985 2.985 -126.675 3.785 ;
        RECT -118.005 2.985 -117.695 3.785 ;
        RECT -117.525 2.985 -117.235 3.710 ;
        RECT -117.065 2.985 -116.755 3.785 ;
        RECT -108.085 2.985 -107.775 3.785 ;
        RECT -107.605 2.985 -107.315 3.710 ;
        RECT -107.145 2.985 -106.835 3.785 ;
        RECT -98.165 2.985 -97.855 3.785 ;
        RECT -97.685 2.985 -97.395 3.710 ;
        RECT -97.225 2.985 -96.915 3.785 ;
        RECT -88.245 2.985 -87.935 3.785 ;
        RECT -87.765 2.985 -87.475 3.710 ;
        RECT -87.305 2.985 -86.995 3.785 ;
        RECT -78.325 2.985 -78.015 3.785 ;
        RECT -77.845 2.985 -77.555 3.710 ;
        RECT -77.385 2.985 -77.075 3.785 ;
        RECT -68.405 2.985 -68.095 3.785 ;
        RECT -67.925 2.985 -67.635 3.710 ;
        RECT -67.465 2.985 -67.155 3.785 ;
        RECT -58.485 2.985 -58.175 3.785 ;
        RECT -58.005 2.985 -57.715 3.710 ;
        RECT -57.545 2.985 -57.235 3.785 ;
        RECT -48.565 2.985 -48.255 3.785 ;
        RECT -48.085 2.985 -47.795 3.710 ;
        RECT -47.625 2.985 -47.315 3.785 ;
        RECT -38.645 2.985 -38.335 3.785 ;
        RECT -38.165 2.985 -37.875 3.710 ;
        RECT -37.705 2.985 -37.395 3.785 ;
        RECT -28.725 2.985 -28.415 3.785 ;
        RECT -28.245 2.985 -27.955 3.710 ;
        RECT -27.785 2.985 -27.475 3.785 ;
        RECT -18.805 2.985 -18.495 3.785 ;
        RECT -18.325 2.985 -18.035 3.710 ;
        RECT -17.865 2.985 -17.555 3.785 ;
        RECT -8.885 2.985 -8.575 3.785 ;
        RECT -8.405 2.985 -8.115 3.710 ;
        RECT -7.945 2.985 -7.635 3.785 ;
        RECT 1.035 2.985 1.345 3.785 ;
        RECT 1.515 2.985 1.805 3.710 ;
        RECT 1.975 2.985 2.285 3.785 ;
        RECT 10.955 2.985 11.265 3.785 ;
        RECT 11.435 2.985 11.725 3.710 ;
        RECT 11.895 2.985 12.205 3.785 ;
        RECT 20.875 2.985 21.185 3.785 ;
        RECT 21.355 2.985 21.645 3.710 ;
        RECT 21.815 2.985 22.125 3.785 ;
        RECT -287.630 2.815 -284.410 2.985 ;
        RECT -277.710 2.815 -274.490 2.985 ;
        RECT -267.790 2.815 -264.570 2.985 ;
        RECT -257.870 2.815 -254.650 2.985 ;
        RECT -247.950 2.815 -244.730 2.985 ;
        RECT -238.030 2.815 -234.810 2.985 ;
        RECT -228.110 2.815 -224.890 2.985 ;
        RECT -218.190 2.815 -214.970 2.985 ;
        RECT -208.270 2.815 -205.050 2.985 ;
        RECT -198.350 2.815 -195.130 2.985 ;
        RECT -188.430 2.815 -185.210 2.985 ;
        RECT -178.510 2.815 -175.290 2.985 ;
        RECT -168.590 2.815 -165.370 2.985 ;
        RECT -158.670 2.815 -155.450 2.985 ;
        RECT -148.750 2.815 -145.530 2.985 ;
        RECT -138.830 2.815 -135.610 2.985 ;
        RECT -128.910 2.815 -125.690 2.985 ;
        RECT -118.990 2.815 -115.770 2.985 ;
        RECT -109.070 2.815 -105.850 2.985 ;
        RECT -99.150 2.815 -95.930 2.985 ;
        RECT -89.230 2.815 -86.010 2.985 ;
        RECT -79.310 2.815 -76.090 2.985 ;
        RECT -69.390 2.815 -66.170 2.985 ;
        RECT -59.470 2.815 -56.250 2.985 ;
        RECT -49.550 2.815 -46.330 2.985 ;
        RECT -39.630 2.815 -36.410 2.985 ;
        RECT -29.710 2.815 -26.490 2.985 ;
        RECT -19.790 2.815 -16.570 2.985 ;
        RECT -9.870 2.815 -6.650 2.985 ;
        RECT 0.050 2.815 3.270 2.985 ;
        RECT 9.970 2.815 13.190 2.985 ;
        RECT 19.890 2.815 23.110 2.985 ;
        RECT -282.915 1.945 -282.745 2.470 ;
        RECT -283.295 1.615 -282.745 1.945 ;
        RECT -282.915 1.090 -282.745 1.615 ;
        RECT -281.205 1.595 -280.915 2.320 ;
        RECT -279.375 1.945 -279.205 2.470 ;
        RECT -272.995 1.945 -272.825 2.470 ;
        RECT -279.375 1.615 -278.825 1.945 ;
        RECT -273.375 1.615 -272.825 1.945 ;
        RECT -281.290 1.425 -280.830 1.595 ;
        RECT -279.375 1.090 -279.205 1.615 ;
        RECT -272.995 1.090 -272.825 1.615 ;
        RECT -271.285 1.595 -270.995 2.320 ;
        RECT -269.455 1.945 -269.285 2.470 ;
        RECT -263.075 1.945 -262.905 2.470 ;
        RECT -269.455 1.615 -268.905 1.945 ;
        RECT -263.455 1.615 -262.905 1.945 ;
        RECT -271.370 1.425 -270.910 1.595 ;
        RECT -269.455 1.090 -269.285 1.615 ;
        RECT -263.075 1.090 -262.905 1.615 ;
        RECT -261.365 1.595 -261.075 2.320 ;
        RECT -259.535 1.945 -259.365 2.470 ;
        RECT -253.155 1.945 -252.985 2.470 ;
        RECT -259.535 1.615 -258.985 1.945 ;
        RECT -253.535 1.615 -252.985 1.945 ;
        RECT -261.450 1.425 -260.990 1.595 ;
        RECT -259.535 1.090 -259.365 1.615 ;
        RECT -253.155 1.090 -252.985 1.615 ;
        RECT -251.445 1.595 -251.155 2.320 ;
        RECT -249.615 1.945 -249.445 2.470 ;
        RECT -243.235 1.945 -243.065 2.470 ;
        RECT -249.615 1.615 -249.065 1.945 ;
        RECT -243.615 1.615 -243.065 1.945 ;
        RECT -251.530 1.425 -251.070 1.595 ;
        RECT -249.615 1.090 -249.445 1.615 ;
        RECT -243.235 1.090 -243.065 1.615 ;
        RECT -241.525 1.595 -241.235 2.320 ;
        RECT -239.695 1.945 -239.525 2.470 ;
        RECT -233.315 1.945 -233.145 2.470 ;
        RECT -239.695 1.615 -239.145 1.945 ;
        RECT -233.695 1.615 -233.145 1.945 ;
        RECT -241.610 1.425 -241.150 1.595 ;
        RECT -239.695 1.090 -239.525 1.615 ;
        RECT -233.315 1.090 -233.145 1.615 ;
        RECT -231.605 1.595 -231.315 2.320 ;
        RECT -229.775 1.945 -229.605 2.470 ;
        RECT -223.395 1.945 -223.225 2.470 ;
        RECT -229.775 1.615 -229.225 1.945 ;
        RECT -223.775 1.615 -223.225 1.945 ;
        RECT -231.690 1.425 -231.230 1.595 ;
        RECT -229.775 1.090 -229.605 1.615 ;
        RECT -223.395 1.090 -223.225 1.615 ;
        RECT -221.685 1.595 -221.395 2.320 ;
        RECT -219.855 1.945 -219.685 2.470 ;
        RECT -213.475 1.945 -213.305 2.470 ;
        RECT -219.855 1.615 -219.305 1.945 ;
        RECT -213.855 1.615 -213.305 1.945 ;
        RECT -221.770 1.425 -221.310 1.595 ;
        RECT -219.855 1.090 -219.685 1.615 ;
        RECT -213.475 1.090 -213.305 1.615 ;
        RECT -211.765 1.595 -211.475 2.320 ;
        RECT -209.935 1.945 -209.765 2.470 ;
        RECT -203.555 1.945 -203.385 2.470 ;
        RECT -209.935 1.615 -209.385 1.945 ;
        RECT -203.935 1.615 -203.385 1.945 ;
        RECT -211.850 1.425 -211.390 1.595 ;
        RECT -209.935 1.090 -209.765 1.615 ;
        RECT -203.555 1.090 -203.385 1.615 ;
        RECT -201.845 1.595 -201.555 2.320 ;
        RECT -200.015 1.945 -199.845 2.470 ;
        RECT -193.635 1.945 -193.465 2.470 ;
        RECT -200.015 1.615 -199.465 1.945 ;
        RECT -194.015 1.615 -193.465 1.945 ;
        RECT -201.930 1.425 -201.470 1.595 ;
        RECT -200.015 1.090 -199.845 1.615 ;
        RECT -193.635 1.090 -193.465 1.615 ;
        RECT -191.925 1.595 -191.635 2.320 ;
        RECT -190.095 1.945 -189.925 2.470 ;
        RECT -183.715 1.945 -183.545 2.470 ;
        RECT -190.095 1.615 -189.545 1.945 ;
        RECT -184.095 1.615 -183.545 1.945 ;
        RECT -192.010 1.425 -191.550 1.595 ;
        RECT -190.095 1.090 -189.925 1.615 ;
        RECT -183.715 1.090 -183.545 1.615 ;
        RECT -182.005 1.595 -181.715 2.320 ;
        RECT -180.175 1.945 -180.005 2.470 ;
        RECT -173.795 1.945 -173.625 2.470 ;
        RECT -180.175 1.615 -179.625 1.945 ;
        RECT -174.175 1.615 -173.625 1.945 ;
        RECT -182.090 1.425 -181.630 1.595 ;
        RECT -180.175 1.090 -180.005 1.615 ;
        RECT -173.795 1.090 -173.625 1.615 ;
        RECT -172.085 1.595 -171.795 2.320 ;
        RECT -170.255 1.945 -170.085 2.470 ;
        RECT -163.875 1.945 -163.705 2.470 ;
        RECT -170.255 1.615 -169.705 1.945 ;
        RECT -164.255 1.615 -163.705 1.945 ;
        RECT -172.170 1.425 -171.710 1.595 ;
        RECT -170.255 1.090 -170.085 1.615 ;
        RECT -163.875 1.090 -163.705 1.615 ;
        RECT -162.165 1.595 -161.875 2.320 ;
        RECT -160.335 1.945 -160.165 2.470 ;
        RECT -153.955 1.945 -153.785 2.470 ;
        RECT -160.335 1.615 -159.785 1.945 ;
        RECT -154.335 1.615 -153.785 1.945 ;
        RECT -162.250 1.425 -161.790 1.595 ;
        RECT -160.335 1.090 -160.165 1.615 ;
        RECT -153.955 1.090 -153.785 1.615 ;
        RECT -152.245 1.595 -151.955 2.320 ;
        RECT -150.415 1.945 -150.245 2.470 ;
        RECT -144.035 1.945 -143.865 2.470 ;
        RECT -150.415 1.615 -149.865 1.945 ;
        RECT -144.415 1.615 -143.865 1.945 ;
        RECT -152.330 1.425 -151.870 1.595 ;
        RECT -150.415 1.090 -150.245 1.615 ;
        RECT -144.035 1.090 -143.865 1.615 ;
        RECT -142.325 1.595 -142.035 2.320 ;
        RECT -140.495 1.945 -140.325 2.470 ;
        RECT -134.115 1.945 -133.945 2.470 ;
        RECT -140.495 1.615 -139.945 1.945 ;
        RECT -134.495 1.615 -133.945 1.945 ;
        RECT -142.410 1.425 -141.950 1.595 ;
        RECT -140.495 1.090 -140.325 1.615 ;
        RECT -134.115 1.090 -133.945 1.615 ;
        RECT -132.405 1.595 -132.115 2.320 ;
        RECT -130.575 1.945 -130.405 2.470 ;
        RECT -124.195 1.945 -124.025 2.470 ;
        RECT -130.575 1.615 -130.025 1.945 ;
        RECT -124.575 1.615 -124.025 1.945 ;
        RECT -132.490 1.425 -132.030 1.595 ;
        RECT -130.575 1.090 -130.405 1.615 ;
        RECT -124.195 1.090 -124.025 1.615 ;
        RECT -122.485 1.595 -122.195 2.320 ;
        RECT -120.655 1.945 -120.485 2.470 ;
        RECT -114.275 1.945 -114.105 2.470 ;
        RECT -120.655 1.615 -120.105 1.945 ;
        RECT -114.655 1.615 -114.105 1.945 ;
        RECT -122.570 1.425 -122.110 1.595 ;
        RECT -120.655 1.090 -120.485 1.615 ;
        RECT -114.275 1.090 -114.105 1.615 ;
        RECT -112.565 1.595 -112.275 2.320 ;
        RECT -110.735 1.945 -110.565 2.470 ;
        RECT -104.355 1.945 -104.185 2.470 ;
        RECT -110.735 1.615 -110.185 1.945 ;
        RECT -104.735 1.615 -104.185 1.945 ;
        RECT -112.650 1.425 -112.190 1.595 ;
        RECT -110.735 1.090 -110.565 1.615 ;
        RECT -104.355 1.090 -104.185 1.615 ;
        RECT -102.645 1.595 -102.355 2.320 ;
        RECT -100.815 1.945 -100.645 2.470 ;
        RECT -94.435 1.945 -94.265 2.470 ;
        RECT -100.815 1.615 -100.265 1.945 ;
        RECT -94.815 1.615 -94.265 1.945 ;
        RECT -102.730 1.425 -102.270 1.595 ;
        RECT -100.815 1.090 -100.645 1.615 ;
        RECT -94.435 1.090 -94.265 1.615 ;
        RECT -92.725 1.595 -92.435 2.320 ;
        RECT -90.895 1.945 -90.725 2.470 ;
        RECT -84.515 1.945 -84.345 2.470 ;
        RECT -90.895 1.615 -90.345 1.945 ;
        RECT -84.895 1.615 -84.345 1.945 ;
        RECT -92.810 1.425 -92.350 1.595 ;
        RECT -90.895 1.090 -90.725 1.615 ;
        RECT -84.515 1.090 -84.345 1.615 ;
        RECT -82.805 1.595 -82.515 2.320 ;
        RECT -80.975 1.945 -80.805 2.470 ;
        RECT -74.595 1.945 -74.425 2.470 ;
        RECT -80.975 1.615 -80.425 1.945 ;
        RECT -74.975 1.615 -74.425 1.945 ;
        RECT -82.890 1.425 -82.430 1.595 ;
        RECT -80.975 1.090 -80.805 1.615 ;
        RECT -74.595 1.090 -74.425 1.615 ;
        RECT -72.885 1.595 -72.595 2.320 ;
        RECT -71.055 1.945 -70.885 2.470 ;
        RECT -64.675 1.945 -64.505 2.470 ;
        RECT -71.055 1.615 -70.505 1.945 ;
        RECT -65.055 1.615 -64.505 1.945 ;
        RECT -72.970 1.425 -72.510 1.595 ;
        RECT -71.055 1.090 -70.885 1.615 ;
        RECT -64.675 1.090 -64.505 1.615 ;
        RECT -62.965 1.595 -62.675 2.320 ;
        RECT -61.135 1.945 -60.965 2.470 ;
        RECT -54.755 1.945 -54.585 2.470 ;
        RECT -61.135 1.615 -60.585 1.945 ;
        RECT -55.135 1.615 -54.585 1.945 ;
        RECT -63.050 1.425 -62.590 1.595 ;
        RECT -61.135 1.090 -60.965 1.615 ;
        RECT -54.755 1.090 -54.585 1.615 ;
        RECT -53.045 1.595 -52.755 2.320 ;
        RECT -51.215 1.945 -51.045 2.470 ;
        RECT -44.835 1.945 -44.665 2.470 ;
        RECT -51.215 1.615 -50.665 1.945 ;
        RECT -45.215 1.615 -44.665 1.945 ;
        RECT -53.130 1.425 -52.670 1.595 ;
        RECT -51.215 1.090 -51.045 1.615 ;
        RECT -44.835 1.090 -44.665 1.615 ;
        RECT -43.125 1.595 -42.835 2.320 ;
        RECT -41.295 1.945 -41.125 2.470 ;
        RECT -34.915 1.945 -34.745 2.470 ;
        RECT -41.295 1.615 -40.745 1.945 ;
        RECT -35.295 1.615 -34.745 1.945 ;
        RECT -43.210 1.425 -42.750 1.595 ;
        RECT -41.295 1.090 -41.125 1.615 ;
        RECT -34.915 1.090 -34.745 1.615 ;
        RECT -33.205 1.595 -32.915 2.320 ;
        RECT -31.375 1.945 -31.205 2.470 ;
        RECT -24.995 1.945 -24.825 2.470 ;
        RECT -31.375 1.615 -30.825 1.945 ;
        RECT -25.375 1.615 -24.825 1.945 ;
        RECT -33.290 1.425 -32.830 1.595 ;
        RECT -31.375 1.090 -31.205 1.615 ;
        RECT -24.995 1.090 -24.825 1.615 ;
        RECT -23.285 1.595 -22.995 2.320 ;
        RECT -21.455 1.945 -21.285 2.470 ;
        RECT -15.075 1.945 -14.905 2.470 ;
        RECT -21.455 1.615 -20.905 1.945 ;
        RECT -15.455 1.615 -14.905 1.945 ;
        RECT -23.370 1.425 -22.910 1.595 ;
        RECT -21.455 1.090 -21.285 1.615 ;
        RECT -15.075 1.090 -14.905 1.615 ;
        RECT -13.365 1.595 -13.075 2.320 ;
        RECT -11.535 1.945 -11.365 2.470 ;
        RECT -5.155 1.945 -4.985 2.470 ;
        RECT -11.535 1.615 -10.985 1.945 ;
        RECT -5.535 1.615 -4.985 1.945 ;
        RECT -13.450 1.425 -12.990 1.595 ;
        RECT -11.535 1.090 -11.365 1.615 ;
        RECT -5.155 1.090 -4.985 1.615 ;
        RECT -3.445 1.595 -3.155 2.320 ;
        RECT -1.615 1.945 -1.445 2.470 ;
        RECT 4.765 1.945 4.935 2.470 ;
        RECT -1.615 1.615 -1.065 1.945 ;
        RECT 4.385 1.615 4.935 1.945 ;
        RECT -3.530 1.425 -3.070 1.595 ;
        RECT -1.615 1.090 -1.445 1.615 ;
        RECT 4.765 1.090 4.935 1.615 ;
        RECT 6.475 1.595 6.765 2.320 ;
        RECT 8.305 1.945 8.475 2.470 ;
        RECT 14.685 1.945 14.855 2.470 ;
        RECT 8.305 1.615 8.855 1.945 ;
        RECT 14.305 1.615 14.855 1.945 ;
        RECT 6.390 1.425 6.850 1.595 ;
        RECT 8.305 1.090 8.475 1.615 ;
        RECT 14.685 1.090 14.855 1.615 ;
        RECT 16.395 1.595 16.685 2.320 ;
        RECT 18.225 1.945 18.395 2.470 ;
        RECT 18.225 1.615 18.775 1.945 ;
        RECT 16.310 1.425 16.770 1.595 ;
        RECT 18.225 1.090 18.395 1.615 ;
        RECT -286.115 -86.445 -285.945 -85.920 ;
        RECT -284.490 -86.335 -284.030 -86.165 ;
        RECT -286.495 -86.775 -285.945 -86.445 ;
        RECT -286.115 -87.300 -285.945 -86.775 ;
        RECT -284.405 -87.060 -284.115 -86.335 ;
        RECT -282.575 -86.445 -282.405 -85.920 ;
        RECT -276.195 -86.445 -276.025 -85.920 ;
        RECT -274.570 -86.335 -274.110 -86.165 ;
        RECT -282.575 -86.775 -282.025 -86.445 ;
        RECT -276.575 -86.775 -276.025 -86.445 ;
        RECT -282.575 -87.300 -282.405 -86.775 ;
        RECT -276.195 -87.300 -276.025 -86.775 ;
        RECT -274.485 -87.060 -274.195 -86.335 ;
        RECT -272.655 -86.445 -272.485 -85.920 ;
        RECT -266.275 -86.445 -266.105 -85.920 ;
        RECT -264.650 -86.335 -264.190 -86.165 ;
        RECT -272.655 -86.775 -272.105 -86.445 ;
        RECT -266.655 -86.775 -266.105 -86.445 ;
        RECT -272.655 -87.300 -272.485 -86.775 ;
        RECT -266.275 -87.300 -266.105 -86.775 ;
        RECT -264.565 -87.060 -264.275 -86.335 ;
        RECT -262.735 -86.445 -262.565 -85.920 ;
        RECT -256.355 -86.445 -256.185 -85.920 ;
        RECT -254.730 -86.335 -254.270 -86.165 ;
        RECT -262.735 -86.775 -262.185 -86.445 ;
        RECT -256.735 -86.775 -256.185 -86.445 ;
        RECT -262.735 -87.300 -262.565 -86.775 ;
        RECT -256.355 -87.300 -256.185 -86.775 ;
        RECT -254.645 -87.060 -254.355 -86.335 ;
        RECT -252.815 -86.445 -252.645 -85.920 ;
        RECT -246.435 -86.445 -246.265 -85.920 ;
        RECT -244.810 -86.335 -244.350 -86.165 ;
        RECT -252.815 -86.775 -252.265 -86.445 ;
        RECT -246.815 -86.775 -246.265 -86.445 ;
        RECT -252.815 -87.300 -252.645 -86.775 ;
        RECT -246.435 -87.300 -246.265 -86.775 ;
        RECT -244.725 -87.060 -244.435 -86.335 ;
        RECT -242.895 -86.445 -242.725 -85.920 ;
        RECT -236.515 -86.445 -236.345 -85.920 ;
        RECT -234.890 -86.335 -234.430 -86.165 ;
        RECT -242.895 -86.775 -242.345 -86.445 ;
        RECT -236.895 -86.775 -236.345 -86.445 ;
        RECT -242.895 -87.300 -242.725 -86.775 ;
        RECT -236.515 -87.300 -236.345 -86.775 ;
        RECT -234.805 -87.060 -234.515 -86.335 ;
        RECT -232.975 -86.445 -232.805 -85.920 ;
        RECT -226.595 -86.445 -226.425 -85.920 ;
        RECT -224.970 -86.335 -224.510 -86.165 ;
        RECT -232.975 -86.775 -232.425 -86.445 ;
        RECT -226.975 -86.775 -226.425 -86.445 ;
        RECT -232.975 -87.300 -232.805 -86.775 ;
        RECT -226.595 -87.300 -226.425 -86.775 ;
        RECT -224.885 -87.060 -224.595 -86.335 ;
        RECT -223.055 -86.445 -222.885 -85.920 ;
        RECT -216.675 -86.445 -216.505 -85.920 ;
        RECT -215.050 -86.335 -214.590 -86.165 ;
        RECT -223.055 -86.775 -222.505 -86.445 ;
        RECT -217.055 -86.775 -216.505 -86.445 ;
        RECT -223.055 -87.300 -222.885 -86.775 ;
        RECT -216.675 -87.300 -216.505 -86.775 ;
        RECT -214.965 -87.060 -214.675 -86.335 ;
        RECT -213.135 -86.445 -212.965 -85.920 ;
        RECT -206.755 -86.445 -206.585 -85.920 ;
        RECT -205.130 -86.335 -204.670 -86.165 ;
        RECT -213.135 -86.775 -212.585 -86.445 ;
        RECT -207.135 -86.775 -206.585 -86.445 ;
        RECT -213.135 -87.300 -212.965 -86.775 ;
        RECT -206.755 -87.300 -206.585 -86.775 ;
        RECT -205.045 -87.060 -204.755 -86.335 ;
        RECT -203.215 -86.445 -203.045 -85.920 ;
        RECT -196.835 -86.445 -196.665 -85.920 ;
        RECT -195.210 -86.335 -194.750 -86.165 ;
        RECT -203.215 -86.775 -202.665 -86.445 ;
        RECT -197.215 -86.775 -196.665 -86.445 ;
        RECT -203.215 -87.300 -203.045 -86.775 ;
        RECT -196.835 -87.300 -196.665 -86.775 ;
        RECT -195.125 -87.060 -194.835 -86.335 ;
        RECT -193.295 -86.445 -193.125 -85.920 ;
        RECT -186.915 -86.445 -186.745 -85.920 ;
        RECT -185.290 -86.335 -184.830 -86.165 ;
        RECT -193.295 -86.775 -192.745 -86.445 ;
        RECT -187.295 -86.775 -186.745 -86.445 ;
        RECT -193.295 -87.300 -193.125 -86.775 ;
        RECT -186.915 -87.300 -186.745 -86.775 ;
        RECT -185.205 -87.060 -184.915 -86.335 ;
        RECT -183.375 -86.445 -183.205 -85.920 ;
        RECT -176.995 -86.445 -176.825 -85.920 ;
        RECT -175.370 -86.335 -174.910 -86.165 ;
        RECT -183.375 -86.775 -182.825 -86.445 ;
        RECT -177.375 -86.775 -176.825 -86.445 ;
        RECT -183.375 -87.300 -183.205 -86.775 ;
        RECT -176.995 -87.300 -176.825 -86.775 ;
        RECT -175.285 -87.060 -174.995 -86.335 ;
        RECT -173.455 -86.445 -173.285 -85.920 ;
        RECT -167.075 -86.445 -166.905 -85.920 ;
        RECT -165.450 -86.335 -164.990 -86.165 ;
        RECT -173.455 -86.775 -172.905 -86.445 ;
        RECT -167.455 -86.775 -166.905 -86.445 ;
        RECT -173.455 -87.300 -173.285 -86.775 ;
        RECT -167.075 -87.300 -166.905 -86.775 ;
        RECT -165.365 -87.060 -165.075 -86.335 ;
        RECT -163.535 -86.445 -163.365 -85.920 ;
        RECT -157.155 -86.445 -156.985 -85.920 ;
        RECT -155.530 -86.335 -155.070 -86.165 ;
        RECT -163.535 -86.775 -162.985 -86.445 ;
        RECT -157.535 -86.775 -156.985 -86.445 ;
        RECT -163.535 -87.300 -163.365 -86.775 ;
        RECT -157.155 -87.300 -156.985 -86.775 ;
        RECT -155.445 -87.060 -155.155 -86.335 ;
        RECT -153.615 -86.445 -153.445 -85.920 ;
        RECT -147.235 -86.445 -147.065 -85.920 ;
        RECT -145.610 -86.335 -145.150 -86.165 ;
        RECT -153.615 -86.775 -153.065 -86.445 ;
        RECT -147.615 -86.775 -147.065 -86.445 ;
        RECT -153.615 -87.300 -153.445 -86.775 ;
        RECT -147.235 -87.300 -147.065 -86.775 ;
        RECT -145.525 -87.060 -145.235 -86.335 ;
        RECT -143.695 -86.445 -143.525 -85.920 ;
        RECT -137.315 -86.445 -137.145 -85.920 ;
        RECT -135.690 -86.335 -135.230 -86.165 ;
        RECT -143.695 -86.775 -143.145 -86.445 ;
        RECT -137.695 -86.775 -137.145 -86.445 ;
        RECT -143.695 -87.300 -143.525 -86.775 ;
        RECT -137.315 -87.300 -137.145 -86.775 ;
        RECT -135.605 -87.060 -135.315 -86.335 ;
        RECT -133.775 -86.445 -133.605 -85.920 ;
        RECT -127.395 -86.445 -127.225 -85.920 ;
        RECT -125.770 -86.335 -125.310 -86.165 ;
        RECT -133.775 -86.775 -133.225 -86.445 ;
        RECT -127.775 -86.775 -127.225 -86.445 ;
        RECT -133.775 -87.300 -133.605 -86.775 ;
        RECT -127.395 -87.300 -127.225 -86.775 ;
        RECT -125.685 -87.060 -125.395 -86.335 ;
        RECT -123.855 -86.445 -123.685 -85.920 ;
        RECT -117.475 -86.445 -117.305 -85.920 ;
        RECT -115.850 -86.335 -115.390 -86.165 ;
        RECT -123.855 -86.775 -123.305 -86.445 ;
        RECT -117.855 -86.775 -117.305 -86.445 ;
        RECT -123.855 -87.300 -123.685 -86.775 ;
        RECT -117.475 -87.300 -117.305 -86.775 ;
        RECT -115.765 -87.060 -115.475 -86.335 ;
        RECT -113.935 -86.445 -113.765 -85.920 ;
        RECT -107.555 -86.445 -107.385 -85.920 ;
        RECT -105.930 -86.335 -105.470 -86.165 ;
        RECT -113.935 -86.775 -113.385 -86.445 ;
        RECT -107.935 -86.775 -107.385 -86.445 ;
        RECT -113.935 -87.300 -113.765 -86.775 ;
        RECT -107.555 -87.300 -107.385 -86.775 ;
        RECT -105.845 -87.060 -105.555 -86.335 ;
        RECT -104.015 -86.445 -103.845 -85.920 ;
        RECT -97.635 -86.445 -97.465 -85.920 ;
        RECT -96.010 -86.335 -95.550 -86.165 ;
        RECT -104.015 -86.775 -103.465 -86.445 ;
        RECT -98.015 -86.775 -97.465 -86.445 ;
        RECT -104.015 -87.300 -103.845 -86.775 ;
        RECT -97.635 -87.300 -97.465 -86.775 ;
        RECT -95.925 -87.060 -95.635 -86.335 ;
        RECT -94.095 -86.445 -93.925 -85.920 ;
        RECT -87.715 -86.445 -87.545 -85.920 ;
        RECT -86.090 -86.335 -85.630 -86.165 ;
        RECT -94.095 -86.775 -93.545 -86.445 ;
        RECT -88.095 -86.775 -87.545 -86.445 ;
        RECT -94.095 -87.300 -93.925 -86.775 ;
        RECT -87.715 -87.300 -87.545 -86.775 ;
        RECT -86.005 -87.060 -85.715 -86.335 ;
        RECT -84.175 -86.445 -84.005 -85.920 ;
        RECT -77.795 -86.445 -77.625 -85.920 ;
        RECT -76.170 -86.335 -75.710 -86.165 ;
        RECT -84.175 -86.775 -83.625 -86.445 ;
        RECT -78.175 -86.775 -77.625 -86.445 ;
        RECT -84.175 -87.300 -84.005 -86.775 ;
        RECT -77.795 -87.300 -77.625 -86.775 ;
        RECT -76.085 -87.060 -75.795 -86.335 ;
        RECT -74.255 -86.445 -74.085 -85.920 ;
        RECT -67.875 -86.445 -67.705 -85.920 ;
        RECT -66.250 -86.335 -65.790 -86.165 ;
        RECT -74.255 -86.775 -73.705 -86.445 ;
        RECT -68.255 -86.775 -67.705 -86.445 ;
        RECT -74.255 -87.300 -74.085 -86.775 ;
        RECT -67.875 -87.300 -67.705 -86.775 ;
        RECT -66.165 -87.060 -65.875 -86.335 ;
        RECT -64.335 -86.445 -64.165 -85.920 ;
        RECT -57.955 -86.445 -57.785 -85.920 ;
        RECT -56.330 -86.335 -55.870 -86.165 ;
        RECT -64.335 -86.775 -63.785 -86.445 ;
        RECT -58.335 -86.775 -57.785 -86.445 ;
        RECT -64.335 -87.300 -64.165 -86.775 ;
        RECT -57.955 -87.300 -57.785 -86.775 ;
        RECT -56.245 -87.060 -55.955 -86.335 ;
        RECT -54.415 -86.445 -54.245 -85.920 ;
        RECT -48.035 -86.445 -47.865 -85.920 ;
        RECT -46.410 -86.335 -45.950 -86.165 ;
        RECT -54.415 -86.775 -53.865 -86.445 ;
        RECT -48.415 -86.775 -47.865 -86.445 ;
        RECT -54.415 -87.300 -54.245 -86.775 ;
        RECT -48.035 -87.300 -47.865 -86.775 ;
        RECT -46.325 -87.060 -46.035 -86.335 ;
        RECT -44.495 -86.445 -44.325 -85.920 ;
        RECT -38.115 -86.445 -37.945 -85.920 ;
        RECT -36.490 -86.335 -36.030 -86.165 ;
        RECT -44.495 -86.775 -43.945 -86.445 ;
        RECT -38.495 -86.775 -37.945 -86.445 ;
        RECT -44.495 -87.300 -44.325 -86.775 ;
        RECT -38.115 -87.300 -37.945 -86.775 ;
        RECT -36.405 -87.060 -36.115 -86.335 ;
        RECT -34.575 -86.445 -34.405 -85.920 ;
        RECT -28.195 -86.445 -28.025 -85.920 ;
        RECT -26.570 -86.335 -26.110 -86.165 ;
        RECT -34.575 -86.775 -34.025 -86.445 ;
        RECT -28.575 -86.775 -28.025 -86.445 ;
        RECT -34.575 -87.300 -34.405 -86.775 ;
        RECT -28.195 -87.300 -28.025 -86.775 ;
        RECT -26.485 -87.060 -26.195 -86.335 ;
        RECT -24.655 -86.445 -24.485 -85.920 ;
        RECT -18.275 -86.445 -18.105 -85.920 ;
        RECT -16.650 -86.335 -16.190 -86.165 ;
        RECT -24.655 -86.775 -24.105 -86.445 ;
        RECT -18.655 -86.775 -18.105 -86.445 ;
        RECT -24.655 -87.300 -24.485 -86.775 ;
        RECT -18.275 -87.300 -18.105 -86.775 ;
        RECT -16.565 -87.060 -16.275 -86.335 ;
        RECT -14.735 -86.445 -14.565 -85.920 ;
        RECT -8.355 -86.445 -8.185 -85.920 ;
        RECT -6.730 -86.335 -6.270 -86.165 ;
        RECT -14.735 -86.775 -14.185 -86.445 ;
        RECT -8.735 -86.775 -8.185 -86.445 ;
        RECT -14.735 -87.300 -14.565 -86.775 ;
        RECT -8.355 -87.300 -8.185 -86.775 ;
        RECT -6.645 -87.060 -6.355 -86.335 ;
        RECT -4.815 -86.445 -4.645 -85.920 ;
        RECT 1.565 -86.445 1.735 -85.920 ;
        RECT 3.190 -86.335 3.650 -86.165 ;
        RECT -4.815 -86.775 -4.265 -86.445 ;
        RECT 1.185 -86.775 1.735 -86.445 ;
        RECT -4.815 -87.300 -4.645 -86.775 ;
        RECT 1.565 -87.300 1.735 -86.775 ;
        RECT 3.275 -87.060 3.565 -86.335 ;
        RECT 5.105 -86.445 5.275 -85.920 ;
        RECT 11.485 -86.445 11.655 -85.920 ;
        RECT 13.110 -86.335 13.570 -86.165 ;
        RECT 5.105 -86.775 5.655 -86.445 ;
        RECT 11.105 -86.775 11.655 -86.445 ;
        RECT 5.105 -87.300 5.275 -86.775 ;
        RECT 11.485 -87.300 11.655 -86.775 ;
        RECT 13.195 -87.060 13.485 -86.335 ;
        RECT 15.025 -86.445 15.195 -85.920 ;
        RECT 21.405 -86.445 21.575 -85.920 ;
        RECT 23.030 -86.335 23.490 -86.165 ;
        RECT 15.025 -86.775 15.575 -86.445 ;
        RECT 21.025 -86.775 21.575 -86.445 ;
        RECT 15.025 -87.300 15.195 -86.775 ;
        RECT 21.405 -87.300 21.575 -86.775 ;
        RECT 23.115 -87.060 23.405 -86.335 ;
        RECT 24.945 -86.445 25.115 -85.920 ;
        RECT 24.945 -86.775 25.495 -86.445 ;
        RECT 24.945 -87.300 25.115 -86.775 ;
        RECT -280.910 -87.815 -277.690 -87.645 ;
        RECT -270.990 -87.815 -267.770 -87.645 ;
        RECT -261.070 -87.815 -257.850 -87.645 ;
        RECT -251.150 -87.815 -247.930 -87.645 ;
        RECT -241.230 -87.815 -238.010 -87.645 ;
        RECT -231.310 -87.815 -228.090 -87.645 ;
        RECT -221.390 -87.815 -218.170 -87.645 ;
        RECT -211.470 -87.815 -208.250 -87.645 ;
        RECT -201.550 -87.815 -198.330 -87.645 ;
        RECT -191.630 -87.815 -188.410 -87.645 ;
        RECT -181.710 -87.815 -178.490 -87.645 ;
        RECT -171.790 -87.815 -168.570 -87.645 ;
        RECT -161.870 -87.815 -158.650 -87.645 ;
        RECT -151.950 -87.815 -148.730 -87.645 ;
        RECT -142.030 -87.815 -138.810 -87.645 ;
        RECT -132.110 -87.815 -128.890 -87.645 ;
        RECT -122.190 -87.815 -118.970 -87.645 ;
        RECT -112.270 -87.815 -109.050 -87.645 ;
        RECT -102.350 -87.815 -99.130 -87.645 ;
        RECT -92.430 -87.815 -89.210 -87.645 ;
        RECT -82.510 -87.815 -79.290 -87.645 ;
        RECT -72.590 -87.815 -69.370 -87.645 ;
        RECT -62.670 -87.815 -59.450 -87.645 ;
        RECT -52.750 -87.815 -49.530 -87.645 ;
        RECT -42.830 -87.815 -39.610 -87.645 ;
        RECT -32.910 -87.815 -29.690 -87.645 ;
        RECT -22.990 -87.815 -19.770 -87.645 ;
        RECT -13.070 -87.815 -9.850 -87.645 ;
        RECT -3.150 -87.815 0.070 -87.645 ;
        RECT 6.770 -87.815 9.990 -87.645 ;
        RECT 16.690 -87.815 19.910 -87.645 ;
        RECT -279.925 -88.615 -279.615 -87.815 ;
        RECT -279.445 -88.540 -279.155 -87.815 ;
        RECT -278.985 -88.615 -278.675 -87.815 ;
        RECT -270.005 -88.615 -269.695 -87.815 ;
        RECT -269.525 -88.540 -269.235 -87.815 ;
        RECT -269.065 -88.615 -268.755 -87.815 ;
        RECT -260.085 -88.615 -259.775 -87.815 ;
        RECT -259.605 -88.540 -259.315 -87.815 ;
        RECT -259.145 -88.615 -258.835 -87.815 ;
        RECT -250.165 -88.615 -249.855 -87.815 ;
        RECT -249.685 -88.540 -249.395 -87.815 ;
        RECT -249.225 -88.615 -248.915 -87.815 ;
        RECT -240.245 -88.615 -239.935 -87.815 ;
        RECT -239.765 -88.540 -239.475 -87.815 ;
        RECT -239.305 -88.615 -238.995 -87.815 ;
        RECT -230.325 -88.615 -230.015 -87.815 ;
        RECT -229.845 -88.540 -229.555 -87.815 ;
        RECT -229.385 -88.615 -229.075 -87.815 ;
        RECT -220.405 -88.615 -220.095 -87.815 ;
        RECT -219.925 -88.540 -219.635 -87.815 ;
        RECT -219.465 -88.615 -219.155 -87.815 ;
        RECT -210.485 -88.615 -210.175 -87.815 ;
        RECT -210.005 -88.540 -209.715 -87.815 ;
        RECT -209.545 -88.615 -209.235 -87.815 ;
        RECT -200.565 -88.615 -200.255 -87.815 ;
        RECT -200.085 -88.540 -199.795 -87.815 ;
        RECT -199.625 -88.615 -199.315 -87.815 ;
        RECT -190.645 -88.615 -190.335 -87.815 ;
        RECT -190.165 -88.540 -189.875 -87.815 ;
        RECT -189.705 -88.615 -189.395 -87.815 ;
        RECT -180.725 -88.615 -180.415 -87.815 ;
        RECT -180.245 -88.540 -179.955 -87.815 ;
        RECT -179.785 -88.615 -179.475 -87.815 ;
        RECT -170.805 -88.615 -170.495 -87.815 ;
        RECT -170.325 -88.540 -170.035 -87.815 ;
        RECT -169.865 -88.615 -169.555 -87.815 ;
        RECT -160.885 -88.615 -160.575 -87.815 ;
        RECT -160.405 -88.540 -160.115 -87.815 ;
        RECT -159.945 -88.615 -159.635 -87.815 ;
        RECT -150.965 -88.615 -150.655 -87.815 ;
        RECT -150.485 -88.540 -150.195 -87.815 ;
        RECT -150.025 -88.615 -149.715 -87.815 ;
        RECT -141.045 -88.615 -140.735 -87.815 ;
        RECT -140.565 -88.540 -140.275 -87.815 ;
        RECT -140.105 -88.615 -139.795 -87.815 ;
        RECT -131.125 -88.615 -130.815 -87.815 ;
        RECT -130.645 -88.540 -130.355 -87.815 ;
        RECT -130.185 -88.615 -129.875 -87.815 ;
        RECT -121.205 -88.615 -120.895 -87.815 ;
        RECT -120.725 -88.540 -120.435 -87.815 ;
        RECT -120.265 -88.615 -119.955 -87.815 ;
        RECT -111.285 -88.615 -110.975 -87.815 ;
        RECT -110.805 -88.540 -110.515 -87.815 ;
        RECT -110.345 -88.615 -110.035 -87.815 ;
        RECT -101.365 -88.615 -101.055 -87.815 ;
        RECT -100.885 -88.540 -100.595 -87.815 ;
        RECT -100.425 -88.615 -100.115 -87.815 ;
        RECT -91.445 -88.615 -91.135 -87.815 ;
        RECT -90.965 -88.540 -90.675 -87.815 ;
        RECT -90.505 -88.615 -90.195 -87.815 ;
        RECT -81.525 -88.615 -81.215 -87.815 ;
        RECT -81.045 -88.540 -80.755 -87.815 ;
        RECT -80.585 -88.615 -80.275 -87.815 ;
        RECT -71.605 -88.615 -71.295 -87.815 ;
        RECT -71.125 -88.540 -70.835 -87.815 ;
        RECT -70.665 -88.615 -70.355 -87.815 ;
        RECT -61.685 -88.615 -61.375 -87.815 ;
        RECT -61.205 -88.540 -60.915 -87.815 ;
        RECT -60.745 -88.615 -60.435 -87.815 ;
        RECT -51.765 -88.615 -51.455 -87.815 ;
        RECT -51.285 -88.540 -50.995 -87.815 ;
        RECT -50.825 -88.615 -50.515 -87.815 ;
        RECT -41.845 -88.615 -41.535 -87.815 ;
        RECT -41.365 -88.540 -41.075 -87.815 ;
        RECT -40.905 -88.615 -40.595 -87.815 ;
        RECT -31.925 -88.615 -31.615 -87.815 ;
        RECT -31.445 -88.540 -31.155 -87.815 ;
        RECT -30.985 -88.615 -30.675 -87.815 ;
        RECT -22.005 -88.615 -21.695 -87.815 ;
        RECT -21.525 -88.540 -21.235 -87.815 ;
        RECT -21.065 -88.615 -20.755 -87.815 ;
        RECT -12.085 -88.615 -11.775 -87.815 ;
        RECT -11.605 -88.540 -11.315 -87.815 ;
        RECT -11.145 -88.615 -10.835 -87.815 ;
        RECT -2.165 -88.615 -1.855 -87.815 ;
        RECT -1.685 -88.540 -1.395 -87.815 ;
        RECT -1.225 -88.615 -0.915 -87.815 ;
        RECT 7.755 -88.615 8.065 -87.815 ;
        RECT 8.235 -88.540 8.525 -87.815 ;
        RECT 8.695 -88.615 9.005 -87.815 ;
        RECT 17.675 -88.615 17.985 -87.815 ;
        RECT 18.155 -88.540 18.445 -87.815 ;
        RECT 18.615 -88.615 18.925 -87.815 ;
        RECT -284.885 -90.365 -284.575 -89.565 ;
        RECT -284.405 -90.365 -284.115 -89.640 ;
        RECT -283.945 -90.365 -283.635 -89.565 ;
        RECT -274.965 -90.365 -274.655 -89.565 ;
        RECT -274.485 -90.365 -274.195 -89.640 ;
        RECT -274.025 -90.365 -273.715 -89.565 ;
        RECT -265.045 -90.365 -264.735 -89.565 ;
        RECT -264.565 -90.365 -264.275 -89.640 ;
        RECT -264.105 -90.365 -263.795 -89.565 ;
        RECT -255.125 -90.365 -254.815 -89.565 ;
        RECT -254.645 -90.365 -254.355 -89.640 ;
        RECT -254.185 -90.365 -253.875 -89.565 ;
        RECT -245.205 -90.365 -244.895 -89.565 ;
        RECT -244.725 -90.365 -244.435 -89.640 ;
        RECT -244.265 -90.365 -243.955 -89.565 ;
        RECT -235.285 -90.365 -234.975 -89.565 ;
        RECT -234.805 -90.365 -234.515 -89.640 ;
        RECT -234.345 -90.365 -234.035 -89.565 ;
        RECT -225.365 -90.365 -225.055 -89.565 ;
        RECT -224.885 -90.365 -224.595 -89.640 ;
        RECT -224.425 -90.365 -224.115 -89.565 ;
        RECT -215.445 -90.365 -215.135 -89.565 ;
        RECT -214.965 -90.365 -214.675 -89.640 ;
        RECT -214.505 -90.365 -214.195 -89.565 ;
        RECT -205.525 -90.365 -205.215 -89.565 ;
        RECT -205.045 -90.365 -204.755 -89.640 ;
        RECT -204.585 -90.365 -204.275 -89.565 ;
        RECT -195.605 -90.365 -195.295 -89.565 ;
        RECT -195.125 -90.365 -194.835 -89.640 ;
        RECT -194.665 -90.365 -194.355 -89.565 ;
        RECT -185.685 -90.365 -185.375 -89.565 ;
        RECT -185.205 -90.365 -184.915 -89.640 ;
        RECT -184.745 -90.365 -184.435 -89.565 ;
        RECT -175.765 -90.365 -175.455 -89.565 ;
        RECT -175.285 -90.365 -174.995 -89.640 ;
        RECT -174.825 -90.365 -174.515 -89.565 ;
        RECT -165.845 -90.365 -165.535 -89.565 ;
        RECT -165.365 -90.365 -165.075 -89.640 ;
        RECT -164.905 -90.365 -164.595 -89.565 ;
        RECT -155.925 -90.365 -155.615 -89.565 ;
        RECT -155.445 -90.365 -155.155 -89.640 ;
        RECT -154.985 -90.365 -154.675 -89.565 ;
        RECT -146.005 -90.365 -145.695 -89.565 ;
        RECT -145.525 -90.365 -145.235 -89.640 ;
        RECT -145.065 -90.365 -144.755 -89.565 ;
        RECT -136.085 -90.365 -135.775 -89.565 ;
        RECT -135.605 -90.365 -135.315 -89.640 ;
        RECT -135.145 -90.365 -134.835 -89.565 ;
        RECT -126.165 -90.365 -125.855 -89.565 ;
        RECT -125.685 -90.365 -125.395 -89.640 ;
        RECT -125.225 -90.365 -124.915 -89.565 ;
        RECT -116.245 -90.365 -115.935 -89.565 ;
        RECT -115.765 -90.365 -115.475 -89.640 ;
        RECT -115.305 -90.365 -114.995 -89.565 ;
        RECT -106.325 -90.365 -106.015 -89.565 ;
        RECT -105.845 -90.365 -105.555 -89.640 ;
        RECT -105.385 -90.365 -105.075 -89.565 ;
        RECT -96.405 -90.365 -96.095 -89.565 ;
        RECT -95.925 -90.365 -95.635 -89.640 ;
        RECT -95.465 -90.365 -95.155 -89.565 ;
        RECT -86.485 -90.365 -86.175 -89.565 ;
        RECT -86.005 -90.365 -85.715 -89.640 ;
        RECT -85.545 -90.365 -85.235 -89.565 ;
        RECT -76.565 -90.365 -76.255 -89.565 ;
        RECT -76.085 -90.365 -75.795 -89.640 ;
        RECT -75.625 -90.365 -75.315 -89.565 ;
        RECT -66.645 -90.365 -66.335 -89.565 ;
        RECT -66.165 -90.365 -65.875 -89.640 ;
        RECT -65.705 -90.365 -65.395 -89.565 ;
        RECT -56.725 -90.365 -56.415 -89.565 ;
        RECT -56.245 -90.365 -55.955 -89.640 ;
        RECT -55.785 -90.365 -55.475 -89.565 ;
        RECT -46.805 -90.365 -46.495 -89.565 ;
        RECT -46.325 -90.365 -46.035 -89.640 ;
        RECT -45.865 -90.365 -45.555 -89.565 ;
        RECT -36.885 -90.365 -36.575 -89.565 ;
        RECT -36.405 -90.365 -36.115 -89.640 ;
        RECT -35.945 -90.365 -35.635 -89.565 ;
        RECT -26.965 -90.365 -26.655 -89.565 ;
        RECT -26.485 -90.365 -26.195 -89.640 ;
        RECT -26.025 -90.365 -25.715 -89.565 ;
        RECT -17.045 -90.365 -16.735 -89.565 ;
        RECT -16.565 -90.365 -16.275 -89.640 ;
        RECT -16.105 -90.365 -15.795 -89.565 ;
        RECT -7.125 -90.365 -6.815 -89.565 ;
        RECT -6.645 -90.365 -6.355 -89.640 ;
        RECT -6.185 -90.365 -5.875 -89.565 ;
        RECT 2.795 -90.365 3.105 -89.565 ;
        RECT 3.275 -90.365 3.565 -89.640 ;
        RECT 3.735 -90.365 4.045 -89.565 ;
        RECT 12.715 -90.365 13.025 -89.565 ;
        RECT 13.195 -90.365 13.485 -89.640 ;
        RECT 13.655 -90.365 13.965 -89.565 ;
        RECT 22.635 -90.365 22.945 -89.565 ;
        RECT 23.115 -90.365 23.405 -89.640 ;
        RECT 23.575 -90.365 23.885 -89.565 ;
        RECT -285.870 -90.535 -282.650 -90.365 ;
        RECT -275.950 -90.535 -272.730 -90.365 ;
        RECT -266.030 -90.535 -262.810 -90.365 ;
        RECT -256.110 -90.535 -252.890 -90.365 ;
        RECT -246.190 -90.535 -242.970 -90.365 ;
        RECT -236.270 -90.535 -233.050 -90.365 ;
        RECT -226.350 -90.535 -223.130 -90.365 ;
        RECT -216.430 -90.535 -213.210 -90.365 ;
        RECT -206.510 -90.535 -203.290 -90.365 ;
        RECT -196.590 -90.535 -193.370 -90.365 ;
        RECT -186.670 -90.535 -183.450 -90.365 ;
        RECT -176.750 -90.535 -173.530 -90.365 ;
        RECT -166.830 -90.535 -163.610 -90.365 ;
        RECT -156.910 -90.535 -153.690 -90.365 ;
        RECT -146.990 -90.535 -143.770 -90.365 ;
        RECT -137.070 -90.535 -133.850 -90.365 ;
        RECT -127.150 -90.535 -123.930 -90.365 ;
        RECT -117.230 -90.535 -114.010 -90.365 ;
        RECT -107.310 -90.535 -104.090 -90.365 ;
        RECT -97.390 -90.535 -94.170 -90.365 ;
        RECT -87.470 -90.535 -84.250 -90.365 ;
        RECT -77.550 -90.535 -74.330 -90.365 ;
        RECT -67.630 -90.535 -64.410 -90.365 ;
        RECT -57.710 -90.535 -54.490 -90.365 ;
        RECT -47.790 -90.535 -44.570 -90.365 ;
        RECT -37.870 -90.535 -34.650 -90.365 ;
        RECT -27.950 -90.535 -24.730 -90.365 ;
        RECT -18.030 -90.535 -14.810 -90.365 ;
        RECT -8.110 -90.535 -4.890 -90.365 ;
        RECT 1.810 -90.535 5.030 -90.365 ;
        RECT 11.730 -90.535 14.950 -90.365 ;
        RECT 21.650 -90.535 24.870 -90.365 ;
        RECT -281.155 -91.405 -280.985 -90.880 ;
        RECT -281.535 -91.735 -280.985 -91.405 ;
        RECT -281.155 -92.260 -280.985 -91.735 ;
        RECT -279.445 -91.755 -279.155 -91.030 ;
        RECT -277.615 -91.405 -277.445 -90.880 ;
        RECT -271.235 -91.405 -271.065 -90.880 ;
        RECT -277.615 -91.735 -277.065 -91.405 ;
        RECT -271.615 -91.735 -271.065 -91.405 ;
        RECT -279.530 -91.925 -279.070 -91.755 ;
        RECT -277.615 -92.260 -277.445 -91.735 ;
        RECT -271.235 -92.260 -271.065 -91.735 ;
        RECT -269.525 -91.755 -269.235 -91.030 ;
        RECT -267.695 -91.405 -267.525 -90.880 ;
        RECT -261.315 -91.405 -261.145 -90.880 ;
        RECT -267.695 -91.735 -267.145 -91.405 ;
        RECT -261.695 -91.735 -261.145 -91.405 ;
        RECT -269.610 -91.925 -269.150 -91.755 ;
        RECT -267.695 -92.260 -267.525 -91.735 ;
        RECT -261.315 -92.260 -261.145 -91.735 ;
        RECT -259.605 -91.755 -259.315 -91.030 ;
        RECT -257.775 -91.405 -257.605 -90.880 ;
        RECT -251.395 -91.405 -251.225 -90.880 ;
        RECT -257.775 -91.735 -257.225 -91.405 ;
        RECT -251.775 -91.735 -251.225 -91.405 ;
        RECT -259.690 -91.925 -259.230 -91.755 ;
        RECT -257.775 -92.260 -257.605 -91.735 ;
        RECT -251.395 -92.260 -251.225 -91.735 ;
        RECT -249.685 -91.755 -249.395 -91.030 ;
        RECT -247.855 -91.405 -247.685 -90.880 ;
        RECT -241.475 -91.405 -241.305 -90.880 ;
        RECT -247.855 -91.735 -247.305 -91.405 ;
        RECT -241.855 -91.735 -241.305 -91.405 ;
        RECT -249.770 -91.925 -249.310 -91.755 ;
        RECT -247.855 -92.260 -247.685 -91.735 ;
        RECT -241.475 -92.260 -241.305 -91.735 ;
        RECT -239.765 -91.755 -239.475 -91.030 ;
        RECT -237.935 -91.405 -237.765 -90.880 ;
        RECT -231.555 -91.405 -231.385 -90.880 ;
        RECT -237.935 -91.735 -237.385 -91.405 ;
        RECT -231.935 -91.735 -231.385 -91.405 ;
        RECT -239.850 -91.925 -239.390 -91.755 ;
        RECT -237.935 -92.260 -237.765 -91.735 ;
        RECT -231.555 -92.260 -231.385 -91.735 ;
        RECT -229.845 -91.755 -229.555 -91.030 ;
        RECT -228.015 -91.405 -227.845 -90.880 ;
        RECT -221.635 -91.405 -221.465 -90.880 ;
        RECT -228.015 -91.735 -227.465 -91.405 ;
        RECT -222.015 -91.735 -221.465 -91.405 ;
        RECT -229.930 -91.925 -229.470 -91.755 ;
        RECT -228.015 -92.260 -227.845 -91.735 ;
        RECT -221.635 -92.260 -221.465 -91.735 ;
        RECT -219.925 -91.755 -219.635 -91.030 ;
        RECT -218.095 -91.405 -217.925 -90.880 ;
        RECT -211.715 -91.405 -211.545 -90.880 ;
        RECT -218.095 -91.735 -217.545 -91.405 ;
        RECT -212.095 -91.735 -211.545 -91.405 ;
        RECT -220.010 -91.925 -219.550 -91.755 ;
        RECT -218.095 -92.260 -217.925 -91.735 ;
        RECT -211.715 -92.260 -211.545 -91.735 ;
        RECT -210.005 -91.755 -209.715 -91.030 ;
        RECT -208.175 -91.405 -208.005 -90.880 ;
        RECT -201.795 -91.405 -201.625 -90.880 ;
        RECT -208.175 -91.735 -207.625 -91.405 ;
        RECT -202.175 -91.735 -201.625 -91.405 ;
        RECT -210.090 -91.925 -209.630 -91.755 ;
        RECT -208.175 -92.260 -208.005 -91.735 ;
        RECT -201.795 -92.260 -201.625 -91.735 ;
        RECT -200.085 -91.755 -199.795 -91.030 ;
        RECT -198.255 -91.405 -198.085 -90.880 ;
        RECT -191.875 -91.405 -191.705 -90.880 ;
        RECT -198.255 -91.735 -197.705 -91.405 ;
        RECT -192.255 -91.735 -191.705 -91.405 ;
        RECT -200.170 -91.925 -199.710 -91.755 ;
        RECT -198.255 -92.260 -198.085 -91.735 ;
        RECT -191.875 -92.260 -191.705 -91.735 ;
        RECT -190.165 -91.755 -189.875 -91.030 ;
        RECT -188.335 -91.405 -188.165 -90.880 ;
        RECT -181.955 -91.405 -181.785 -90.880 ;
        RECT -188.335 -91.735 -187.785 -91.405 ;
        RECT -182.335 -91.735 -181.785 -91.405 ;
        RECT -190.250 -91.925 -189.790 -91.755 ;
        RECT -188.335 -92.260 -188.165 -91.735 ;
        RECT -181.955 -92.260 -181.785 -91.735 ;
        RECT -180.245 -91.755 -179.955 -91.030 ;
        RECT -178.415 -91.405 -178.245 -90.880 ;
        RECT -172.035 -91.405 -171.865 -90.880 ;
        RECT -178.415 -91.735 -177.865 -91.405 ;
        RECT -172.415 -91.735 -171.865 -91.405 ;
        RECT -180.330 -91.925 -179.870 -91.755 ;
        RECT -178.415 -92.260 -178.245 -91.735 ;
        RECT -172.035 -92.260 -171.865 -91.735 ;
        RECT -170.325 -91.755 -170.035 -91.030 ;
        RECT -168.495 -91.405 -168.325 -90.880 ;
        RECT -162.115 -91.405 -161.945 -90.880 ;
        RECT -168.495 -91.735 -167.945 -91.405 ;
        RECT -162.495 -91.735 -161.945 -91.405 ;
        RECT -170.410 -91.925 -169.950 -91.755 ;
        RECT -168.495 -92.260 -168.325 -91.735 ;
        RECT -162.115 -92.260 -161.945 -91.735 ;
        RECT -160.405 -91.755 -160.115 -91.030 ;
        RECT -158.575 -91.405 -158.405 -90.880 ;
        RECT -152.195 -91.405 -152.025 -90.880 ;
        RECT -158.575 -91.735 -158.025 -91.405 ;
        RECT -152.575 -91.735 -152.025 -91.405 ;
        RECT -160.490 -91.925 -160.030 -91.755 ;
        RECT -158.575 -92.260 -158.405 -91.735 ;
        RECT -152.195 -92.260 -152.025 -91.735 ;
        RECT -150.485 -91.755 -150.195 -91.030 ;
        RECT -148.655 -91.405 -148.485 -90.880 ;
        RECT -142.275 -91.405 -142.105 -90.880 ;
        RECT -148.655 -91.735 -148.105 -91.405 ;
        RECT -142.655 -91.735 -142.105 -91.405 ;
        RECT -150.570 -91.925 -150.110 -91.755 ;
        RECT -148.655 -92.260 -148.485 -91.735 ;
        RECT -142.275 -92.260 -142.105 -91.735 ;
        RECT -140.565 -91.755 -140.275 -91.030 ;
        RECT -138.735 -91.405 -138.565 -90.880 ;
        RECT -132.355 -91.405 -132.185 -90.880 ;
        RECT -138.735 -91.735 -138.185 -91.405 ;
        RECT -132.735 -91.735 -132.185 -91.405 ;
        RECT -140.650 -91.925 -140.190 -91.755 ;
        RECT -138.735 -92.260 -138.565 -91.735 ;
        RECT -132.355 -92.260 -132.185 -91.735 ;
        RECT -130.645 -91.755 -130.355 -91.030 ;
        RECT -128.815 -91.405 -128.645 -90.880 ;
        RECT -122.435 -91.405 -122.265 -90.880 ;
        RECT -128.815 -91.735 -128.265 -91.405 ;
        RECT -122.815 -91.735 -122.265 -91.405 ;
        RECT -130.730 -91.925 -130.270 -91.755 ;
        RECT -128.815 -92.260 -128.645 -91.735 ;
        RECT -122.435 -92.260 -122.265 -91.735 ;
        RECT -120.725 -91.755 -120.435 -91.030 ;
        RECT -118.895 -91.405 -118.725 -90.880 ;
        RECT -112.515 -91.405 -112.345 -90.880 ;
        RECT -118.895 -91.735 -118.345 -91.405 ;
        RECT -112.895 -91.735 -112.345 -91.405 ;
        RECT -120.810 -91.925 -120.350 -91.755 ;
        RECT -118.895 -92.260 -118.725 -91.735 ;
        RECT -112.515 -92.260 -112.345 -91.735 ;
        RECT -110.805 -91.755 -110.515 -91.030 ;
        RECT -108.975 -91.405 -108.805 -90.880 ;
        RECT -102.595 -91.405 -102.425 -90.880 ;
        RECT -108.975 -91.735 -108.425 -91.405 ;
        RECT -102.975 -91.735 -102.425 -91.405 ;
        RECT -110.890 -91.925 -110.430 -91.755 ;
        RECT -108.975 -92.260 -108.805 -91.735 ;
        RECT -102.595 -92.260 -102.425 -91.735 ;
        RECT -100.885 -91.755 -100.595 -91.030 ;
        RECT -99.055 -91.405 -98.885 -90.880 ;
        RECT -92.675 -91.405 -92.505 -90.880 ;
        RECT -99.055 -91.735 -98.505 -91.405 ;
        RECT -93.055 -91.735 -92.505 -91.405 ;
        RECT -100.970 -91.925 -100.510 -91.755 ;
        RECT -99.055 -92.260 -98.885 -91.735 ;
        RECT -92.675 -92.260 -92.505 -91.735 ;
        RECT -90.965 -91.755 -90.675 -91.030 ;
        RECT -89.135 -91.405 -88.965 -90.880 ;
        RECT -82.755 -91.405 -82.585 -90.880 ;
        RECT -89.135 -91.735 -88.585 -91.405 ;
        RECT -83.135 -91.735 -82.585 -91.405 ;
        RECT -91.050 -91.925 -90.590 -91.755 ;
        RECT -89.135 -92.260 -88.965 -91.735 ;
        RECT -82.755 -92.260 -82.585 -91.735 ;
        RECT -81.045 -91.755 -80.755 -91.030 ;
        RECT -79.215 -91.405 -79.045 -90.880 ;
        RECT -72.835 -91.405 -72.665 -90.880 ;
        RECT -79.215 -91.735 -78.665 -91.405 ;
        RECT -73.215 -91.735 -72.665 -91.405 ;
        RECT -81.130 -91.925 -80.670 -91.755 ;
        RECT -79.215 -92.260 -79.045 -91.735 ;
        RECT -72.835 -92.260 -72.665 -91.735 ;
        RECT -71.125 -91.755 -70.835 -91.030 ;
        RECT -69.295 -91.405 -69.125 -90.880 ;
        RECT -62.915 -91.405 -62.745 -90.880 ;
        RECT -69.295 -91.735 -68.745 -91.405 ;
        RECT -63.295 -91.735 -62.745 -91.405 ;
        RECT -71.210 -91.925 -70.750 -91.755 ;
        RECT -69.295 -92.260 -69.125 -91.735 ;
        RECT -62.915 -92.260 -62.745 -91.735 ;
        RECT -61.205 -91.755 -60.915 -91.030 ;
        RECT -59.375 -91.405 -59.205 -90.880 ;
        RECT -52.995 -91.405 -52.825 -90.880 ;
        RECT -59.375 -91.735 -58.825 -91.405 ;
        RECT -53.375 -91.735 -52.825 -91.405 ;
        RECT -61.290 -91.925 -60.830 -91.755 ;
        RECT -59.375 -92.260 -59.205 -91.735 ;
        RECT -52.995 -92.260 -52.825 -91.735 ;
        RECT -51.285 -91.755 -50.995 -91.030 ;
        RECT -49.455 -91.405 -49.285 -90.880 ;
        RECT -43.075 -91.405 -42.905 -90.880 ;
        RECT -49.455 -91.735 -48.905 -91.405 ;
        RECT -43.455 -91.735 -42.905 -91.405 ;
        RECT -51.370 -91.925 -50.910 -91.755 ;
        RECT -49.455 -92.260 -49.285 -91.735 ;
        RECT -43.075 -92.260 -42.905 -91.735 ;
        RECT -41.365 -91.755 -41.075 -91.030 ;
        RECT -39.535 -91.405 -39.365 -90.880 ;
        RECT -33.155 -91.405 -32.985 -90.880 ;
        RECT -39.535 -91.735 -38.985 -91.405 ;
        RECT -33.535 -91.735 -32.985 -91.405 ;
        RECT -41.450 -91.925 -40.990 -91.755 ;
        RECT -39.535 -92.260 -39.365 -91.735 ;
        RECT -33.155 -92.260 -32.985 -91.735 ;
        RECT -31.445 -91.755 -31.155 -91.030 ;
        RECT -29.615 -91.405 -29.445 -90.880 ;
        RECT -23.235 -91.405 -23.065 -90.880 ;
        RECT -29.615 -91.735 -29.065 -91.405 ;
        RECT -23.615 -91.735 -23.065 -91.405 ;
        RECT -31.530 -91.925 -31.070 -91.755 ;
        RECT -29.615 -92.260 -29.445 -91.735 ;
        RECT -23.235 -92.260 -23.065 -91.735 ;
        RECT -21.525 -91.755 -21.235 -91.030 ;
        RECT -19.695 -91.405 -19.525 -90.880 ;
        RECT -13.315 -91.405 -13.145 -90.880 ;
        RECT -19.695 -91.735 -19.145 -91.405 ;
        RECT -13.695 -91.735 -13.145 -91.405 ;
        RECT -21.610 -91.925 -21.150 -91.755 ;
        RECT -19.695 -92.260 -19.525 -91.735 ;
        RECT -13.315 -92.260 -13.145 -91.735 ;
        RECT -11.605 -91.755 -11.315 -91.030 ;
        RECT -9.775 -91.405 -9.605 -90.880 ;
        RECT -3.395 -91.405 -3.225 -90.880 ;
        RECT -9.775 -91.735 -9.225 -91.405 ;
        RECT -3.775 -91.735 -3.225 -91.405 ;
        RECT -11.690 -91.925 -11.230 -91.755 ;
        RECT -9.775 -92.260 -9.605 -91.735 ;
        RECT -3.395 -92.260 -3.225 -91.735 ;
        RECT -1.685 -91.755 -1.395 -91.030 ;
        RECT 0.145 -91.405 0.315 -90.880 ;
        RECT 6.525 -91.405 6.695 -90.880 ;
        RECT 0.145 -91.735 0.695 -91.405 ;
        RECT 6.145 -91.735 6.695 -91.405 ;
        RECT -1.770 -91.925 -1.310 -91.755 ;
        RECT 0.145 -92.260 0.315 -91.735 ;
        RECT 6.525 -92.260 6.695 -91.735 ;
        RECT 8.235 -91.755 8.525 -91.030 ;
        RECT 10.065 -91.405 10.235 -90.880 ;
        RECT 16.445 -91.405 16.615 -90.880 ;
        RECT 10.065 -91.735 10.615 -91.405 ;
        RECT 16.065 -91.735 16.615 -91.405 ;
        RECT 8.150 -91.925 8.610 -91.755 ;
        RECT 10.065 -92.260 10.235 -91.735 ;
        RECT 16.445 -92.260 16.615 -91.735 ;
        RECT 18.155 -91.755 18.445 -91.030 ;
        RECT 19.985 -91.405 20.155 -90.880 ;
        RECT 19.985 -91.735 20.535 -91.405 ;
        RECT 18.070 -91.925 18.530 -91.755 ;
        RECT 19.985 -92.260 20.155 -91.735 ;
        RECT -285.865 -174.155 -285.695 -173.630 ;
        RECT -284.240 -174.045 -283.780 -173.875 ;
        RECT -286.245 -174.485 -285.695 -174.155 ;
        RECT -285.865 -175.010 -285.695 -174.485 ;
        RECT -284.155 -174.770 -283.865 -174.045 ;
        RECT -282.325 -174.155 -282.155 -173.630 ;
        RECT -275.945 -174.155 -275.775 -173.630 ;
        RECT -274.320 -174.045 -273.860 -173.875 ;
        RECT -282.325 -174.485 -281.775 -174.155 ;
        RECT -276.325 -174.485 -275.775 -174.155 ;
        RECT -282.325 -175.010 -282.155 -174.485 ;
        RECT -275.945 -175.010 -275.775 -174.485 ;
        RECT -274.235 -174.770 -273.945 -174.045 ;
        RECT -272.405 -174.155 -272.235 -173.630 ;
        RECT -266.025 -174.155 -265.855 -173.630 ;
        RECT -264.400 -174.045 -263.940 -173.875 ;
        RECT -272.405 -174.485 -271.855 -174.155 ;
        RECT -266.405 -174.485 -265.855 -174.155 ;
        RECT -272.405 -175.010 -272.235 -174.485 ;
        RECT -266.025 -175.010 -265.855 -174.485 ;
        RECT -264.315 -174.770 -264.025 -174.045 ;
        RECT -262.485 -174.155 -262.315 -173.630 ;
        RECT -256.105 -174.155 -255.935 -173.630 ;
        RECT -254.480 -174.045 -254.020 -173.875 ;
        RECT -262.485 -174.485 -261.935 -174.155 ;
        RECT -256.485 -174.485 -255.935 -174.155 ;
        RECT -262.485 -175.010 -262.315 -174.485 ;
        RECT -256.105 -175.010 -255.935 -174.485 ;
        RECT -254.395 -174.770 -254.105 -174.045 ;
        RECT -252.565 -174.155 -252.395 -173.630 ;
        RECT -246.185 -174.155 -246.015 -173.630 ;
        RECT -244.560 -174.045 -244.100 -173.875 ;
        RECT -252.565 -174.485 -252.015 -174.155 ;
        RECT -246.565 -174.485 -246.015 -174.155 ;
        RECT -252.565 -175.010 -252.395 -174.485 ;
        RECT -246.185 -175.010 -246.015 -174.485 ;
        RECT -244.475 -174.770 -244.185 -174.045 ;
        RECT -242.645 -174.155 -242.475 -173.630 ;
        RECT -236.265 -174.155 -236.095 -173.630 ;
        RECT -234.640 -174.045 -234.180 -173.875 ;
        RECT -242.645 -174.485 -242.095 -174.155 ;
        RECT -236.645 -174.485 -236.095 -174.155 ;
        RECT -242.645 -175.010 -242.475 -174.485 ;
        RECT -236.265 -175.010 -236.095 -174.485 ;
        RECT -234.555 -174.770 -234.265 -174.045 ;
        RECT -232.725 -174.155 -232.555 -173.630 ;
        RECT -226.345 -174.155 -226.175 -173.630 ;
        RECT -224.720 -174.045 -224.260 -173.875 ;
        RECT -232.725 -174.485 -232.175 -174.155 ;
        RECT -226.725 -174.485 -226.175 -174.155 ;
        RECT -232.725 -175.010 -232.555 -174.485 ;
        RECT -226.345 -175.010 -226.175 -174.485 ;
        RECT -224.635 -174.770 -224.345 -174.045 ;
        RECT -222.805 -174.155 -222.635 -173.630 ;
        RECT -216.425 -174.155 -216.255 -173.630 ;
        RECT -214.800 -174.045 -214.340 -173.875 ;
        RECT -222.805 -174.485 -222.255 -174.155 ;
        RECT -216.805 -174.485 -216.255 -174.155 ;
        RECT -222.805 -175.010 -222.635 -174.485 ;
        RECT -216.425 -175.010 -216.255 -174.485 ;
        RECT -214.715 -174.770 -214.425 -174.045 ;
        RECT -212.885 -174.155 -212.715 -173.630 ;
        RECT -206.505 -174.155 -206.335 -173.630 ;
        RECT -204.880 -174.045 -204.420 -173.875 ;
        RECT -212.885 -174.485 -212.335 -174.155 ;
        RECT -206.885 -174.485 -206.335 -174.155 ;
        RECT -212.885 -175.010 -212.715 -174.485 ;
        RECT -206.505 -175.010 -206.335 -174.485 ;
        RECT -204.795 -174.770 -204.505 -174.045 ;
        RECT -202.965 -174.155 -202.795 -173.630 ;
        RECT -196.585 -174.155 -196.415 -173.630 ;
        RECT -194.960 -174.045 -194.500 -173.875 ;
        RECT -202.965 -174.485 -202.415 -174.155 ;
        RECT -196.965 -174.485 -196.415 -174.155 ;
        RECT -202.965 -175.010 -202.795 -174.485 ;
        RECT -196.585 -175.010 -196.415 -174.485 ;
        RECT -194.875 -174.770 -194.585 -174.045 ;
        RECT -193.045 -174.155 -192.875 -173.630 ;
        RECT -186.665 -174.155 -186.495 -173.630 ;
        RECT -185.040 -174.045 -184.580 -173.875 ;
        RECT -193.045 -174.485 -192.495 -174.155 ;
        RECT -187.045 -174.485 -186.495 -174.155 ;
        RECT -193.045 -175.010 -192.875 -174.485 ;
        RECT -186.665 -175.010 -186.495 -174.485 ;
        RECT -184.955 -174.770 -184.665 -174.045 ;
        RECT -183.125 -174.155 -182.955 -173.630 ;
        RECT -176.745 -174.155 -176.575 -173.630 ;
        RECT -175.120 -174.045 -174.660 -173.875 ;
        RECT -183.125 -174.485 -182.575 -174.155 ;
        RECT -177.125 -174.485 -176.575 -174.155 ;
        RECT -183.125 -175.010 -182.955 -174.485 ;
        RECT -176.745 -175.010 -176.575 -174.485 ;
        RECT -175.035 -174.770 -174.745 -174.045 ;
        RECT -173.205 -174.155 -173.035 -173.630 ;
        RECT -166.825 -174.155 -166.655 -173.630 ;
        RECT -165.200 -174.045 -164.740 -173.875 ;
        RECT -173.205 -174.485 -172.655 -174.155 ;
        RECT -167.205 -174.485 -166.655 -174.155 ;
        RECT -173.205 -175.010 -173.035 -174.485 ;
        RECT -166.825 -175.010 -166.655 -174.485 ;
        RECT -165.115 -174.770 -164.825 -174.045 ;
        RECT -163.285 -174.155 -163.115 -173.630 ;
        RECT -156.905 -174.155 -156.735 -173.630 ;
        RECT -155.280 -174.045 -154.820 -173.875 ;
        RECT -163.285 -174.485 -162.735 -174.155 ;
        RECT -157.285 -174.485 -156.735 -174.155 ;
        RECT -163.285 -175.010 -163.115 -174.485 ;
        RECT -156.905 -175.010 -156.735 -174.485 ;
        RECT -155.195 -174.770 -154.905 -174.045 ;
        RECT -153.365 -174.155 -153.195 -173.630 ;
        RECT -146.985 -174.155 -146.815 -173.630 ;
        RECT -145.360 -174.045 -144.900 -173.875 ;
        RECT -153.365 -174.485 -152.815 -174.155 ;
        RECT -147.365 -174.485 -146.815 -174.155 ;
        RECT -153.365 -175.010 -153.195 -174.485 ;
        RECT -146.985 -175.010 -146.815 -174.485 ;
        RECT -145.275 -174.770 -144.985 -174.045 ;
        RECT -143.445 -174.155 -143.275 -173.630 ;
        RECT -137.065 -174.155 -136.895 -173.630 ;
        RECT -135.440 -174.045 -134.980 -173.875 ;
        RECT -143.445 -174.485 -142.895 -174.155 ;
        RECT -137.445 -174.485 -136.895 -174.155 ;
        RECT -143.445 -175.010 -143.275 -174.485 ;
        RECT -137.065 -175.010 -136.895 -174.485 ;
        RECT -135.355 -174.770 -135.065 -174.045 ;
        RECT -133.525 -174.155 -133.355 -173.630 ;
        RECT -127.145 -174.155 -126.975 -173.630 ;
        RECT -125.520 -174.045 -125.060 -173.875 ;
        RECT -133.525 -174.485 -132.975 -174.155 ;
        RECT -127.525 -174.485 -126.975 -174.155 ;
        RECT -133.525 -175.010 -133.355 -174.485 ;
        RECT -127.145 -175.010 -126.975 -174.485 ;
        RECT -125.435 -174.770 -125.145 -174.045 ;
        RECT -123.605 -174.155 -123.435 -173.630 ;
        RECT -117.225 -174.155 -117.055 -173.630 ;
        RECT -115.600 -174.045 -115.140 -173.875 ;
        RECT -123.605 -174.485 -123.055 -174.155 ;
        RECT -117.605 -174.485 -117.055 -174.155 ;
        RECT -123.605 -175.010 -123.435 -174.485 ;
        RECT -117.225 -175.010 -117.055 -174.485 ;
        RECT -115.515 -174.770 -115.225 -174.045 ;
        RECT -113.685 -174.155 -113.515 -173.630 ;
        RECT -107.305 -174.155 -107.135 -173.630 ;
        RECT -105.680 -174.045 -105.220 -173.875 ;
        RECT -113.685 -174.485 -113.135 -174.155 ;
        RECT -107.685 -174.485 -107.135 -174.155 ;
        RECT -113.685 -175.010 -113.515 -174.485 ;
        RECT -107.305 -175.010 -107.135 -174.485 ;
        RECT -105.595 -174.770 -105.305 -174.045 ;
        RECT -103.765 -174.155 -103.595 -173.630 ;
        RECT -97.385 -174.155 -97.215 -173.630 ;
        RECT -95.760 -174.045 -95.300 -173.875 ;
        RECT -103.765 -174.485 -103.215 -174.155 ;
        RECT -97.765 -174.485 -97.215 -174.155 ;
        RECT -103.765 -175.010 -103.595 -174.485 ;
        RECT -97.385 -175.010 -97.215 -174.485 ;
        RECT -95.675 -174.770 -95.385 -174.045 ;
        RECT -93.845 -174.155 -93.675 -173.630 ;
        RECT -87.465 -174.155 -87.295 -173.630 ;
        RECT -85.840 -174.045 -85.380 -173.875 ;
        RECT -93.845 -174.485 -93.295 -174.155 ;
        RECT -87.845 -174.485 -87.295 -174.155 ;
        RECT -93.845 -175.010 -93.675 -174.485 ;
        RECT -87.465 -175.010 -87.295 -174.485 ;
        RECT -85.755 -174.770 -85.465 -174.045 ;
        RECT -83.925 -174.155 -83.755 -173.630 ;
        RECT -77.545 -174.155 -77.375 -173.630 ;
        RECT -75.920 -174.045 -75.460 -173.875 ;
        RECT -83.925 -174.485 -83.375 -174.155 ;
        RECT -77.925 -174.485 -77.375 -174.155 ;
        RECT -83.925 -175.010 -83.755 -174.485 ;
        RECT -77.545 -175.010 -77.375 -174.485 ;
        RECT -75.835 -174.770 -75.545 -174.045 ;
        RECT -74.005 -174.155 -73.835 -173.630 ;
        RECT -67.625 -174.155 -67.455 -173.630 ;
        RECT -66.000 -174.045 -65.540 -173.875 ;
        RECT -74.005 -174.485 -73.455 -174.155 ;
        RECT -68.005 -174.485 -67.455 -174.155 ;
        RECT -74.005 -175.010 -73.835 -174.485 ;
        RECT -67.625 -175.010 -67.455 -174.485 ;
        RECT -65.915 -174.770 -65.625 -174.045 ;
        RECT -64.085 -174.155 -63.915 -173.630 ;
        RECT -57.705 -174.155 -57.535 -173.630 ;
        RECT -56.080 -174.045 -55.620 -173.875 ;
        RECT -64.085 -174.485 -63.535 -174.155 ;
        RECT -58.085 -174.485 -57.535 -174.155 ;
        RECT -64.085 -175.010 -63.915 -174.485 ;
        RECT -57.705 -175.010 -57.535 -174.485 ;
        RECT -55.995 -174.770 -55.705 -174.045 ;
        RECT -54.165 -174.155 -53.995 -173.630 ;
        RECT -47.785 -174.155 -47.615 -173.630 ;
        RECT -46.160 -174.045 -45.700 -173.875 ;
        RECT -54.165 -174.485 -53.615 -174.155 ;
        RECT -48.165 -174.485 -47.615 -174.155 ;
        RECT -54.165 -175.010 -53.995 -174.485 ;
        RECT -47.785 -175.010 -47.615 -174.485 ;
        RECT -46.075 -174.770 -45.785 -174.045 ;
        RECT -44.245 -174.155 -44.075 -173.630 ;
        RECT -37.865 -174.155 -37.695 -173.630 ;
        RECT -36.240 -174.045 -35.780 -173.875 ;
        RECT -44.245 -174.485 -43.695 -174.155 ;
        RECT -38.245 -174.485 -37.695 -174.155 ;
        RECT -44.245 -175.010 -44.075 -174.485 ;
        RECT -37.865 -175.010 -37.695 -174.485 ;
        RECT -36.155 -174.770 -35.865 -174.045 ;
        RECT -34.325 -174.155 -34.155 -173.630 ;
        RECT -27.945 -174.155 -27.775 -173.630 ;
        RECT -26.320 -174.045 -25.860 -173.875 ;
        RECT -34.325 -174.485 -33.775 -174.155 ;
        RECT -28.325 -174.485 -27.775 -174.155 ;
        RECT -34.325 -175.010 -34.155 -174.485 ;
        RECT -27.945 -175.010 -27.775 -174.485 ;
        RECT -26.235 -174.770 -25.945 -174.045 ;
        RECT -24.405 -174.155 -24.235 -173.630 ;
        RECT -18.025 -174.155 -17.855 -173.630 ;
        RECT -16.400 -174.045 -15.940 -173.875 ;
        RECT -24.405 -174.485 -23.855 -174.155 ;
        RECT -18.405 -174.485 -17.855 -174.155 ;
        RECT -24.405 -175.010 -24.235 -174.485 ;
        RECT -18.025 -175.010 -17.855 -174.485 ;
        RECT -16.315 -174.770 -16.025 -174.045 ;
        RECT -14.485 -174.155 -14.315 -173.630 ;
        RECT -8.105 -174.155 -7.935 -173.630 ;
        RECT -6.480 -174.045 -6.020 -173.875 ;
        RECT -14.485 -174.485 -13.935 -174.155 ;
        RECT -8.485 -174.485 -7.935 -174.155 ;
        RECT -14.485 -175.010 -14.315 -174.485 ;
        RECT -8.105 -175.010 -7.935 -174.485 ;
        RECT -6.395 -174.770 -6.105 -174.045 ;
        RECT -4.565 -174.155 -4.395 -173.630 ;
        RECT 1.815 -174.155 1.985 -173.630 ;
        RECT 3.440 -174.045 3.900 -173.875 ;
        RECT -4.565 -174.485 -4.015 -174.155 ;
        RECT 1.435 -174.485 1.985 -174.155 ;
        RECT -4.565 -175.010 -4.395 -174.485 ;
        RECT 1.815 -175.010 1.985 -174.485 ;
        RECT 3.525 -174.770 3.815 -174.045 ;
        RECT 5.355 -174.155 5.525 -173.630 ;
        RECT 11.735 -174.155 11.905 -173.630 ;
        RECT 13.360 -174.045 13.820 -173.875 ;
        RECT 5.355 -174.485 5.905 -174.155 ;
        RECT 11.355 -174.485 11.905 -174.155 ;
        RECT 5.355 -175.010 5.525 -174.485 ;
        RECT 11.735 -175.010 11.905 -174.485 ;
        RECT 13.445 -174.770 13.735 -174.045 ;
        RECT 15.275 -174.155 15.445 -173.630 ;
        RECT 21.655 -174.155 21.825 -173.630 ;
        RECT 23.280 -174.045 23.740 -173.875 ;
        RECT 15.275 -174.485 15.825 -174.155 ;
        RECT 21.275 -174.485 21.825 -174.155 ;
        RECT 15.275 -175.010 15.445 -174.485 ;
        RECT 21.655 -175.010 21.825 -174.485 ;
        RECT 23.365 -174.770 23.655 -174.045 ;
        RECT 25.195 -174.155 25.365 -173.630 ;
        RECT 25.195 -174.485 25.745 -174.155 ;
        RECT 25.195 -175.010 25.365 -174.485 ;
        RECT -280.660 -175.525 -277.440 -175.355 ;
        RECT -270.740 -175.525 -267.520 -175.355 ;
        RECT -260.820 -175.525 -257.600 -175.355 ;
        RECT -250.900 -175.525 -247.680 -175.355 ;
        RECT -240.980 -175.525 -237.760 -175.355 ;
        RECT -231.060 -175.525 -227.840 -175.355 ;
        RECT -221.140 -175.525 -217.920 -175.355 ;
        RECT -211.220 -175.525 -208.000 -175.355 ;
        RECT -201.300 -175.525 -198.080 -175.355 ;
        RECT -191.380 -175.525 -188.160 -175.355 ;
        RECT -181.460 -175.525 -178.240 -175.355 ;
        RECT -171.540 -175.525 -168.320 -175.355 ;
        RECT -161.620 -175.525 -158.400 -175.355 ;
        RECT -151.700 -175.525 -148.480 -175.355 ;
        RECT -141.780 -175.525 -138.560 -175.355 ;
        RECT -131.860 -175.525 -128.640 -175.355 ;
        RECT -121.940 -175.525 -118.720 -175.355 ;
        RECT -112.020 -175.525 -108.800 -175.355 ;
        RECT -102.100 -175.525 -98.880 -175.355 ;
        RECT -92.180 -175.525 -88.960 -175.355 ;
        RECT -82.260 -175.525 -79.040 -175.355 ;
        RECT -72.340 -175.525 -69.120 -175.355 ;
        RECT -62.420 -175.525 -59.200 -175.355 ;
        RECT -52.500 -175.525 -49.280 -175.355 ;
        RECT -42.580 -175.525 -39.360 -175.355 ;
        RECT -32.660 -175.525 -29.440 -175.355 ;
        RECT -22.740 -175.525 -19.520 -175.355 ;
        RECT -12.820 -175.525 -9.600 -175.355 ;
        RECT -2.900 -175.525 0.320 -175.355 ;
        RECT 7.020 -175.525 10.240 -175.355 ;
        RECT 16.940 -175.525 20.160 -175.355 ;
        RECT -279.675 -176.325 -279.365 -175.525 ;
        RECT -279.195 -176.250 -278.905 -175.525 ;
        RECT -278.735 -176.325 -278.425 -175.525 ;
        RECT -269.755 -176.325 -269.445 -175.525 ;
        RECT -269.275 -176.250 -268.985 -175.525 ;
        RECT -268.815 -176.325 -268.505 -175.525 ;
        RECT -259.835 -176.325 -259.525 -175.525 ;
        RECT -259.355 -176.250 -259.065 -175.525 ;
        RECT -258.895 -176.325 -258.585 -175.525 ;
        RECT -249.915 -176.325 -249.605 -175.525 ;
        RECT -249.435 -176.250 -249.145 -175.525 ;
        RECT -248.975 -176.325 -248.665 -175.525 ;
        RECT -239.995 -176.325 -239.685 -175.525 ;
        RECT -239.515 -176.250 -239.225 -175.525 ;
        RECT -239.055 -176.325 -238.745 -175.525 ;
        RECT -230.075 -176.325 -229.765 -175.525 ;
        RECT -229.595 -176.250 -229.305 -175.525 ;
        RECT -229.135 -176.325 -228.825 -175.525 ;
        RECT -220.155 -176.325 -219.845 -175.525 ;
        RECT -219.675 -176.250 -219.385 -175.525 ;
        RECT -219.215 -176.325 -218.905 -175.525 ;
        RECT -210.235 -176.325 -209.925 -175.525 ;
        RECT -209.755 -176.250 -209.465 -175.525 ;
        RECT -209.295 -176.325 -208.985 -175.525 ;
        RECT -200.315 -176.325 -200.005 -175.525 ;
        RECT -199.835 -176.250 -199.545 -175.525 ;
        RECT -199.375 -176.325 -199.065 -175.525 ;
        RECT -190.395 -176.325 -190.085 -175.525 ;
        RECT -189.915 -176.250 -189.625 -175.525 ;
        RECT -189.455 -176.325 -189.145 -175.525 ;
        RECT -180.475 -176.325 -180.165 -175.525 ;
        RECT -179.995 -176.250 -179.705 -175.525 ;
        RECT -179.535 -176.325 -179.225 -175.525 ;
        RECT -170.555 -176.325 -170.245 -175.525 ;
        RECT -170.075 -176.250 -169.785 -175.525 ;
        RECT -169.615 -176.325 -169.305 -175.525 ;
        RECT -160.635 -176.325 -160.325 -175.525 ;
        RECT -160.155 -176.250 -159.865 -175.525 ;
        RECT -159.695 -176.325 -159.385 -175.525 ;
        RECT -150.715 -176.325 -150.405 -175.525 ;
        RECT -150.235 -176.250 -149.945 -175.525 ;
        RECT -149.775 -176.325 -149.465 -175.525 ;
        RECT -140.795 -176.325 -140.485 -175.525 ;
        RECT -140.315 -176.250 -140.025 -175.525 ;
        RECT -139.855 -176.325 -139.545 -175.525 ;
        RECT -130.875 -176.325 -130.565 -175.525 ;
        RECT -130.395 -176.250 -130.105 -175.525 ;
        RECT -129.935 -176.325 -129.625 -175.525 ;
        RECT -120.955 -176.325 -120.645 -175.525 ;
        RECT -120.475 -176.250 -120.185 -175.525 ;
        RECT -120.015 -176.325 -119.705 -175.525 ;
        RECT -111.035 -176.325 -110.725 -175.525 ;
        RECT -110.555 -176.250 -110.265 -175.525 ;
        RECT -110.095 -176.325 -109.785 -175.525 ;
        RECT -101.115 -176.325 -100.805 -175.525 ;
        RECT -100.635 -176.250 -100.345 -175.525 ;
        RECT -100.175 -176.325 -99.865 -175.525 ;
        RECT -91.195 -176.325 -90.885 -175.525 ;
        RECT -90.715 -176.250 -90.425 -175.525 ;
        RECT -90.255 -176.325 -89.945 -175.525 ;
        RECT -81.275 -176.325 -80.965 -175.525 ;
        RECT -80.795 -176.250 -80.505 -175.525 ;
        RECT -80.335 -176.325 -80.025 -175.525 ;
        RECT -71.355 -176.325 -71.045 -175.525 ;
        RECT -70.875 -176.250 -70.585 -175.525 ;
        RECT -70.415 -176.325 -70.105 -175.525 ;
        RECT -61.435 -176.325 -61.125 -175.525 ;
        RECT -60.955 -176.250 -60.665 -175.525 ;
        RECT -60.495 -176.325 -60.185 -175.525 ;
        RECT -51.515 -176.325 -51.205 -175.525 ;
        RECT -51.035 -176.250 -50.745 -175.525 ;
        RECT -50.575 -176.325 -50.265 -175.525 ;
        RECT -41.595 -176.325 -41.285 -175.525 ;
        RECT -41.115 -176.250 -40.825 -175.525 ;
        RECT -40.655 -176.325 -40.345 -175.525 ;
        RECT -31.675 -176.325 -31.365 -175.525 ;
        RECT -31.195 -176.250 -30.905 -175.525 ;
        RECT -30.735 -176.325 -30.425 -175.525 ;
        RECT -21.755 -176.325 -21.445 -175.525 ;
        RECT -21.275 -176.250 -20.985 -175.525 ;
        RECT -20.815 -176.325 -20.505 -175.525 ;
        RECT -11.835 -176.325 -11.525 -175.525 ;
        RECT -11.355 -176.250 -11.065 -175.525 ;
        RECT -10.895 -176.325 -10.585 -175.525 ;
        RECT -1.915 -176.325 -1.605 -175.525 ;
        RECT -1.435 -176.250 -1.145 -175.525 ;
        RECT -0.975 -176.325 -0.665 -175.525 ;
        RECT 8.005 -176.325 8.315 -175.525 ;
        RECT 8.485 -176.250 8.775 -175.525 ;
        RECT 8.945 -176.325 9.255 -175.525 ;
        RECT 17.925 -176.325 18.235 -175.525 ;
        RECT 18.405 -176.250 18.695 -175.525 ;
        RECT 18.865 -176.325 19.175 -175.525 ;
        RECT -284.635 -178.075 -284.325 -177.275 ;
        RECT -284.155 -178.075 -283.865 -177.350 ;
        RECT -283.695 -178.075 -283.385 -177.275 ;
        RECT -274.715 -178.075 -274.405 -177.275 ;
        RECT -274.235 -178.075 -273.945 -177.350 ;
        RECT -273.775 -178.075 -273.465 -177.275 ;
        RECT -264.795 -178.075 -264.485 -177.275 ;
        RECT -264.315 -178.075 -264.025 -177.350 ;
        RECT -263.855 -178.075 -263.545 -177.275 ;
        RECT -254.875 -178.075 -254.565 -177.275 ;
        RECT -254.395 -178.075 -254.105 -177.350 ;
        RECT -253.935 -178.075 -253.625 -177.275 ;
        RECT -244.955 -178.075 -244.645 -177.275 ;
        RECT -244.475 -178.075 -244.185 -177.350 ;
        RECT -244.015 -178.075 -243.705 -177.275 ;
        RECT -235.035 -178.075 -234.725 -177.275 ;
        RECT -234.555 -178.075 -234.265 -177.350 ;
        RECT -234.095 -178.075 -233.785 -177.275 ;
        RECT -225.115 -178.075 -224.805 -177.275 ;
        RECT -224.635 -178.075 -224.345 -177.350 ;
        RECT -224.175 -178.075 -223.865 -177.275 ;
        RECT -215.195 -178.075 -214.885 -177.275 ;
        RECT -214.715 -178.075 -214.425 -177.350 ;
        RECT -214.255 -178.075 -213.945 -177.275 ;
        RECT -205.275 -178.075 -204.965 -177.275 ;
        RECT -204.795 -178.075 -204.505 -177.350 ;
        RECT -204.335 -178.075 -204.025 -177.275 ;
        RECT -195.355 -178.075 -195.045 -177.275 ;
        RECT -194.875 -178.075 -194.585 -177.350 ;
        RECT -194.415 -178.075 -194.105 -177.275 ;
        RECT -185.435 -178.075 -185.125 -177.275 ;
        RECT -184.955 -178.075 -184.665 -177.350 ;
        RECT -184.495 -178.075 -184.185 -177.275 ;
        RECT -175.515 -178.075 -175.205 -177.275 ;
        RECT -175.035 -178.075 -174.745 -177.350 ;
        RECT -174.575 -178.075 -174.265 -177.275 ;
        RECT -165.595 -178.075 -165.285 -177.275 ;
        RECT -165.115 -178.075 -164.825 -177.350 ;
        RECT -164.655 -178.075 -164.345 -177.275 ;
        RECT -155.675 -178.075 -155.365 -177.275 ;
        RECT -155.195 -178.075 -154.905 -177.350 ;
        RECT -154.735 -178.075 -154.425 -177.275 ;
        RECT -145.755 -178.075 -145.445 -177.275 ;
        RECT -145.275 -178.075 -144.985 -177.350 ;
        RECT -144.815 -178.075 -144.505 -177.275 ;
        RECT -135.835 -178.075 -135.525 -177.275 ;
        RECT -135.355 -178.075 -135.065 -177.350 ;
        RECT -134.895 -178.075 -134.585 -177.275 ;
        RECT -125.915 -178.075 -125.605 -177.275 ;
        RECT -125.435 -178.075 -125.145 -177.350 ;
        RECT -124.975 -178.075 -124.665 -177.275 ;
        RECT -115.995 -178.075 -115.685 -177.275 ;
        RECT -115.515 -178.075 -115.225 -177.350 ;
        RECT -115.055 -178.075 -114.745 -177.275 ;
        RECT -106.075 -178.075 -105.765 -177.275 ;
        RECT -105.595 -178.075 -105.305 -177.350 ;
        RECT -105.135 -178.075 -104.825 -177.275 ;
        RECT -96.155 -178.075 -95.845 -177.275 ;
        RECT -95.675 -178.075 -95.385 -177.350 ;
        RECT -95.215 -178.075 -94.905 -177.275 ;
        RECT -86.235 -178.075 -85.925 -177.275 ;
        RECT -85.755 -178.075 -85.465 -177.350 ;
        RECT -85.295 -178.075 -84.985 -177.275 ;
        RECT -76.315 -178.075 -76.005 -177.275 ;
        RECT -75.835 -178.075 -75.545 -177.350 ;
        RECT -75.375 -178.075 -75.065 -177.275 ;
        RECT -66.395 -178.075 -66.085 -177.275 ;
        RECT -65.915 -178.075 -65.625 -177.350 ;
        RECT -65.455 -178.075 -65.145 -177.275 ;
        RECT -56.475 -178.075 -56.165 -177.275 ;
        RECT -55.995 -178.075 -55.705 -177.350 ;
        RECT -55.535 -178.075 -55.225 -177.275 ;
        RECT -46.555 -178.075 -46.245 -177.275 ;
        RECT -46.075 -178.075 -45.785 -177.350 ;
        RECT -45.615 -178.075 -45.305 -177.275 ;
        RECT -36.635 -178.075 -36.325 -177.275 ;
        RECT -36.155 -178.075 -35.865 -177.350 ;
        RECT -35.695 -178.075 -35.385 -177.275 ;
        RECT -26.715 -178.075 -26.405 -177.275 ;
        RECT -26.235 -178.075 -25.945 -177.350 ;
        RECT -25.775 -178.075 -25.465 -177.275 ;
        RECT -16.795 -178.075 -16.485 -177.275 ;
        RECT -16.315 -178.075 -16.025 -177.350 ;
        RECT -15.855 -178.075 -15.545 -177.275 ;
        RECT -6.875 -178.075 -6.565 -177.275 ;
        RECT -6.395 -178.075 -6.105 -177.350 ;
        RECT -5.935 -178.075 -5.625 -177.275 ;
        RECT 3.045 -178.075 3.355 -177.275 ;
        RECT 3.525 -178.075 3.815 -177.350 ;
        RECT 3.985 -178.075 4.295 -177.275 ;
        RECT 12.965 -178.075 13.275 -177.275 ;
        RECT 13.445 -178.075 13.735 -177.350 ;
        RECT 13.905 -178.075 14.215 -177.275 ;
        RECT 22.885 -178.075 23.195 -177.275 ;
        RECT 23.365 -178.075 23.655 -177.350 ;
        RECT 23.825 -178.075 24.135 -177.275 ;
        RECT -285.620 -178.245 -282.400 -178.075 ;
        RECT -275.700 -178.245 -272.480 -178.075 ;
        RECT -265.780 -178.245 -262.560 -178.075 ;
        RECT -255.860 -178.245 -252.640 -178.075 ;
        RECT -245.940 -178.245 -242.720 -178.075 ;
        RECT -236.020 -178.245 -232.800 -178.075 ;
        RECT -226.100 -178.245 -222.880 -178.075 ;
        RECT -216.180 -178.245 -212.960 -178.075 ;
        RECT -206.260 -178.245 -203.040 -178.075 ;
        RECT -196.340 -178.245 -193.120 -178.075 ;
        RECT -186.420 -178.245 -183.200 -178.075 ;
        RECT -176.500 -178.245 -173.280 -178.075 ;
        RECT -166.580 -178.245 -163.360 -178.075 ;
        RECT -156.660 -178.245 -153.440 -178.075 ;
        RECT -146.740 -178.245 -143.520 -178.075 ;
        RECT -136.820 -178.245 -133.600 -178.075 ;
        RECT -126.900 -178.245 -123.680 -178.075 ;
        RECT -116.980 -178.245 -113.760 -178.075 ;
        RECT -107.060 -178.245 -103.840 -178.075 ;
        RECT -97.140 -178.245 -93.920 -178.075 ;
        RECT -87.220 -178.245 -84.000 -178.075 ;
        RECT -77.300 -178.245 -74.080 -178.075 ;
        RECT -67.380 -178.245 -64.160 -178.075 ;
        RECT -57.460 -178.245 -54.240 -178.075 ;
        RECT -47.540 -178.245 -44.320 -178.075 ;
        RECT -37.620 -178.245 -34.400 -178.075 ;
        RECT -27.700 -178.245 -24.480 -178.075 ;
        RECT -17.780 -178.245 -14.560 -178.075 ;
        RECT -7.860 -178.245 -4.640 -178.075 ;
        RECT 2.060 -178.245 5.280 -178.075 ;
        RECT 11.980 -178.245 15.200 -178.075 ;
        RECT 21.900 -178.245 25.120 -178.075 ;
        RECT -280.905 -179.115 -280.735 -178.590 ;
        RECT -281.285 -179.445 -280.735 -179.115 ;
        RECT -280.905 -179.970 -280.735 -179.445 ;
        RECT -279.195 -179.465 -278.905 -178.740 ;
        RECT -277.365 -179.115 -277.195 -178.590 ;
        RECT -270.985 -179.115 -270.815 -178.590 ;
        RECT -277.365 -179.445 -276.815 -179.115 ;
        RECT -271.365 -179.445 -270.815 -179.115 ;
        RECT -279.280 -179.635 -278.820 -179.465 ;
        RECT -277.365 -179.970 -277.195 -179.445 ;
        RECT -270.985 -179.970 -270.815 -179.445 ;
        RECT -269.275 -179.465 -268.985 -178.740 ;
        RECT -267.445 -179.115 -267.275 -178.590 ;
        RECT -261.065 -179.115 -260.895 -178.590 ;
        RECT -267.445 -179.445 -266.895 -179.115 ;
        RECT -261.445 -179.445 -260.895 -179.115 ;
        RECT -269.360 -179.635 -268.900 -179.465 ;
        RECT -267.445 -179.970 -267.275 -179.445 ;
        RECT -261.065 -179.970 -260.895 -179.445 ;
        RECT -259.355 -179.465 -259.065 -178.740 ;
        RECT -257.525 -179.115 -257.355 -178.590 ;
        RECT -251.145 -179.115 -250.975 -178.590 ;
        RECT -257.525 -179.445 -256.975 -179.115 ;
        RECT -251.525 -179.445 -250.975 -179.115 ;
        RECT -259.440 -179.635 -258.980 -179.465 ;
        RECT -257.525 -179.970 -257.355 -179.445 ;
        RECT -251.145 -179.970 -250.975 -179.445 ;
        RECT -249.435 -179.465 -249.145 -178.740 ;
        RECT -247.605 -179.115 -247.435 -178.590 ;
        RECT -241.225 -179.115 -241.055 -178.590 ;
        RECT -247.605 -179.445 -247.055 -179.115 ;
        RECT -241.605 -179.445 -241.055 -179.115 ;
        RECT -249.520 -179.635 -249.060 -179.465 ;
        RECT -247.605 -179.970 -247.435 -179.445 ;
        RECT -241.225 -179.970 -241.055 -179.445 ;
        RECT -239.515 -179.465 -239.225 -178.740 ;
        RECT -237.685 -179.115 -237.515 -178.590 ;
        RECT -231.305 -179.115 -231.135 -178.590 ;
        RECT -237.685 -179.445 -237.135 -179.115 ;
        RECT -231.685 -179.445 -231.135 -179.115 ;
        RECT -239.600 -179.635 -239.140 -179.465 ;
        RECT -237.685 -179.970 -237.515 -179.445 ;
        RECT -231.305 -179.970 -231.135 -179.445 ;
        RECT -229.595 -179.465 -229.305 -178.740 ;
        RECT -227.765 -179.115 -227.595 -178.590 ;
        RECT -221.385 -179.115 -221.215 -178.590 ;
        RECT -227.765 -179.445 -227.215 -179.115 ;
        RECT -221.765 -179.445 -221.215 -179.115 ;
        RECT -229.680 -179.635 -229.220 -179.465 ;
        RECT -227.765 -179.970 -227.595 -179.445 ;
        RECT -221.385 -179.970 -221.215 -179.445 ;
        RECT -219.675 -179.465 -219.385 -178.740 ;
        RECT -217.845 -179.115 -217.675 -178.590 ;
        RECT -211.465 -179.115 -211.295 -178.590 ;
        RECT -217.845 -179.445 -217.295 -179.115 ;
        RECT -211.845 -179.445 -211.295 -179.115 ;
        RECT -219.760 -179.635 -219.300 -179.465 ;
        RECT -217.845 -179.970 -217.675 -179.445 ;
        RECT -211.465 -179.970 -211.295 -179.445 ;
        RECT -209.755 -179.465 -209.465 -178.740 ;
        RECT -207.925 -179.115 -207.755 -178.590 ;
        RECT -201.545 -179.115 -201.375 -178.590 ;
        RECT -207.925 -179.445 -207.375 -179.115 ;
        RECT -201.925 -179.445 -201.375 -179.115 ;
        RECT -209.840 -179.635 -209.380 -179.465 ;
        RECT -207.925 -179.970 -207.755 -179.445 ;
        RECT -201.545 -179.970 -201.375 -179.445 ;
        RECT -199.835 -179.465 -199.545 -178.740 ;
        RECT -198.005 -179.115 -197.835 -178.590 ;
        RECT -191.625 -179.115 -191.455 -178.590 ;
        RECT -198.005 -179.445 -197.455 -179.115 ;
        RECT -192.005 -179.445 -191.455 -179.115 ;
        RECT -199.920 -179.635 -199.460 -179.465 ;
        RECT -198.005 -179.970 -197.835 -179.445 ;
        RECT -191.625 -179.970 -191.455 -179.445 ;
        RECT -189.915 -179.465 -189.625 -178.740 ;
        RECT -188.085 -179.115 -187.915 -178.590 ;
        RECT -181.705 -179.115 -181.535 -178.590 ;
        RECT -188.085 -179.445 -187.535 -179.115 ;
        RECT -182.085 -179.445 -181.535 -179.115 ;
        RECT -190.000 -179.635 -189.540 -179.465 ;
        RECT -188.085 -179.970 -187.915 -179.445 ;
        RECT -181.705 -179.970 -181.535 -179.445 ;
        RECT -179.995 -179.465 -179.705 -178.740 ;
        RECT -178.165 -179.115 -177.995 -178.590 ;
        RECT -171.785 -179.115 -171.615 -178.590 ;
        RECT -178.165 -179.445 -177.615 -179.115 ;
        RECT -172.165 -179.445 -171.615 -179.115 ;
        RECT -180.080 -179.635 -179.620 -179.465 ;
        RECT -178.165 -179.970 -177.995 -179.445 ;
        RECT -171.785 -179.970 -171.615 -179.445 ;
        RECT -170.075 -179.465 -169.785 -178.740 ;
        RECT -168.245 -179.115 -168.075 -178.590 ;
        RECT -161.865 -179.115 -161.695 -178.590 ;
        RECT -168.245 -179.445 -167.695 -179.115 ;
        RECT -162.245 -179.445 -161.695 -179.115 ;
        RECT -170.160 -179.635 -169.700 -179.465 ;
        RECT -168.245 -179.970 -168.075 -179.445 ;
        RECT -161.865 -179.970 -161.695 -179.445 ;
        RECT -160.155 -179.465 -159.865 -178.740 ;
        RECT -158.325 -179.115 -158.155 -178.590 ;
        RECT -151.945 -179.115 -151.775 -178.590 ;
        RECT -158.325 -179.445 -157.775 -179.115 ;
        RECT -152.325 -179.445 -151.775 -179.115 ;
        RECT -160.240 -179.635 -159.780 -179.465 ;
        RECT -158.325 -179.970 -158.155 -179.445 ;
        RECT -151.945 -179.970 -151.775 -179.445 ;
        RECT -150.235 -179.465 -149.945 -178.740 ;
        RECT -148.405 -179.115 -148.235 -178.590 ;
        RECT -142.025 -179.115 -141.855 -178.590 ;
        RECT -148.405 -179.445 -147.855 -179.115 ;
        RECT -142.405 -179.445 -141.855 -179.115 ;
        RECT -150.320 -179.635 -149.860 -179.465 ;
        RECT -148.405 -179.970 -148.235 -179.445 ;
        RECT -142.025 -179.970 -141.855 -179.445 ;
        RECT -140.315 -179.465 -140.025 -178.740 ;
        RECT -138.485 -179.115 -138.315 -178.590 ;
        RECT -132.105 -179.115 -131.935 -178.590 ;
        RECT -138.485 -179.445 -137.935 -179.115 ;
        RECT -132.485 -179.445 -131.935 -179.115 ;
        RECT -140.400 -179.635 -139.940 -179.465 ;
        RECT -138.485 -179.970 -138.315 -179.445 ;
        RECT -132.105 -179.970 -131.935 -179.445 ;
        RECT -130.395 -179.465 -130.105 -178.740 ;
        RECT -128.565 -179.115 -128.395 -178.590 ;
        RECT -122.185 -179.115 -122.015 -178.590 ;
        RECT -128.565 -179.445 -128.015 -179.115 ;
        RECT -122.565 -179.445 -122.015 -179.115 ;
        RECT -130.480 -179.635 -130.020 -179.465 ;
        RECT -128.565 -179.970 -128.395 -179.445 ;
        RECT -122.185 -179.970 -122.015 -179.445 ;
        RECT -120.475 -179.465 -120.185 -178.740 ;
        RECT -118.645 -179.115 -118.475 -178.590 ;
        RECT -112.265 -179.115 -112.095 -178.590 ;
        RECT -118.645 -179.445 -118.095 -179.115 ;
        RECT -112.645 -179.445 -112.095 -179.115 ;
        RECT -120.560 -179.635 -120.100 -179.465 ;
        RECT -118.645 -179.970 -118.475 -179.445 ;
        RECT -112.265 -179.970 -112.095 -179.445 ;
        RECT -110.555 -179.465 -110.265 -178.740 ;
        RECT -108.725 -179.115 -108.555 -178.590 ;
        RECT -102.345 -179.115 -102.175 -178.590 ;
        RECT -108.725 -179.445 -108.175 -179.115 ;
        RECT -102.725 -179.445 -102.175 -179.115 ;
        RECT -110.640 -179.635 -110.180 -179.465 ;
        RECT -108.725 -179.970 -108.555 -179.445 ;
        RECT -102.345 -179.970 -102.175 -179.445 ;
        RECT -100.635 -179.465 -100.345 -178.740 ;
        RECT -98.805 -179.115 -98.635 -178.590 ;
        RECT -92.425 -179.115 -92.255 -178.590 ;
        RECT -98.805 -179.445 -98.255 -179.115 ;
        RECT -92.805 -179.445 -92.255 -179.115 ;
        RECT -100.720 -179.635 -100.260 -179.465 ;
        RECT -98.805 -179.970 -98.635 -179.445 ;
        RECT -92.425 -179.970 -92.255 -179.445 ;
        RECT -90.715 -179.465 -90.425 -178.740 ;
        RECT -88.885 -179.115 -88.715 -178.590 ;
        RECT -82.505 -179.115 -82.335 -178.590 ;
        RECT -88.885 -179.445 -88.335 -179.115 ;
        RECT -82.885 -179.445 -82.335 -179.115 ;
        RECT -90.800 -179.635 -90.340 -179.465 ;
        RECT -88.885 -179.970 -88.715 -179.445 ;
        RECT -82.505 -179.970 -82.335 -179.445 ;
        RECT -80.795 -179.465 -80.505 -178.740 ;
        RECT -78.965 -179.115 -78.795 -178.590 ;
        RECT -72.585 -179.115 -72.415 -178.590 ;
        RECT -78.965 -179.445 -78.415 -179.115 ;
        RECT -72.965 -179.445 -72.415 -179.115 ;
        RECT -80.880 -179.635 -80.420 -179.465 ;
        RECT -78.965 -179.970 -78.795 -179.445 ;
        RECT -72.585 -179.970 -72.415 -179.445 ;
        RECT -70.875 -179.465 -70.585 -178.740 ;
        RECT -69.045 -179.115 -68.875 -178.590 ;
        RECT -62.665 -179.115 -62.495 -178.590 ;
        RECT -69.045 -179.445 -68.495 -179.115 ;
        RECT -63.045 -179.445 -62.495 -179.115 ;
        RECT -70.960 -179.635 -70.500 -179.465 ;
        RECT -69.045 -179.970 -68.875 -179.445 ;
        RECT -62.665 -179.970 -62.495 -179.445 ;
        RECT -60.955 -179.465 -60.665 -178.740 ;
        RECT -59.125 -179.115 -58.955 -178.590 ;
        RECT -52.745 -179.115 -52.575 -178.590 ;
        RECT -59.125 -179.445 -58.575 -179.115 ;
        RECT -53.125 -179.445 -52.575 -179.115 ;
        RECT -61.040 -179.635 -60.580 -179.465 ;
        RECT -59.125 -179.970 -58.955 -179.445 ;
        RECT -52.745 -179.970 -52.575 -179.445 ;
        RECT -51.035 -179.465 -50.745 -178.740 ;
        RECT -49.205 -179.115 -49.035 -178.590 ;
        RECT -42.825 -179.115 -42.655 -178.590 ;
        RECT -49.205 -179.445 -48.655 -179.115 ;
        RECT -43.205 -179.445 -42.655 -179.115 ;
        RECT -51.120 -179.635 -50.660 -179.465 ;
        RECT -49.205 -179.970 -49.035 -179.445 ;
        RECT -42.825 -179.970 -42.655 -179.445 ;
        RECT -41.115 -179.465 -40.825 -178.740 ;
        RECT -39.285 -179.115 -39.115 -178.590 ;
        RECT -32.905 -179.115 -32.735 -178.590 ;
        RECT -39.285 -179.445 -38.735 -179.115 ;
        RECT -33.285 -179.445 -32.735 -179.115 ;
        RECT -41.200 -179.635 -40.740 -179.465 ;
        RECT -39.285 -179.970 -39.115 -179.445 ;
        RECT -32.905 -179.970 -32.735 -179.445 ;
        RECT -31.195 -179.465 -30.905 -178.740 ;
        RECT -29.365 -179.115 -29.195 -178.590 ;
        RECT -22.985 -179.115 -22.815 -178.590 ;
        RECT -29.365 -179.445 -28.815 -179.115 ;
        RECT -23.365 -179.445 -22.815 -179.115 ;
        RECT -31.280 -179.635 -30.820 -179.465 ;
        RECT -29.365 -179.970 -29.195 -179.445 ;
        RECT -22.985 -179.970 -22.815 -179.445 ;
        RECT -21.275 -179.465 -20.985 -178.740 ;
        RECT -19.445 -179.115 -19.275 -178.590 ;
        RECT -13.065 -179.115 -12.895 -178.590 ;
        RECT -19.445 -179.445 -18.895 -179.115 ;
        RECT -13.445 -179.445 -12.895 -179.115 ;
        RECT -21.360 -179.635 -20.900 -179.465 ;
        RECT -19.445 -179.970 -19.275 -179.445 ;
        RECT -13.065 -179.970 -12.895 -179.445 ;
        RECT -11.355 -179.465 -11.065 -178.740 ;
        RECT -9.525 -179.115 -9.355 -178.590 ;
        RECT -3.145 -179.115 -2.975 -178.590 ;
        RECT -9.525 -179.445 -8.975 -179.115 ;
        RECT -3.525 -179.445 -2.975 -179.115 ;
        RECT -11.440 -179.635 -10.980 -179.465 ;
        RECT -9.525 -179.970 -9.355 -179.445 ;
        RECT -3.145 -179.970 -2.975 -179.445 ;
        RECT -1.435 -179.465 -1.145 -178.740 ;
        RECT 0.395 -179.115 0.565 -178.590 ;
        RECT 6.775 -179.115 6.945 -178.590 ;
        RECT 0.395 -179.445 0.945 -179.115 ;
        RECT 6.395 -179.445 6.945 -179.115 ;
        RECT -1.520 -179.635 -1.060 -179.465 ;
        RECT 0.395 -179.970 0.565 -179.445 ;
        RECT 6.775 -179.970 6.945 -179.445 ;
        RECT 8.485 -179.465 8.775 -178.740 ;
        RECT 10.315 -179.115 10.485 -178.590 ;
        RECT 16.695 -179.115 16.865 -178.590 ;
        RECT 10.315 -179.445 10.865 -179.115 ;
        RECT 16.315 -179.445 16.865 -179.115 ;
        RECT 8.400 -179.635 8.860 -179.465 ;
        RECT 10.315 -179.970 10.485 -179.445 ;
        RECT 16.695 -179.970 16.865 -179.445 ;
        RECT 18.405 -179.465 18.695 -178.740 ;
        RECT 20.235 -179.115 20.405 -178.590 ;
        RECT 20.235 -179.445 20.785 -179.115 ;
        RECT 18.320 -179.635 18.780 -179.465 ;
        RECT 20.235 -179.970 20.405 -179.445 ;
      LAYER mcon ;
        RECT -288.125 94.825 -287.955 94.995 ;
        RECT -286.355 94.725 -286.185 94.895 ;
        RECT -284.585 94.825 -284.415 94.995 ;
        RECT -288.125 94.365 -287.955 94.535 ;
        RECT -288.125 93.905 -287.955 94.075 ;
        RECT -278.205 94.825 -278.035 94.995 ;
        RECT -276.435 94.725 -276.265 94.895 ;
        RECT -274.665 94.825 -274.495 94.995 ;
        RECT -284.585 94.365 -284.415 94.535 ;
        RECT -278.205 94.365 -278.035 94.535 ;
        RECT -284.585 93.905 -284.415 94.075 ;
        RECT -278.205 93.905 -278.035 94.075 ;
        RECT -268.285 94.825 -268.115 94.995 ;
        RECT -266.515 94.725 -266.345 94.895 ;
        RECT -264.745 94.825 -264.575 94.995 ;
        RECT -274.665 94.365 -274.495 94.535 ;
        RECT -268.285 94.365 -268.115 94.535 ;
        RECT -274.665 93.905 -274.495 94.075 ;
        RECT -268.285 93.905 -268.115 94.075 ;
        RECT -258.365 94.825 -258.195 94.995 ;
        RECT -256.595 94.725 -256.425 94.895 ;
        RECT -254.825 94.825 -254.655 94.995 ;
        RECT -264.745 94.365 -264.575 94.535 ;
        RECT -258.365 94.365 -258.195 94.535 ;
        RECT -264.745 93.905 -264.575 94.075 ;
        RECT -258.365 93.905 -258.195 94.075 ;
        RECT -248.445 94.825 -248.275 94.995 ;
        RECT -246.675 94.725 -246.505 94.895 ;
        RECT -244.905 94.825 -244.735 94.995 ;
        RECT -254.825 94.365 -254.655 94.535 ;
        RECT -248.445 94.365 -248.275 94.535 ;
        RECT -254.825 93.905 -254.655 94.075 ;
        RECT -248.445 93.905 -248.275 94.075 ;
        RECT -238.525 94.825 -238.355 94.995 ;
        RECT -236.755 94.725 -236.585 94.895 ;
        RECT -234.985 94.825 -234.815 94.995 ;
        RECT -244.905 94.365 -244.735 94.535 ;
        RECT -238.525 94.365 -238.355 94.535 ;
        RECT -244.905 93.905 -244.735 94.075 ;
        RECT -238.525 93.905 -238.355 94.075 ;
        RECT -228.605 94.825 -228.435 94.995 ;
        RECT -226.835 94.725 -226.665 94.895 ;
        RECT -225.065 94.825 -224.895 94.995 ;
        RECT -234.985 94.365 -234.815 94.535 ;
        RECT -228.605 94.365 -228.435 94.535 ;
        RECT -234.985 93.905 -234.815 94.075 ;
        RECT -228.605 93.905 -228.435 94.075 ;
        RECT -218.685 94.825 -218.515 94.995 ;
        RECT -216.915 94.725 -216.745 94.895 ;
        RECT -215.145 94.825 -214.975 94.995 ;
        RECT -225.065 94.365 -224.895 94.535 ;
        RECT -218.685 94.365 -218.515 94.535 ;
        RECT -225.065 93.905 -224.895 94.075 ;
        RECT -218.685 93.905 -218.515 94.075 ;
        RECT -208.765 94.825 -208.595 94.995 ;
        RECT -206.995 94.725 -206.825 94.895 ;
        RECT -205.225 94.825 -205.055 94.995 ;
        RECT -215.145 94.365 -214.975 94.535 ;
        RECT -208.765 94.365 -208.595 94.535 ;
        RECT -215.145 93.905 -214.975 94.075 ;
        RECT -208.765 93.905 -208.595 94.075 ;
        RECT -198.845 94.825 -198.675 94.995 ;
        RECT -197.075 94.725 -196.905 94.895 ;
        RECT -195.305 94.825 -195.135 94.995 ;
        RECT -205.225 94.365 -205.055 94.535 ;
        RECT -198.845 94.365 -198.675 94.535 ;
        RECT -205.225 93.905 -205.055 94.075 ;
        RECT -198.845 93.905 -198.675 94.075 ;
        RECT -188.925 94.825 -188.755 94.995 ;
        RECT -187.155 94.725 -186.985 94.895 ;
        RECT -185.385 94.825 -185.215 94.995 ;
        RECT -195.305 94.365 -195.135 94.535 ;
        RECT -188.925 94.365 -188.755 94.535 ;
        RECT -195.305 93.905 -195.135 94.075 ;
        RECT -188.925 93.905 -188.755 94.075 ;
        RECT -179.005 94.825 -178.835 94.995 ;
        RECT -177.235 94.725 -177.065 94.895 ;
        RECT -175.465 94.825 -175.295 94.995 ;
        RECT -185.385 94.365 -185.215 94.535 ;
        RECT -179.005 94.365 -178.835 94.535 ;
        RECT -185.385 93.905 -185.215 94.075 ;
        RECT -179.005 93.905 -178.835 94.075 ;
        RECT -169.085 94.825 -168.915 94.995 ;
        RECT -167.315 94.725 -167.145 94.895 ;
        RECT -165.545 94.825 -165.375 94.995 ;
        RECT -175.465 94.365 -175.295 94.535 ;
        RECT -169.085 94.365 -168.915 94.535 ;
        RECT -175.465 93.905 -175.295 94.075 ;
        RECT -169.085 93.905 -168.915 94.075 ;
        RECT -159.165 94.825 -158.995 94.995 ;
        RECT -157.395 94.725 -157.225 94.895 ;
        RECT -155.625 94.825 -155.455 94.995 ;
        RECT -165.545 94.365 -165.375 94.535 ;
        RECT -159.165 94.365 -158.995 94.535 ;
        RECT -165.545 93.905 -165.375 94.075 ;
        RECT -159.165 93.905 -158.995 94.075 ;
        RECT -149.245 94.825 -149.075 94.995 ;
        RECT -147.475 94.725 -147.305 94.895 ;
        RECT -145.705 94.825 -145.535 94.995 ;
        RECT -155.625 94.365 -155.455 94.535 ;
        RECT -149.245 94.365 -149.075 94.535 ;
        RECT -155.625 93.905 -155.455 94.075 ;
        RECT -149.245 93.905 -149.075 94.075 ;
        RECT -139.325 94.825 -139.155 94.995 ;
        RECT -137.555 94.725 -137.385 94.895 ;
        RECT -135.785 94.825 -135.615 94.995 ;
        RECT -145.705 94.365 -145.535 94.535 ;
        RECT -139.325 94.365 -139.155 94.535 ;
        RECT -145.705 93.905 -145.535 94.075 ;
        RECT -139.325 93.905 -139.155 94.075 ;
        RECT -129.405 94.825 -129.235 94.995 ;
        RECT -127.635 94.725 -127.465 94.895 ;
        RECT -125.865 94.825 -125.695 94.995 ;
        RECT -135.785 94.365 -135.615 94.535 ;
        RECT -129.405 94.365 -129.235 94.535 ;
        RECT -135.785 93.905 -135.615 94.075 ;
        RECT -129.405 93.905 -129.235 94.075 ;
        RECT -119.485 94.825 -119.315 94.995 ;
        RECT -117.715 94.725 -117.545 94.895 ;
        RECT -115.945 94.825 -115.775 94.995 ;
        RECT -125.865 94.365 -125.695 94.535 ;
        RECT -119.485 94.365 -119.315 94.535 ;
        RECT -125.865 93.905 -125.695 94.075 ;
        RECT -119.485 93.905 -119.315 94.075 ;
        RECT -109.565 94.825 -109.395 94.995 ;
        RECT -107.795 94.725 -107.625 94.895 ;
        RECT -106.025 94.825 -105.855 94.995 ;
        RECT -115.945 94.365 -115.775 94.535 ;
        RECT -109.565 94.365 -109.395 94.535 ;
        RECT -115.945 93.905 -115.775 94.075 ;
        RECT -109.565 93.905 -109.395 94.075 ;
        RECT -99.645 94.825 -99.475 94.995 ;
        RECT -97.875 94.725 -97.705 94.895 ;
        RECT -96.105 94.825 -95.935 94.995 ;
        RECT -106.025 94.365 -105.855 94.535 ;
        RECT -99.645 94.365 -99.475 94.535 ;
        RECT -106.025 93.905 -105.855 94.075 ;
        RECT -99.645 93.905 -99.475 94.075 ;
        RECT -89.725 94.825 -89.555 94.995 ;
        RECT -87.955 94.725 -87.785 94.895 ;
        RECT -86.185 94.825 -86.015 94.995 ;
        RECT -96.105 94.365 -95.935 94.535 ;
        RECT -89.725 94.365 -89.555 94.535 ;
        RECT -96.105 93.905 -95.935 94.075 ;
        RECT -89.725 93.905 -89.555 94.075 ;
        RECT -79.805 94.825 -79.635 94.995 ;
        RECT -78.035 94.725 -77.865 94.895 ;
        RECT -76.265 94.825 -76.095 94.995 ;
        RECT -86.185 94.365 -86.015 94.535 ;
        RECT -79.805 94.365 -79.635 94.535 ;
        RECT -86.185 93.905 -86.015 94.075 ;
        RECT -79.805 93.905 -79.635 94.075 ;
        RECT -69.885 94.825 -69.715 94.995 ;
        RECT -68.115 94.725 -67.945 94.895 ;
        RECT -66.345 94.825 -66.175 94.995 ;
        RECT -76.265 94.365 -76.095 94.535 ;
        RECT -69.885 94.365 -69.715 94.535 ;
        RECT -76.265 93.905 -76.095 94.075 ;
        RECT -69.885 93.905 -69.715 94.075 ;
        RECT -59.965 94.825 -59.795 94.995 ;
        RECT -58.195 94.725 -58.025 94.895 ;
        RECT -56.425 94.825 -56.255 94.995 ;
        RECT -66.345 94.365 -66.175 94.535 ;
        RECT -59.965 94.365 -59.795 94.535 ;
        RECT -66.345 93.905 -66.175 94.075 ;
        RECT -59.965 93.905 -59.795 94.075 ;
        RECT -50.045 94.825 -49.875 94.995 ;
        RECT -48.275 94.725 -48.105 94.895 ;
        RECT -46.505 94.825 -46.335 94.995 ;
        RECT -56.425 94.365 -56.255 94.535 ;
        RECT -50.045 94.365 -49.875 94.535 ;
        RECT -56.425 93.905 -56.255 94.075 ;
        RECT -50.045 93.905 -49.875 94.075 ;
        RECT -40.125 94.825 -39.955 94.995 ;
        RECT -38.355 94.725 -38.185 94.895 ;
        RECT -36.585 94.825 -36.415 94.995 ;
        RECT -46.505 94.365 -46.335 94.535 ;
        RECT -40.125 94.365 -39.955 94.535 ;
        RECT -46.505 93.905 -46.335 94.075 ;
        RECT -40.125 93.905 -39.955 94.075 ;
        RECT -30.205 94.825 -30.035 94.995 ;
        RECT -28.435 94.725 -28.265 94.895 ;
        RECT -26.665 94.825 -26.495 94.995 ;
        RECT -36.585 94.365 -36.415 94.535 ;
        RECT -30.205 94.365 -30.035 94.535 ;
        RECT -36.585 93.905 -36.415 94.075 ;
        RECT -30.205 93.905 -30.035 94.075 ;
        RECT -20.285 94.825 -20.115 94.995 ;
        RECT -18.515 94.725 -18.345 94.895 ;
        RECT -16.745 94.825 -16.575 94.995 ;
        RECT -26.665 94.365 -26.495 94.535 ;
        RECT -20.285 94.365 -20.115 94.535 ;
        RECT -26.665 93.905 -26.495 94.075 ;
        RECT -20.285 93.905 -20.115 94.075 ;
        RECT -10.365 94.825 -10.195 94.995 ;
        RECT -8.595 94.725 -8.425 94.895 ;
        RECT -6.825 94.825 -6.655 94.995 ;
        RECT -16.745 94.365 -16.575 94.535 ;
        RECT -10.365 94.365 -10.195 94.535 ;
        RECT -16.745 93.905 -16.575 94.075 ;
        RECT -10.365 93.905 -10.195 94.075 ;
        RECT -0.445 94.825 -0.275 94.995 ;
        RECT 1.325 94.725 1.495 94.895 ;
        RECT 3.095 94.825 3.265 94.995 ;
        RECT -6.825 94.365 -6.655 94.535 ;
        RECT -0.445 94.365 -0.275 94.535 ;
        RECT -6.825 93.905 -6.655 94.075 ;
        RECT -0.445 93.905 -0.275 94.075 ;
        RECT 9.475 94.825 9.645 94.995 ;
        RECT 11.245 94.725 11.415 94.895 ;
        RECT 13.015 94.825 13.185 94.995 ;
        RECT 3.095 94.365 3.265 94.535 ;
        RECT 9.475 94.365 9.645 94.535 ;
        RECT 3.095 93.905 3.265 94.075 ;
        RECT 9.475 93.905 9.645 94.075 ;
        RECT 19.395 94.825 19.565 94.995 ;
        RECT 21.165 94.725 21.335 94.895 ;
        RECT 22.935 94.825 23.105 94.995 ;
        RECT 13.015 94.365 13.185 94.535 ;
        RECT 19.395 94.365 19.565 94.535 ;
        RECT 13.015 93.905 13.185 94.075 ;
        RECT 19.395 93.905 19.565 94.075 ;
        RECT 22.935 94.365 23.105 94.535 ;
        RECT 22.935 93.905 23.105 94.075 ;
        RECT -282.775 93.245 -282.605 93.415 ;
        RECT -282.315 93.245 -282.145 93.415 ;
        RECT -281.855 93.245 -281.685 93.415 ;
        RECT -281.395 93.245 -281.225 93.415 ;
        RECT -280.935 93.245 -280.765 93.415 ;
        RECT -280.475 93.245 -280.305 93.415 ;
        RECT -280.015 93.245 -279.845 93.415 ;
        RECT -272.855 93.245 -272.685 93.415 ;
        RECT -272.395 93.245 -272.225 93.415 ;
        RECT -271.935 93.245 -271.765 93.415 ;
        RECT -271.475 93.245 -271.305 93.415 ;
        RECT -271.015 93.245 -270.845 93.415 ;
        RECT -270.555 93.245 -270.385 93.415 ;
        RECT -270.095 93.245 -269.925 93.415 ;
        RECT -262.935 93.245 -262.765 93.415 ;
        RECT -262.475 93.245 -262.305 93.415 ;
        RECT -262.015 93.245 -261.845 93.415 ;
        RECT -261.555 93.245 -261.385 93.415 ;
        RECT -261.095 93.245 -260.925 93.415 ;
        RECT -260.635 93.245 -260.465 93.415 ;
        RECT -260.175 93.245 -260.005 93.415 ;
        RECT -253.015 93.245 -252.845 93.415 ;
        RECT -252.555 93.245 -252.385 93.415 ;
        RECT -252.095 93.245 -251.925 93.415 ;
        RECT -251.635 93.245 -251.465 93.415 ;
        RECT -251.175 93.245 -251.005 93.415 ;
        RECT -250.715 93.245 -250.545 93.415 ;
        RECT -250.255 93.245 -250.085 93.415 ;
        RECT -243.095 93.245 -242.925 93.415 ;
        RECT -242.635 93.245 -242.465 93.415 ;
        RECT -242.175 93.245 -242.005 93.415 ;
        RECT -241.715 93.245 -241.545 93.415 ;
        RECT -241.255 93.245 -241.085 93.415 ;
        RECT -240.795 93.245 -240.625 93.415 ;
        RECT -240.335 93.245 -240.165 93.415 ;
        RECT -233.175 93.245 -233.005 93.415 ;
        RECT -232.715 93.245 -232.545 93.415 ;
        RECT -232.255 93.245 -232.085 93.415 ;
        RECT -231.795 93.245 -231.625 93.415 ;
        RECT -231.335 93.245 -231.165 93.415 ;
        RECT -230.875 93.245 -230.705 93.415 ;
        RECT -230.415 93.245 -230.245 93.415 ;
        RECT -223.255 93.245 -223.085 93.415 ;
        RECT -222.795 93.245 -222.625 93.415 ;
        RECT -222.335 93.245 -222.165 93.415 ;
        RECT -221.875 93.245 -221.705 93.415 ;
        RECT -221.415 93.245 -221.245 93.415 ;
        RECT -220.955 93.245 -220.785 93.415 ;
        RECT -220.495 93.245 -220.325 93.415 ;
        RECT -213.335 93.245 -213.165 93.415 ;
        RECT -212.875 93.245 -212.705 93.415 ;
        RECT -212.415 93.245 -212.245 93.415 ;
        RECT -211.955 93.245 -211.785 93.415 ;
        RECT -211.495 93.245 -211.325 93.415 ;
        RECT -211.035 93.245 -210.865 93.415 ;
        RECT -210.575 93.245 -210.405 93.415 ;
        RECT -203.415 93.245 -203.245 93.415 ;
        RECT -202.955 93.245 -202.785 93.415 ;
        RECT -202.495 93.245 -202.325 93.415 ;
        RECT -202.035 93.245 -201.865 93.415 ;
        RECT -201.575 93.245 -201.405 93.415 ;
        RECT -201.115 93.245 -200.945 93.415 ;
        RECT -200.655 93.245 -200.485 93.415 ;
        RECT -193.495 93.245 -193.325 93.415 ;
        RECT -193.035 93.245 -192.865 93.415 ;
        RECT -192.575 93.245 -192.405 93.415 ;
        RECT -192.115 93.245 -191.945 93.415 ;
        RECT -191.655 93.245 -191.485 93.415 ;
        RECT -191.195 93.245 -191.025 93.415 ;
        RECT -190.735 93.245 -190.565 93.415 ;
        RECT -183.575 93.245 -183.405 93.415 ;
        RECT -183.115 93.245 -182.945 93.415 ;
        RECT -182.655 93.245 -182.485 93.415 ;
        RECT -182.195 93.245 -182.025 93.415 ;
        RECT -181.735 93.245 -181.565 93.415 ;
        RECT -181.275 93.245 -181.105 93.415 ;
        RECT -180.815 93.245 -180.645 93.415 ;
        RECT -173.655 93.245 -173.485 93.415 ;
        RECT -173.195 93.245 -173.025 93.415 ;
        RECT -172.735 93.245 -172.565 93.415 ;
        RECT -172.275 93.245 -172.105 93.415 ;
        RECT -171.815 93.245 -171.645 93.415 ;
        RECT -171.355 93.245 -171.185 93.415 ;
        RECT -170.895 93.245 -170.725 93.415 ;
        RECT -163.735 93.245 -163.565 93.415 ;
        RECT -163.275 93.245 -163.105 93.415 ;
        RECT -162.815 93.245 -162.645 93.415 ;
        RECT -162.355 93.245 -162.185 93.415 ;
        RECT -161.895 93.245 -161.725 93.415 ;
        RECT -161.435 93.245 -161.265 93.415 ;
        RECT -160.975 93.245 -160.805 93.415 ;
        RECT -153.815 93.245 -153.645 93.415 ;
        RECT -153.355 93.245 -153.185 93.415 ;
        RECT -152.895 93.245 -152.725 93.415 ;
        RECT -152.435 93.245 -152.265 93.415 ;
        RECT -151.975 93.245 -151.805 93.415 ;
        RECT -151.515 93.245 -151.345 93.415 ;
        RECT -151.055 93.245 -150.885 93.415 ;
        RECT -143.895 93.245 -143.725 93.415 ;
        RECT -143.435 93.245 -143.265 93.415 ;
        RECT -142.975 93.245 -142.805 93.415 ;
        RECT -142.515 93.245 -142.345 93.415 ;
        RECT -142.055 93.245 -141.885 93.415 ;
        RECT -141.595 93.245 -141.425 93.415 ;
        RECT -141.135 93.245 -140.965 93.415 ;
        RECT -133.975 93.245 -133.805 93.415 ;
        RECT -133.515 93.245 -133.345 93.415 ;
        RECT -133.055 93.245 -132.885 93.415 ;
        RECT -132.595 93.245 -132.425 93.415 ;
        RECT -132.135 93.245 -131.965 93.415 ;
        RECT -131.675 93.245 -131.505 93.415 ;
        RECT -131.215 93.245 -131.045 93.415 ;
        RECT -124.055 93.245 -123.885 93.415 ;
        RECT -123.595 93.245 -123.425 93.415 ;
        RECT -123.135 93.245 -122.965 93.415 ;
        RECT -122.675 93.245 -122.505 93.415 ;
        RECT -122.215 93.245 -122.045 93.415 ;
        RECT -121.755 93.245 -121.585 93.415 ;
        RECT -121.295 93.245 -121.125 93.415 ;
        RECT -114.135 93.245 -113.965 93.415 ;
        RECT -113.675 93.245 -113.505 93.415 ;
        RECT -113.215 93.245 -113.045 93.415 ;
        RECT -112.755 93.245 -112.585 93.415 ;
        RECT -112.295 93.245 -112.125 93.415 ;
        RECT -111.835 93.245 -111.665 93.415 ;
        RECT -111.375 93.245 -111.205 93.415 ;
        RECT -104.215 93.245 -104.045 93.415 ;
        RECT -103.755 93.245 -103.585 93.415 ;
        RECT -103.295 93.245 -103.125 93.415 ;
        RECT -102.835 93.245 -102.665 93.415 ;
        RECT -102.375 93.245 -102.205 93.415 ;
        RECT -101.915 93.245 -101.745 93.415 ;
        RECT -101.455 93.245 -101.285 93.415 ;
        RECT -94.295 93.245 -94.125 93.415 ;
        RECT -93.835 93.245 -93.665 93.415 ;
        RECT -93.375 93.245 -93.205 93.415 ;
        RECT -92.915 93.245 -92.745 93.415 ;
        RECT -92.455 93.245 -92.285 93.415 ;
        RECT -91.995 93.245 -91.825 93.415 ;
        RECT -91.535 93.245 -91.365 93.415 ;
        RECT -84.375 93.245 -84.205 93.415 ;
        RECT -83.915 93.245 -83.745 93.415 ;
        RECT -83.455 93.245 -83.285 93.415 ;
        RECT -82.995 93.245 -82.825 93.415 ;
        RECT -82.535 93.245 -82.365 93.415 ;
        RECT -82.075 93.245 -81.905 93.415 ;
        RECT -81.615 93.245 -81.445 93.415 ;
        RECT -74.455 93.245 -74.285 93.415 ;
        RECT -73.995 93.245 -73.825 93.415 ;
        RECT -73.535 93.245 -73.365 93.415 ;
        RECT -73.075 93.245 -72.905 93.415 ;
        RECT -72.615 93.245 -72.445 93.415 ;
        RECT -72.155 93.245 -71.985 93.415 ;
        RECT -71.695 93.245 -71.525 93.415 ;
        RECT -64.535 93.245 -64.365 93.415 ;
        RECT -64.075 93.245 -63.905 93.415 ;
        RECT -63.615 93.245 -63.445 93.415 ;
        RECT -63.155 93.245 -62.985 93.415 ;
        RECT -62.695 93.245 -62.525 93.415 ;
        RECT -62.235 93.245 -62.065 93.415 ;
        RECT -61.775 93.245 -61.605 93.415 ;
        RECT -54.615 93.245 -54.445 93.415 ;
        RECT -54.155 93.245 -53.985 93.415 ;
        RECT -53.695 93.245 -53.525 93.415 ;
        RECT -53.235 93.245 -53.065 93.415 ;
        RECT -52.775 93.245 -52.605 93.415 ;
        RECT -52.315 93.245 -52.145 93.415 ;
        RECT -51.855 93.245 -51.685 93.415 ;
        RECT -44.695 93.245 -44.525 93.415 ;
        RECT -44.235 93.245 -44.065 93.415 ;
        RECT -43.775 93.245 -43.605 93.415 ;
        RECT -43.315 93.245 -43.145 93.415 ;
        RECT -42.855 93.245 -42.685 93.415 ;
        RECT -42.395 93.245 -42.225 93.415 ;
        RECT -41.935 93.245 -41.765 93.415 ;
        RECT -34.775 93.245 -34.605 93.415 ;
        RECT -34.315 93.245 -34.145 93.415 ;
        RECT -33.855 93.245 -33.685 93.415 ;
        RECT -33.395 93.245 -33.225 93.415 ;
        RECT -32.935 93.245 -32.765 93.415 ;
        RECT -32.475 93.245 -32.305 93.415 ;
        RECT -32.015 93.245 -31.845 93.415 ;
        RECT -24.855 93.245 -24.685 93.415 ;
        RECT -24.395 93.245 -24.225 93.415 ;
        RECT -23.935 93.245 -23.765 93.415 ;
        RECT -23.475 93.245 -23.305 93.415 ;
        RECT -23.015 93.245 -22.845 93.415 ;
        RECT -22.555 93.245 -22.385 93.415 ;
        RECT -22.095 93.245 -21.925 93.415 ;
        RECT -14.935 93.245 -14.765 93.415 ;
        RECT -14.475 93.245 -14.305 93.415 ;
        RECT -14.015 93.245 -13.845 93.415 ;
        RECT -13.555 93.245 -13.385 93.415 ;
        RECT -13.095 93.245 -12.925 93.415 ;
        RECT -12.635 93.245 -12.465 93.415 ;
        RECT -12.175 93.245 -12.005 93.415 ;
        RECT -5.015 93.245 -4.845 93.415 ;
        RECT -4.555 93.245 -4.385 93.415 ;
        RECT -4.095 93.245 -3.925 93.415 ;
        RECT -3.635 93.245 -3.465 93.415 ;
        RECT -3.175 93.245 -3.005 93.415 ;
        RECT -2.715 93.245 -2.545 93.415 ;
        RECT -2.255 93.245 -2.085 93.415 ;
        RECT 4.905 93.245 5.075 93.415 ;
        RECT 5.365 93.245 5.535 93.415 ;
        RECT 5.825 93.245 5.995 93.415 ;
        RECT 6.285 93.245 6.455 93.415 ;
        RECT 6.745 93.245 6.915 93.415 ;
        RECT 7.205 93.245 7.375 93.415 ;
        RECT 7.665 93.245 7.835 93.415 ;
        RECT 14.825 93.245 14.995 93.415 ;
        RECT 15.285 93.245 15.455 93.415 ;
        RECT 15.745 93.245 15.915 93.415 ;
        RECT 16.205 93.245 16.375 93.415 ;
        RECT 16.665 93.245 16.835 93.415 ;
        RECT 17.125 93.245 17.295 93.415 ;
        RECT 17.585 93.245 17.755 93.415 ;
        RECT -287.735 90.525 -287.565 90.695 ;
        RECT -287.275 90.525 -287.105 90.695 ;
        RECT -286.815 90.525 -286.645 90.695 ;
        RECT -286.355 90.525 -286.185 90.695 ;
        RECT -285.895 90.525 -285.725 90.695 ;
        RECT -285.435 90.525 -285.265 90.695 ;
        RECT -284.975 90.525 -284.805 90.695 ;
        RECT -277.815 90.525 -277.645 90.695 ;
        RECT -277.355 90.525 -277.185 90.695 ;
        RECT -276.895 90.525 -276.725 90.695 ;
        RECT -276.435 90.525 -276.265 90.695 ;
        RECT -275.975 90.525 -275.805 90.695 ;
        RECT -275.515 90.525 -275.345 90.695 ;
        RECT -275.055 90.525 -274.885 90.695 ;
        RECT -267.895 90.525 -267.725 90.695 ;
        RECT -267.435 90.525 -267.265 90.695 ;
        RECT -266.975 90.525 -266.805 90.695 ;
        RECT -266.515 90.525 -266.345 90.695 ;
        RECT -266.055 90.525 -265.885 90.695 ;
        RECT -265.595 90.525 -265.425 90.695 ;
        RECT -265.135 90.525 -264.965 90.695 ;
        RECT -257.975 90.525 -257.805 90.695 ;
        RECT -257.515 90.525 -257.345 90.695 ;
        RECT -257.055 90.525 -256.885 90.695 ;
        RECT -256.595 90.525 -256.425 90.695 ;
        RECT -256.135 90.525 -255.965 90.695 ;
        RECT -255.675 90.525 -255.505 90.695 ;
        RECT -255.215 90.525 -255.045 90.695 ;
        RECT -248.055 90.525 -247.885 90.695 ;
        RECT -247.595 90.525 -247.425 90.695 ;
        RECT -247.135 90.525 -246.965 90.695 ;
        RECT -246.675 90.525 -246.505 90.695 ;
        RECT -246.215 90.525 -246.045 90.695 ;
        RECT -245.755 90.525 -245.585 90.695 ;
        RECT -245.295 90.525 -245.125 90.695 ;
        RECT -238.135 90.525 -237.965 90.695 ;
        RECT -237.675 90.525 -237.505 90.695 ;
        RECT -237.215 90.525 -237.045 90.695 ;
        RECT -236.755 90.525 -236.585 90.695 ;
        RECT -236.295 90.525 -236.125 90.695 ;
        RECT -235.835 90.525 -235.665 90.695 ;
        RECT -235.375 90.525 -235.205 90.695 ;
        RECT -228.215 90.525 -228.045 90.695 ;
        RECT -227.755 90.525 -227.585 90.695 ;
        RECT -227.295 90.525 -227.125 90.695 ;
        RECT -226.835 90.525 -226.665 90.695 ;
        RECT -226.375 90.525 -226.205 90.695 ;
        RECT -225.915 90.525 -225.745 90.695 ;
        RECT -225.455 90.525 -225.285 90.695 ;
        RECT -218.295 90.525 -218.125 90.695 ;
        RECT -217.835 90.525 -217.665 90.695 ;
        RECT -217.375 90.525 -217.205 90.695 ;
        RECT -216.915 90.525 -216.745 90.695 ;
        RECT -216.455 90.525 -216.285 90.695 ;
        RECT -215.995 90.525 -215.825 90.695 ;
        RECT -215.535 90.525 -215.365 90.695 ;
        RECT -208.375 90.525 -208.205 90.695 ;
        RECT -207.915 90.525 -207.745 90.695 ;
        RECT -207.455 90.525 -207.285 90.695 ;
        RECT -206.995 90.525 -206.825 90.695 ;
        RECT -206.535 90.525 -206.365 90.695 ;
        RECT -206.075 90.525 -205.905 90.695 ;
        RECT -205.615 90.525 -205.445 90.695 ;
        RECT -198.455 90.525 -198.285 90.695 ;
        RECT -197.995 90.525 -197.825 90.695 ;
        RECT -197.535 90.525 -197.365 90.695 ;
        RECT -197.075 90.525 -196.905 90.695 ;
        RECT -196.615 90.525 -196.445 90.695 ;
        RECT -196.155 90.525 -195.985 90.695 ;
        RECT -195.695 90.525 -195.525 90.695 ;
        RECT -188.535 90.525 -188.365 90.695 ;
        RECT -188.075 90.525 -187.905 90.695 ;
        RECT -187.615 90.525 -187.445 90.695 ;
        RECT -187.155 90.525 -186.985 90.695 ;
        RECT -186.695 90.525 -186.525 90.695 ;
        RECT -186.235 90.525 -186.065 90.695 ;
        RECT -185.775 90.525 -185.605 90.695 ;
        RECT -178.615 90.525 -178.445 90.695 ;
        RECT -178.155 90.525 -177.985 90.695 ;
        RECT -177.695 90.525 -177.525 90.695 ;
        RECT -177.235 90.525 -177.065 90.695 ;
        RECT -176.775 90.525 -176.605 90.695 ;
        RECT -176.315 90.525 -176.145 90.695 ;
        RECT -175.855 90.525 -175.685 90.695 ;
        RECT -168.695 90.525 -168.525 90.695 ;
        RECT -168.235 90.525 -168.065 90.695 ;
        RECT -167.775 90.525 -167.605 90.695 ;
        RECT -167.315 90.525 -167.145 90.695 ;
        RECT -166.855 90.525 -166.685 90.695 ;
        RECT -166.395 90.525 -166.225 90.695 ;
        RECT -165.935 90.525 -165.765 90.695 ;
        RECT -158.775 90.525 -158.605 90.695 ;
        RECT -158.315 90.525 -158.145 90.695 ;
        RECT -157.855 90.525 -157.685 90.695 ;
        RECT -157.395 90.525 -157.225 90.695 ;
        RECT -156.935 90.525 -156.765 90.695 ;
        RECT -156.475 90.525 -156.305 90.695 ;
        RECT -156.015 90.525 -155.845 90.695 ;
        RECT -148.855 90.525 -148.685 90.695 ;
        RECT -148.395 90.525 -148.225 90.695 ;
        RECT -147.935 90.525 -147.765 90.695 ;
        RECT -147.475 90.525 -147.305 90.695 ;
        RECT -147.015 90.525 -146.845 90.695 ;
        RECT -146.555 90.525 -146.385 90.695 ;
        RECT -146.095 90.525 -145.925 90.695 ;
        RECT -138.935 90.525 -138.765 90.695 ;
        RECT -138.475 90.525 -138.305 90.695 ;
        RECT -138.015 90.525 -137.845 90.695 ;
        RECT -137.555 90.525 -137.385 90.695 ;
        RECT -137.095 90.525 -136.925 90.695 ;
        RECT -136.635 90.525 -136.465 90.695 ;
        RECT -136.175 90.525 -136.005 90.695 ;
        RECT -129.015 90.525 -128.845 90.695 ;
        RECT -128.555 90.525 -128.385 90.695 ;
        RECT -128.095 90.525 -127.925 90.695 ;
        RECT -127.635 90.525 -127.465 90.695 ;
        RECT -127.175 90.525 -127.005 90.695 ;
        RECT -126.715 90.525 -126.545 90.695 ;
        RECT -126.255 90.525 -126.085 90.695 ;
        RECT -119.095 90.525 -118.925 90.695 ;
        RECT -118.635 90.525 -118.465 90.695 ;
        RECT -118.175 90.525 -118.005 90.695 ;
        RECT -117.715 90.525 -117.545 90.695 ;
        RECT -117.255 90.525 -117.085 90.695 ;
        RECT -116.795 90.525 -116.625 90.695 ;
        RECT -116.335 90.525 -116.165 90.695 ;
        RECT -109.175 90.525 -109.005 90.695 ;
        RECT -108.715 90.525 -108.545 90.695 ;
        RECT -108.255 90.525 -108.085 90.695 ;
        RECT -107.795 90.525 -107.625 90.695 ;
        RECT -107.335 90.525 -107.165 90.695 ;
        RECT -106.875 90.525 -106.705 90.695 ;
        RECT -106.415 90.525 -106.245 90.695 ;
        RECT -99.255 90.525 -99.085 90.695 ;
        RECT -98.795 90.525 -98.625 90.695 ;
        RECT -98.335 90.525 -98.165 90.695 ;
        RECT -97.875 90.525 -97.705 90.695 ;
        RECT -97.415 90.525 -97.245 90.695 ;
        RECT -96.955 90.525 -96.785 90.695 ;
        RECT -96.495 90.525 -96.325 90.695 ;
        RECT -89.335 90.525 -89.165 90.695 ;
        RECT -88.875 90.525 -88.705 90.695 ;
        RECT -88.415 90.525 -88.245 90.695 ;
        RECT -87.955 90.525 -87.785 90.695 ;
        RECT -87.495 90.525 -87.325 90.695 ;
        RECT -87.035 90.525 -86.865 90.695 ;
        RECT -86.575 90.525 -86.405 90.695 ;
        RECT -79.415 90.525 -79.245 90.695 ;
        RECT -78.955 90.525 -78.785 90.695 ;
        RECT -78.495 90.525 -78.325 90.695 ;
        RECT -78.035 90.525 -77.865 90.695 ;
        RECT -77.575 90.525 -77.405 90.695 ;
        RECT -77.115 90.525 -76.945 90.695 ;
        RECT -76.655 90.525 -76.485 90.695 ;
        RECT -69.495 90.525 -69.325 90.695 ;
        RECT -69.035 90.525 -68.865 90.695 ;
        RECT -68.575 90.525 -68.405 90.695 ;
        RECT -68.115 90.525 -67.945 90.695 ;
        RECT -67.655 90.525 -67.485 90.695 ;
        RECT -67.195 90.525 -67.025 90.695 ;
        RECT -66.735 90.525 -66.565 90.695 ;
        RECT -59.575 90.525 -59.405 90.695 ;
        RECT -59.115 90.525 -58.945 90.695 ;
        RECT -58.655 90.525 -58.485 90.695 ;
        RECT -58.195 90.525 -58.025 90.695 ;
        RECT -57.735 90.525 -57.565 90.695 ;
        RECT -57.275 90.525 -57.105 90.695 ;
        RECT -56.815 90.525 -56.645 90.695 ;
        RECT -49.655 90.525 -49.485 90.695 ;
        RECT -49.195 90.525 -49.025 90.695 ;
        RECT -48.735 90.525 -48.565 90.695 ;
        RECT -48.275 90.525 -48.105 90.695 ;
        RECT -47.815 90.525 -47.645 90.695 ;
        RECT -47.355 90.525 -47.185 90.695 ;
        RECT -46.895 90.525 -46.725 90.695 ;
        RECT -39.735 90.525 -39.565 90.695 ;
        RECT -39.275 90.525 -39.105 90.695 ;
        RECT -38.815 90.525 -38.645 90.695 ;
        RECT -38.355 90.525 -38.185 90.695 ;
        RECT -37.895 90.525 -37.725 90.695 ;
        RECT -37.435 90.525 -37.265 90.695 ;
        RECT -36.975 90.525 -36.805 90.695 ;
        RECT -29.815 90.525 -29.645 90.695 ;
        RECT -29.355 90.525 -29.185 90.695 ;
        RECT -28.895 90.525 -28.725 90.695 ;
        RECT -28.435 90.525 -28.265 90.695 ;
        RECT -27.975 90.525 -27.805 90.695 ;
        RECT -27.515 90.525 -27.345 90.695 ;
        RECT -27.055 90.525 -26.885 90.695 ;
        RECT -19.895 90.525 -19.725 90.695 ;
        RECT -19.435 90.525 -19.265 90.695 ;
        RECT -18.975 90.525 -18.805 90.695 ;
        RECT -18.515 90.525 -18.345 90.695 ;
        RECT -18.055 90.525 -17.885 90.695 ;
        RECT -17.595 90.525 -17.425 90.695 ;
        RECT -17.135 90.525 -16.965 90.695 ;
        RECT -9.975 90.525 -9.805 90.695 ;
        RECT -9.515 90.525 -9.345 90.695 ;
        RECT -9.055 90.525 -8.885 90.695 ;
        RECT -8.595 90.525 -8.425 90.695 ;
        RECT -8.135 90.525 -7.965 90.695 ;
        RECT -7.675 90.525 -7.505 90.695 ;
        RECT -7.215 90.525 -7.045 90.695 ;
        RECT -0.055 90.525 0.115 90.695 ;
        RECT 0.405 90.525 0.575 90.695 ;
        RECT 0.865 90.525 1.035 90.695 ;
        RECT 1.325 90.525 1.495 90.695 ;
        RECT 1.785 90.525 1.955 90.695 ;
        RECT 2.245 90.525 2.415 90.695 ;
        RECT 2.705 90.525 2.875 90.695 ;
        RECT 9.865 90.525 10.035 90.695 ;
        RECT 10.325 90.525 10.495 90.695 ;
        RECT 10.785 90.525 10.955 90.695 ;
        RECT 11.245 90.525 11.415 90.695 ;
        RECT 11.705 90.525 11.875 90.695 ;
        RECT 12.165 90.525 12.335 90.695 ;
        RECT 12.625 90.525 12.795 90.695 ;
        RECT 19.785 90.525 19.955 90.695 ;
        RECT 20.245 90.525 20.415 90.695 ;
        RECT 20.705 90.525 20.875 90.695 ;
        RECT 21.165 90.525 21.335 90.695 ;
        RECT 21.625 90.525 21.795 90.695 ;
        RECT 22.085 90.525 22.255 90.695 ;
        RECT 22.545 90.525 22.715 90.695 ;
        RECT -283.165 89.865 -282.995 90.035 ;
        RECT -283.165 89.405 -282.995 89.575 ;
        RECT -279.625 89.865 -279.455 90.035 ;
        RECT -273.245 89.865 -273.075 90.035 ;
        RECT -279.625 89.405 -279.455 89.575 ;
        RECT -273.245 89.405 -273.075 89.575 ;
        RECT -281.395 89.135 -281.225 89.305 ;
        RECT -283.165 88.945 -282.995 89.115 ;
        RECT -279.625 88.945 -279.455 89.115 ;
        RECT -269.705 89.865 -269.535 90.035 ;
        RECT -263.325 89.865 -263.155 90.035 ;
        RECT -269.705 89.405 -269.535 89.575 ;
        RECT -263.325 89.405 -263.155 89.575 ;
        RECT -271.475 89.135 -271.305 89.305 ;
        RECT -273.245 88.945 -273.075 89.115 ;
        RECT -269.705 88.945 -269.535 89.115 ;
        RECT -259.785 89.865 -259.615 90.035 ;
        RECT -253.405 89.865 -253.235 90.035 ;
        RECT -259.785 89.405 -259.615 89.575 ;
        RECT -253.405 89.405 -253.235 89.575 ;
        RECT -261.555 89.135 -261.385 89.305 ;
        RECT -263.325 88.945 -263.155 89.115 ;
        RECT -259.785 88.945 -259.615 89.115 ;
        RECT -249.865 89.865 -249.695 90.035 ;
        RECT -243.485 89.865 -243.315 90.035 ;
        RECT -249.865 89.405 -249.695 89.575 ;
        RECT -243.485 89.405 -243.315 89.575 ;
        RECT -251.635 89.135 -251.465 89.305 ;
        RECT -253.405 88.945 -253.235 89.115 ;
        RECT -249.865 88.945 -249.695 89.115 ;
        RECT -239.945 89.865 -239.775 90.035 ;
        RECT -233.565 89.865 -233.395 90.035 ;
        RECT -239.945 89.405 -239.775 89.575 ;
        RECT -233.565 89.405 -233.395 89.575 ;
        RECT -241.715 89.135 -241.545 89.305 ;
        RECT -243.485 88.945 -243.315 89.115 ;
        RECT -239.945 88.945 -239.775 89.115 ;
        RECT -230.025 89.865 -229.855 90.035 ;
        RECT -223.645 89.865 -223.475 90.035 ;
        RECT -230.025 89.405 -229.855 89.575 ;
        RECT -223.645 89.405 -223.475 89.575 ;
        RECT -231.795 89.135 -231.625 89.305 ;
        RECT -233.565 88.945 -233.395 89.115 ;
        RECT -230.025 88.945 -229.855 89.115 ;
        RECT -220.105 89.865 -219.935 90.035 ;
        RECT -213.725 89.865 -213.555 90.035 ;
        RECT -220.105 89.405 -219.935 89.575 ;
        RECT -213.725 89.405 -213.555 89.575 ;
        RECT -221.875 89.135 -221.705 89.305 ;
        RECT -223.645 88.945 -223.475 89.115 ;
        RECT -220.105 88.945 -219.935 89.115 ;
        RECT -210.185 89.865 -210.015 90.035 ;
        RECT -203.805 89.865 -203.635 90.035 ;
        RECT -210.185 89.405 -210.015 89.575 ;
        RECT -203.805 89.405 -203.635 89.575 ;
        RECT -211.955 89.135 -211.785 89.305 ;
        RECT -213.725 88.945 -213.555 89.115 ;
        RECT -210.185 88.945 -210.015 89.115 ;
        RECT -200.265 89.865 -200.095 90.035 ;
        RECT -193.885 89.865 -193.715 90.035 ;
        RECT -200.265 89.405 -200.095 89.575 ;
        RECT -193.885 89.405 -193.715 89.575 ;
        RECT -202.035 89.135 -201.865 89.305 ;
        RECT -203.805 88.945 -203.635 89.115 ;
        RECT -200.265 88.945 -200.095 89.115 ;
        RECT -190.345 89.865 -190.175 90.035 ;
        RECT -183.965 89.865 -183.795 90.035 ;
        RECT -190.345 89.405 -190.175 89.575 ;
        RECT -183.965 89.405 -183.795 89.575 ;
        RECT -192.115 89.135 -191.945 89.305 ;
        RECT -193.885 88.945 -193.715 89.115 ;
        RECT -190.345 88.945 -190.175 89.115 ;
        RECT -180.425 89.865 -180.255 90.035 ;
        RECT -174.045 89.865 -173.875 90.035 ;
        RECT -180.425 89.405 -180.255 89.575 ;
        RECT -174.045 89.405 -173.875 89.575 ;
        RECT -182.195 89.135 -182.025 89.305 ;
        RECT -183.965 88.945 -183.795 89.115 ;
        RECT -180.425 88.945 -180.255 89.115 ;
        RECT -170.505 89.865 -170.335 90.035 ;
        RECT -164.125 89.865 -163.955 90.035 ;
        RECT -170.505 89.405 -170.335 89.575 ;
        RECT -164.125 89.405 -163.955 89.575 ;
        RECT -172.275 89.135 -172.105 89.305 ;
        RECT -174.045 88.945 -173.875 89.115 ;
        RECT -170.505 88.945 -170.335 89.115 ;
        RECT -160.585 89.865 -160.415 90.035 ;
        RECT -154.205 89.865 -154.035 90.035 ;
        RECT -160.585 89.405 -160.415 89.575 ;
        RECT -154.205 89.405 -154.035 89.575 ;
        RECT -162.355 89.135 -162.185 89.305 ;
        RECT -164.125 88.945 -163.955 89.115 ;
        RECT -160.585 88.945 -160.415 89.115 ;
        RECT -150.665 89.865 -150.495 90.035 ;
        RECT -144.285 89.865 -144.115 90.035 ;
        RECT -150.665 89.405 -150.495 89.575 ;
        RECT -144.285 89.405 -144.115 89.575 ;
        RECT -152.435 89.135 -152.265 89.305 ;
        RECT -154.205 88.945 -154.035 89.115 ;
        RECT -150.665 88.945 -150.495 89.115 ;
        RECT -140.745 89.865 -140.575 90.035 ;
        RECT -134.365 89.865 -134.195 90.035 ;
        RECT -140.745 89.405 -140.575 89.575 ;
        RECT -134.365 89.405 -134.195 89.575 ;
        RECT -142.515 89.135 -142.345 89.305 ;
        RECT -144.285 88.945 -144.115 89.115 ;
        RECT -140.745 88.945 -140.575 89.115 ;
        RECT -130.825 89.865 -130.655 90.035 ;
        RECT -124.445 89.865 -124.275 90.035 ;
        RECT -130.825 89.405 -130.655 89.575 ;
        RECT -124.445 89.405 -124.275 89.575 ;
        RECT -132.595 89.135 -132.425 89.305 ;
        RECT -134.365 88.945 -134.195 89.115 ;
        RECT -130.825 88.945 -130.655 89.115 ;
        RECT -120.905 89.865 -120.735 90.035 ;
        RECT -114.525 89.865 -114.355 90.035 ;
        RECT -120.905 89.405 -120.735 89.575 ;
        RECT -114.525 89.405 -114.355 89.575 ;
        RECT -122.675 89.135 -122.505 89.305 ;
        RECT -124.445 88.945 -124.275 89.115 ;
        RECT -120.905 88.945 -120.735 89.115 ;
        RECT -110.985 89.865 -110.815 90.035 ;
        RECT -104.605 89.865 -104.435 90.035 ;
        RECT -110.985 89.405 -110.815 89.575 ;
        RECT -104.605 89.405 -104.435 89.575 ;
        RECT -112.755 89.135 -112.585 89.305 ;
        RECT -114.525 88.945 -114.355 89.115 ;
        RECT -110.985 88.945 -110.815 89.115 ;
        RECT -101.065 89.865 -100.895 90.035 ;
        RECT -94.685 89.865 -94.515 90.035 ;
        RECT -101.065 89.405 -100.895 89.575 ;
        RECT -94.685 89.405 -94.515 89.575 ;
        RECT -102.835 89.135 -102.665 89.305 ;
        RECT -104.605 88.945 -104.435 89.115 ;
        RECT -101.065 88.945 -100.895 89.115 ;
        RECT -91.145 89.865 -90.975 90.035 ;
        RECT -84.765 89.865 -84.595 90.035 ;
        RECT -91.145 89.405 -90.975 89.575 ;
        RECT -84.765 89.405 -84.595 89.575 ;
        RECT -92.915 89.135 -92.745 89.305 ;
        RECT -94.685 88.945 -94.515 89.115 ;
        RECT -91.145 88.945 -90.975 89.115 ;
        RECT -81.225 89.865 -81.055 90.035 ;
        RECT -74.845 89.865 -74.675 90.035 ;
        RECT -81.225 89.405 -81.055 89.575 ;
        RECT -74.845 89.405 -74.675 89.575 ;
        RECT -82.995 89.135 -82.825 89.305 ;
        RECT -84.765 88.945 -84.595 89.115 ;
        RECT -81.225 88.945 -81.055 89.115 ;
        RECT -71.305 89.865 -71.135 90.035 ;
        RECT -64.925 89.865 -64.755 90.035 ;
        RECT -71.305 89.405 -71.135 89.575 ;
        RECT -64.925 89.405 -64.755 89.575 ;
        RECT -73.075 89.135 -72.905 89.305 ;
        RECT -74.845 88.945 -74.675 89.115 ;
        RECT -71.305 88.945 -71.135 89.115 ;
        RECT -61.385 89.865 -61.215 90.035 ;
        RECT -55.005 89.865 -54.835 90.035 ;
        RECT -61.385 89.405 -61.215 89.575 ;
        RECT -55.005 89.405 -54.835 89.575 ;
        RECT -63.155 89.135 -62.985 89.305 ;
        RECT -64.925 88.945 -64.755 89.115 ;
        RECT -61.385 88.945 -61.215 89.115 ;
        RECT -51.465 89.865 -51.295 90.035 ;
        RECT -45.085 89.865 -44.915 90.035 ;
        RECT -51.465 89.405 -51.295 89.575 ;
        RECT -45.085 89.405 -44.915 89.575 ;
        RECT -53.235 89.135 -53.065 89.305 ;
        RECT -55.005 88.945 -54.835 89.115 ;
        RECT -51.465 88.945 -51.295 89.115 ;
        RECT -41.545 89.865 -41.375 90.035 ;
        RECT -35.165 89.865 -34.995 90.035 ;
        RECT -41.545 89.405 -41.375 89.575 ;
        RECT -35.165 89.405 -34.995 89.575 ;
        RECT -43.315 89.135 -43.145 89.305 ;
        RECT -45.085 88.945 -44.915 89.115 ;
        RECT -41.545 88.945 -41.375 89.115 ;
        RECT -31.625 89.865 -31.455 90.035 ;
        RECT -25.245 89.865 -25.075 90.035 ;
        RECT -31.625 89.405 -31.455 89.575 ;
        RECT -25.245 89.405 -25.075 89.575 ;
        RECT -33.395 89.135 -33.225 89.305 ;
        RECT -35.165 88.945 -34.995 89.115 ;
        RECT -31.625 88.945 -31.455 89.115 ;
        RECT -21.705 89.865 -21.535 90.035 ;
        RECT -15.325 89.865 -15.155 90.035 ;
        RECT -21.705 89.405 -21.535 89.575 ;
        RECT -15.325 89.405 -15.155 89.575 ;
        RECT -23.475 89.135 -23.305 89.305 ;
        RECT -25.245 88.945 -25.075 89.115 ;
        RECT -21.705 88.945 -21.535 89.115 ;
        RECT -11.785 89.865 -11.615 90.035 ;
        RECT -5.405 89.865 -5.235 90.035 ;
        RECT -11.785 89.405 -11.615 89.575 ;
        RECT -5.405 89.405 -5.235 89.575 ;
        RECT -13.555 89.135 -13.385 89.305 ;
        RECT -15.325 88.945 -15.155 89.115 ;
        RECT -11.785 88.945 -11.615 89.115 ;
        RECT -1.865 89.865 -1.695 90.035 ;
        RECT 4.515 89.865 4.685 90.035 ;
        RECT -1.865 89.405 -1.695 89.575 ;
        RECT 4.515 89.405 4.685 89.575 ;
        RECT -3.635 89.135 -3.465 89.305 ;
        RECT -5.405 88.945 -5.235 89.115 ;
        RECT -1.865 88.945 -1.695 89.115 ;
        RECT 8.055 89.865 8.225 90.035 ;
        RECT 14.435 89.865 14.605 90.035 ;
        RECT 8.055 89.405 8.225 89.575 ;
        RECT 14.435 89.405 14.605 89.575 ;
        RECT 6.285 89.135 6.455 89.305 ;
        RECT 4.515 88.945 4.685 89.115 ;
        RECT 8.055 88.945 8.225 89.115 ;
        RECT 17.975 89.865 18.145 90.035 ;
        RECT 17.975 89.405 18.145 89.575 ;
        RECT 16.205 89.135 16.375 89.305 ;
        RECT 14.435 88.945 14.605 89.115 ;
        RECT 17.975 88.945 18.145 89.115 ;
        RECT -287.875 7.115 -287.705 7.285 ;
        RECT -286.105 7.015 -285.935 7.185 ;
        RECT -284.335 7.115 -284.165 7.285 ;
        RECT -287.875 6.655 -287.705 6.825 ;
        RECT -287.875 6.195 -287.705 6.365 ;
        RECT -277.955 7.115 -277.785 7.285 ;
        RECT -276.185 7.015 -276.015 7.185 ;
        RECT -274.415 7.115 -274.245 7.285 ;
        RECT -284.335 6.655 -284.165 6.825 ;
        RECT -277.955 6.655 -277.785 6.825 ;
        RECT -284.335 6.195 -284.165 6.365 ;
        RECT -277.955 6.195 -277.785 6.365 ;
        RECT -268.035 7.115 -267.865 7.285 ;
        RECT -266.265 7.015 -266.095 7.185 ;
        RECT -264.495 7.115 -264.325 7.285 ;
        RECT -274.415 6.655 -274.245 6.825 ;
        RECT -268.035 6.655 -267.865 6.825 ;
        RECT -274.415 6.195 -274.245 6.365 ;
        RECT -268.035 6.195 -267.865 6.365 ;
        RECT -258.115 7.115 -257.945 7.285 ;
        RECT -256.345 7.015 -256.175 7.185 ;
        RECT -254.575 7.115 -254.405 7.285 ;
        RECT -264.495 6.655 -264.325 6.825 ;
        RECT -258.115 6.655 -257.945 6.825 ;
        RECT -264.495 6.195 -264.325 6.365 ;
        RECT -258.115 6.195 -257.945 6.365 ;
        RECT -248.195 7.115 -248.025 7.285 ;
        RECT -246.425 7.015 -246.255 7.185 ;
        RECT -244.655 7.115 -244.485 7.285 ;
        RECT -254.575 6.655 -254.405 6.825 ;
        RECT -248.195 6.655 -248.025 6.825 ;
        RECT -254.575 6.195 -254.405 6.365 ;
        RECT -248.195 6.195 -248.025 6.365 ;
        RECT -238.275 7.115 -238.105 7.285 ;
        RECT -236.505 7.015 -236.335 7.185 ;
        RECT -234.735 7.115 -234.565 7.285 ;
        RECT -244.655 6.655 -244.485 6.825 ;
        RECT -238.275 6.655 -238.105 6.825 ;
        RECT -244.655 6.195 -244.485 6.365 ;
        RECT -238.275 6.195 -238.105 6.365 ;
        RECT -228.355 7.115 -228.185 7.285 ;
        RECT -226.585 7.015 -226.415 7.185 ;
        RECT -224.815 7.115 -224.645 7.285 ;
        RECT -234.735 6.655 -234.565 6.825 ;
        RECT -228.355 6.655 -228.185 6.825 ;
        RECT -234.735 6.195 -234.565 6.365 ;
        RECT -228.355 6.195 -228.185 6.365 ;
        RECT -218.435 7.115 -218.265 7.285 ;
        RECT -216.665 7.015 -216.495 7.185 ;
        RECT -214.895 7.115 -214.725 7.285 ;
        RECT -224.815 6.655 -224.645 6.825 ;
        RECT -218.435 6.655 -218.265 6.825 ;
        RECT -224.815 6.195 -224.645 6.365 ;
        RECT -218.435 6.195 -218.265 6.365 ;
        RECT -208.515 7.115 -208.345 7.285 ;
        RECT -206.745 7.015 -206.575 7.185 ;
        RECT -204.975 7.115 -204.805 7.285 ;
        RECT -214.895 6.655 -214.725 6.825 ;
        RECT -208.515 6.655 -208.345 6.825 ;
        RECT -214.895 6.195 -214.725 6.365 ;
        RECT -208.515 6.195 -208.345 6.365 ;
        RECT -198.595 7.115 -198.425 7.285 ;
        RECT -196.825 7.015 -196.655 7.185 ;
        RECT -195.055 7.115 -194.885 7.285 ;
        RECT -204.975 6.655 -204.805 6.825 ;
        RECT -198.595 6.655 -198.425 6.825 ;
        RECT -204.975 6.195 -204.805 6.365 ;
        RECT -198.595 6.195 -198.425 6.365 ;
        RECT -188.675 7.115 -188.505 7.285 ;
        RECT -186.905 7.015 -186.735 7.185 ;
        RECT -185.135 7.115 -184.965 7.285 ;
        RECT -195.055 6.655 -194.885 6.825 ;
        RECT -188.675 6.655 -188.505 6.825 ;
        RECT -195.055 6.195 -194.885 6.365 ;
        RECT -188.675 6.195 -188.505 6.365 ;
        RECT -178.755 7.115 -178.585 7.285 ;
        RECT -176.985 7.015 -176.815 7.185 ;
        RECT -175.215 7.115 -175.045 7.285 ;
        RECT -185.135 6.655 -184.965 6.825 ;
        RECT -178.755 6.655 -178.585 6.825 ;
        RECT -185.135 6.195 -184.965 6.365 ;
        RECT -178.755 6.195 -178.585 6.365 ;
        RECT -168.835 7.115 -168.665 7.285 ;
        RECT -167.065 7.015 -166.895 7.185 ;
        RECT -165.295 7.115 -165.125 7.285 ;
        RECT -175.215 6.655 -175.045 6.825 ;
        RECT -168.835 6.655 -168.665 6.825 ;
        RECT -175.215 6.195 -175.045 6.365 ;
        RECT -168.835 6.195 -168.665 6.365 ;
        RECT -158.915 7.115 -158.745 7.285 ;
        RECT -157.145 7.015 -156.975 7.185 ;
        RECT -155.375 7.115 -155.205 7.285 ;
        RECT -165.295 6.655 -165.125 6.825 ;
        RECT -158.915 6.655 -158.745 6.825 ;
        RECT -165.295 6.195 -165.125 6.365 ;
        RECT -158.915 6.195 -158.745 6.365 ;
        RECT -148.995 7.115 -148.825 7.285 ;
        RECT -147.225 7.015 -147.055 7.185 ;
        RECT -145.455 7.115 -145.285 7.285 ;
        RECT -155.375 6.655 -155.205 6.825 ;
        RECT -148.995 6.655 -148.825 6.825 ;
        RECT -155.375 6.195 -155.205 6.365 ;
        RECT -148.995 6.195 -148.825 6.365 ;
        RECT -139.075 7.115 -138.905 7.285 ;
        RECT -137.305 7.015 -137.135 7.185 ;
        RECT -135.535 7.115 -135.365 7.285 ;
        RECT -145.455 6.655 -145.285 6.825 ;
        RECT -139.075 6.655 -138.905 6.825 ;
        RECT -145.455 6.195 -145.285 6.365 ;
        RECT -139.075 6.195 -138.905 6.365 ;
        RECT -129.155 7.115 -128.985 7.285 ;
        RECT -127.385 7.015 -127.215 7.185 ;
        RECT -125.615 7.115 -125.445 7.285 ;
        RECT -135.535 6.655 -135.365 6.825 ;
        RECT -129.155 6.655 -128.985 6.825 ;
        RECT -135.535 6.195 -135.365 6.365 ;
        RECT -129.155 6.195 -128.985 6.365 ;
        RECT -119.235 7.115 -119.065 7.285 ;
        RECT -117.465 7.015 -117.295 7.185 ;
        RECT -115.695 7.115 -115.525 7.285 ;
        RECT -125.615 6.655 -125.445 6.825 ;
        RECT -119.235 6.655 -119.065 6.825 ;
        RECT -125.615 6.195 -125.445 6.365 ;
        RECT -119.235 6.195 -119.065 6.365 ;
        RECT -109.315 7.115 -109.145 7.285 ;
        RECT -107.545 7.015 -107.375 7.185 ;
        RECT -105.775 7.115 -105.605 7.285 ;
        RECT -115.695 6.655 -115.525 6.825 ;
        RECT -109.315 6.655 -109.145 6.825 ;
        RECT -115.695 6.195 -115.525 6.365 ;
        RECT -109.315 6.195 -109.145 6.365 ;
        RECT -99.395 7.115 -99.225 7.285 ;
        RECT -97.625 7.015 -97.455 7.185 ;
        RECT -95.855 7.115 -95.685 7.285 ;
        RECT -105.775 6.655 -105.605 6.825 ;
        RECT -99.395 6.655 -99.225 6.825 ;
        RECT -105.775 6.195 -105.605 6.365 ;
        RECT -99.395 6.195 -99.225 6.365 ;
        RECT -89.475 7.115 -89.305 7.285 ;
        RECT -87.705 7.015 -87.535 7.185 ;
        RECT -85.935 7.115 -85.765 7.285 ;
        RECT -95.855 6.655 -95.685 6.825 ;
        RECT -89.475 6.655 -89.305 6.825 ;
        RECT -95.855 6.195 -95.685 6.365 ;
        RECT -89.475 6.195 -89.305 6.365 ;
        RECT -79.555 7.115 -79.385 7.285 ;
        RECT -77.785 7.015 -77.615 7.185 ;
        RECT -76.015 7.115 -75.845 7.285 ;
        RECT -85.935 6.655 -85.765 6.825 ;
        RECT -79.555 6.655 -79.385 6.825 ;
        RECT -85.935 6.195 -85.765 6.365 ;
        RECT -79.555 6.195 -79.385 6.365 ;
        RECT -69.635 7.115 -69.465 7.285 ;
        RECT -67.865 7.015 -67.695 7.185 ;
        RECT -66.095 7.115 -65.925 7.285 ;
        RECT -76.015 6.655 -75.845 6.825 ;
        RECT -69.635 6.655 -69.465 6.825 ;
        RECT -76.015 6.195 -75.845 6.365 ;
        RECT -69.635 6.195 -69.465 6.365 ;
        RECT -59.715 7.115 -59.545 7.285 ;
        RECT -57.945 7.015 -57.775 7.185 ;
        RECT -56.175 7.115 -56.005 7.285 ;
        RECT -66.095 6.655 -65.925 6.825 ;
        RECT -59.715 6.655 -59.545 6.825 ;
        RECT -66.095 6.195 -65.925 6.365 ;
        RECT -59.715 6.195 -59.545 6.365 ;
        RECT -49.795 7.115 -49.625 7.285 ;
        RECT -48.025 7.015 -47.855 7.185 ;
        RECT -46.255 7.115 -46.085 7.285 ;
        RECT -56.175 6.655 -56.005 6.825 ;
        RECT -49.795 6.655 -49.625 6.825 ;
        RECT -56.175 6.195 -56.005 6.365 ;
        RECT -49.795 6.195 -49.625 6.365 ;
        RECT -39.875 7.115 -39.705 7.285 ;
        RECT -38.105 7.015 -37.935 7.185 ;
        RECT -36.335 7.115 -36.165 7.285 ;
        RECT -46.255 6.655 -46.085 6.825 ;
        RECT -39.875 6.655 -39.705 6.825 ;
        RECT -46.255 6.195 -46.085 6.365 ;
        RECT -39.875 6.195 -39.705 6.365 ;
        RECT -29.955 7.115 -29.785 7.285 ;
        RECT -28.185 7.015 -28.015 7.185 ;
        RECT -26.415 7.115 -26.245 7.285 ;
        RECT -36.335 6.655 -36.165 6.825 ;
        RECT -29.955 6.655 -29.785 6.825 ;
        RECT -36.335 6.195 -36.165 6.365 ;
        RECT -29.955 6.195 -29.785 6.365 ;
        RECT -20.035 7.115 -19.865 7.285 ;
        RECT -18.265 7.015 -18.095 7.185 ;
        RECT -16.495 7.115 -16.325 7.285 ;
        RECT -26.415 6.655 -26.245 6.825 ;
        RECT -20.035 6.655 -19.865 6.825 ;
        RECT -26.415 6.195 -26.245 6.365 ;
        RECT -20.035 6.195 -19.865 6.365 ;
        RECT -10.115 7.115 -9.945 7.285 ;
        RECT -8.345 7.015 -8.175 7.185 ;
        RECT -6.575 7.115 -6.405 7.285 ;
        RECT -16.495 6.655 -16.325 6.825 ;
        RECT -10.115 6.655 -9.945 6.825 ;
        RECT -16.495 6.195 -16.325 6.365 ;
        RECT -10.115 6.195 -9.945 6.365 ;
        RECT -0.195 7.115 -0.025 7.285 ;
        RECT 1.575 7.015 1.745 7.185 ;
        RECT 3.345 7.115 3.515 7.285 ;
        RECT -6.575 6.655 -6.405 6.825 ;
        RECT -0.195 6.655 -0.025 6.825 ;
        RECT -6.575 6.195 -6.405 6.365 ;
        RECT -0.195 6.195 -0.025 6.365 ;
        RECT 9.725 7.115 9.895 7.285 ;
        RECT 11.495 7.015 11.665 7.185 ;
        RECT 13.265 7.115 13.435 7.285 ;
        RECT 3.345 6.655 3.515 6.825 ;
        RECT 9.725 6.655 9.895 6.825 ;
        RECT 3.345 6.195 3.515 6.365 ;
        RECT 9.725 6.195 9.895 6.365 ;
        RECT 19.645 7.115 19.815 7.285 ;
        RECT 21.415 7.015 21.585 7.185 ;
        RECT 23.185 7.115 23.355 7.285 ;
        RECT 13.265 6.655 13.435 6.825 ;
        RECT 19.645 6.655 19.815 6.825 ;
        RECT 13.265 6.195 13.435 6.365 ;
        RECT 19.645 6.195 19.815 6.365 ;
        RECT 23.185 6.655 23.355 6.825 ;
        RECT 23.185 6.195 23.355 6.365 ;
        RECT -282.525 5.535 -282.355 5.705 ;
        RECT -282.065 5.535 -281.895 5.705 ;
        RECT -281.605 5.535 -281.435 5.705 ;
        RECT -281.145 5.535 -280.975 5.705 ;
        RECT -280.685 5.535 -280.515 5.705 ;
        RECT -280.225 5.535 -280.055 5.705 ;
        RECT -279.765 5.535 -279.595 5.705 ;
        RECT -272.605 5.535 -272.435 5.705 ;
        RECT -272.145 5.535 -271.975 5.705 ;
        RECT -271.685 5.535 -271.515 5.705 ;
        RECT -271.225 5.535 -271.055 5.705 ;
        RECT -270.765 5.535 -270.595 5.705 ;
        RECT -270.305 5.535 -270.135 5.705 ;
        RECT -269.845 5.535 -269.675 5.705 ;
        RECT -262.685 5.535 -262.515 5.705 ;
        RECT -262.225 5.535 -262.055 5.705 ;
        RECT -261.765 5.535 -261.595 5.705 ;
        RECT -261.305 5.535 -261.135 5.705 ;
        RECT -260.845 5.535 -260.675 5.705 ;
        RECT -260.385 5.535 -260.215 5.705 ;
        RECT -259.925 5.535 -259.755 5.705 ;
        RECT -252.765 5.535 -252.595 5.705 ;
        RECT -252.305 5.535 -252.135 5.705 ;
        RECT -251.845 5.535 -251.675 5.705 ;
        RECT -251.385 5.535 -251.215 5.705 ;
        RECT -250.925 5.535 -250.755 5.705 ;
        RECT -250.465 5.535 -250.295 5.705 ;
        RECT -250.005 5.535 -249.835 5.705 ;
        RECT -242.845 5.535 -242.675 5.705 ;
        RECT -242.385 5.535 -242.215 5.705 ;
        RECT -241.925 5.535 -241.755 5.705 ;
        RECT -241.465 5.535 -241.295 5.705 ;
        RECT -241.005 5.535 -240.835 5.705 ;
        RECT -240.545 5.535 -240.375 5.705 ;
        RECT -240.085 5.535 -239.915 5.705 ;
        RECT -232.925 5.535 -232.755 5.705 ;
        RECT -232.465 5.535 -232.295 5.705 ;
        RECT -232.005 5.535 -231.835 5.705 ;
        RECT -231.545 5.535 -231.375 5.705 ;
        RECT -231.085 5.535 -230.915 5.705 ;
        RECT -230.625 5.535 -230.455 5.705 ;
        RECT -230.165 5.535 -229.995 5.705 ;
        RECT -223.005 5.535 -222.835 5.705 ;
        RECT -222.545 5.535 -222.375 5.705 ;
        RECT -222.085 5.535 -221.915 5.705 ;
        RECT -221.625 5.535 -221.455 5.705 ;
        RECT -221.165 5.535 -220.995 5.705 ;
        RECT -220.705 5.535 -220.535 5.705 ;
        RECT -220.245 5.535 -220.075 5.705 ;
        RECT -213.085 5.535 -212.915 5.705 ;
        RECT -212.625 5.535 -212.455 5.705 ;
        RECT -212.165 5.535 -211.995 5.705 ;
        RECT -211.705 5.535 -211.535 5.705 ;
        RECT -211.245 5.535 -211.075 5.705 ;
        RECT -210.785 5.535 -210.615 5.705 ;
        RECT -210.325 5.535 -210.155 5.705 ;
        RECT -203.165 5.535 -202.995 5.705 ;
        RECT -202.705 5.535 -202.535 5.705 ;
        RECT -202.245 5.535 -202.075 5.705 ;
        RECT -201.785 5.535 -201.615 5.705 ;
        RECT -201.325 5.535 -201.155 5.705 ;
        RECT -200.865 5.535 -200.695 5.705 ;
        RECT -200.405 5.535 -200.235 5.705 ;
        RECT -193.245 5.535 -193.075 5.705 ;
        RECT -192.785 5.535 -192.615 5.705 ;
        RECT -192.325 5.535 -192.155 5.705 ;
        RECT -191.865 5.535 -191.695 5.705 ;
        RECT -191.405 5.535 -191.235 5.705 ;
        RECT -190.945 5.535 -190.775 5.705 ;
        RECT -190.485 5.535 -190.315 5.705 ;
        RECT -183.325 5.535 -183.155 5.705 ;
        RECT -182.865 5.535 -182.695 5.705 ;
        RECT -182.405 5.535 -182.235 5.705 ;
        RECT -181.945 5.535 -181.775 5.705 ;
        RECT -181.485 5.535 -181.315 5.705 ;
        RECT -181.025 5.535 -180.855 5.705 ;
        RECT -180.565 5.535 -180.395 5.705 ;
        RECT -173.405 5.535 -173.235 5.705 ;
        RECT -172.945 5.535 -172.775 5.705 ;
        RECT -172.485 5.535 -172.315 5.705 ;
        RECT -172.025 5.535 -171.855 5.705 ;
        RECT -171.565 5.535 -171.395 5.705 ;
        RECT -171.105 5.535 -170.935 5.705 ;
        RECT -170.645 5.535 -170.475 5.705 ;
        RECT -163.485 5.535 -163.315 5.705 ;
        RECT -163.025 5.535 -162.855 5.705 ;
        RECT -162.565 5.535 -162.395 5.705 ;
        RECT -162.105 5.535 -161.935 5.705 ;
        RECT -161.645 5.535 -161.475 5.705 ;
        RECT -161.185 5.535 -161.015 5.705 ;
        RECT -160.725 5.535 -160.555 5.705 ;
        RECT -153.565 5.535 -153.395 5.705 ;
        RECT -153.105 5.535 -152.935 5.705 ;
        RECT -152.645 5.535 -152.475 5.705 ;
        RECT -152.185 5.535 -152.015 5.705 ;
        RECT -151.725 5.535 -151.555 5.705 ;
        RECT -151.265 5.535 -151.095 5.705 ;
        RECT -150.805 5.535 -150.635 5.705 ;
        RECT -143.645 5.535 -143.475 5.705 ;
        RECT -143.185 5.535 -143.015 5.705 ;
        RECT -142.725 5.535 -142.555 5.705 ;
        RECT -142.265 5.535 -142.095 5.705 ;
        RECT -141.805 5.535 -141.635 5.705 ;
        RECT -141.345 5.535 -141.175 5.705 ;
        RECT -140.885 5.535 -140.715 5.705 ;
        RECT -133.725 5.535 -133.555 5.705 ;
        RECT -133.265 5.535 -133.095 5.705 ;
        RECT -132.805 5.535 -132.635 5.705 ;
        RECT -132.345 5.535 -132.175 5.705 ;
        RECT -131.885 5.535 -131.715 5.705 ;
        RECT -131.425 5.535 -131.255 5.705 ;
        RECT -130.965 5.535 -130.795 5.705 ;
        RECT -123.805 5.535 -123.635 5.705 ;
        RECT -123.345 5.535 -123.175 5.705 ;
        RECT -122.885 5.535 -122.715 5.705 ;
        RECT -122.425 5.535 -122.255 5.705 ;
        RECT -121.965 5.535 -121.795 5.705 ;
        RECT -121.505 5.535 -121.335 5.705 ;
        RECT -121.045 5.535 -120.875 5.705 ;
        RECT -113.885 5.535 -113.715 5.705 ;
        RECT -113.425 5.535 -113.255 5.705 ;
        RECT -112.965 5.535 -112.795 5.705 ;
        RECT -112.505 5.535 -112.335 5.705 ;
        RECT -112.045 5.535 -111.875 5.705 ;
        RECT -111.585 5.535 -111.415 5.705 ;
        RECT -111.125 5.535 -110.955 5.705 ;
        RECT -103.965 5.535 -103.795 5.705 ;
        RECT -103.505 5.535 -103.335 5.705 ;
        RECT -103.045 5.535 -102.875 5.705 ;
        RECT -102.585 5.535 -102.415 5.705 ;
        RECT -102.125 5.535 -101.955 5.705 ;
        RECT -101.665 5.535 -101.495 5.705 ;
        RECT -101.205 5.535 -101.035 5.705 ;
        RECT -94.045 5.535 -93.875 5.705 ;
        RECT -93.585 5.535 -93.415 5.705 ;
        RECT -93.125 5.535 -92.955 5.705 ;
        RECT -92.665 5.535 -92.495 5.705 ;
        RECT -92.205 5.535 -92.035 5.705 ;
        RECT -91.745 5.535 -91.575 5.705 ;
        RECT -91.285 5.535 -91.115 5.705 ;
        RECT -84.125 5.535 -83.955 5.705 ;
        RECT -83.665 5.535 -83.495 5.705 ;
        RECT -83.205 5.535 -83.035 5.705 ;
        RECT -82.745 5.535 -82.575 5.705 ;
        RECT -82.285 5.535 -82.115 5.705 ;
        RECT -81.825 5.535 -81.655 5.705 ;
        RECT -81.365 5.535 -81.195 5.705 ;
        RECT -74.205 5.535 -74.035 5.705 ;
        RECT -73.745 5.535 -73.575 5.705 ;
        RECT -73.285 5.535 -73.115 5.705 ;
        RECT -72.825 5.535 -72.655 5.705 ;
        RECT -72.365 5.535 -72.195 5.705 ;
        RECT -71.905 5.535 -71.735 5.705 ;
        RECT -71.445 5.535 -71.275 5.705 ;
        RECT -64.285 5.535 -64.115 5.705 ;
        RECT -63.825 5.535 -63.655 5.705 ;
        RECT -63.365 5.535 -63.195 5.705 ;
        RECT -62.905 5.535 -62.735 5.705 ;
        RECT -62.445 5.535 -62.275 5.705 ;
        RECT -61.985 5.535 -61.815 5.705 ;
        RECT -61.525 5.535 -61.355 5.705 ;
        RECT -54.365 5.535 -54.195 5.705 ;
        RECT -53.905 5.535 -53.735 5.705 ;
        RECT -53.445 5.535 -53.275 5.705 ;
        RECT -52.985 5.535 -52.815 5.705 ;
        RECT -52.525 5.535 -52.355 5.705 ;
        RECT -52.065 5.535 -51.895 5.705 ;
        RECT -51.605 5.535 -51.435 5.705 ;
        RECT -44.445 5.535 -44.275 5.705 ;
        RECT -43.985 5.535 -43.815 5.705 ;
        RECT -43.525 5.535 -43.355 5.705 ;
        RECT -43.065 5.535 -42.895 5.705 ;
        RECT -42.605 5.535 -42.435 5.705 ;
        RECT -42.145 5.535 -41.975 5.705 ;
        RECT -41.685 5.535 -41.515 5.705 ;
        RECT -34.525 5.535 -34.355 5.705 ;
        RECT -34.065 5.535 -33.895 5.705 ;
        RECT -33.605 5.535 -33.435 5.705 ;
        RECT -33.145 5.535 -32.975 5.705 ;
        RECT -32.685 5.535 -32.515 5.705 ;
        RECT -32.225 5.535 -32.055 5.705 ;
        RECT -31.765 5.535 -31.595 5.705 ;
        RECT -24.605 5.535 -24.435 5.705 ;
        RECT -24.145 5.535 -23.975 5.705 ;
        RECT -23.685 5.535 -23.515 5.705 ;
        RECT -23.225 5.535 -23.055 5.705 ;
        RECT -22.765 5.535 -22.595 5.705 ;
        RECT -22.305 5.535 -22.135 5.705 ;
        RECT -21.845 5.535 -21.675 5.705 ;
        RECT -14.685 5.535 -14.515 5.705 ;
        RECT -14.225 5.535 -14.055 5.705 ;
        RECT -13.765 5.535 -13.595 5.705 ;
        RECT -13.305 5.535 -13.135 5.705 ;
        RECT -12.845 5.535 -12.675 5.705 ;
        RECT -12.385 5.535 -12.215 5.705 ;
        RECT -11.925 5.535 -11.755 5.705 ;
        RECT -4.765 5.535 -4.595 5.705 ;
        RECT -4.305 5.535 -4.135 5.705 ;
        RECT -3.845 5.535 -3.675 5.705 ;
        RECT -3.385 5.535 -3.215 5.705 ;
        RECT -2.925 5.535 -2.755 5.705 ;
        RECT -2.465 5.535 -2.295 5.705 ;
        RECT -2.005 5.535 -1.835 5.705 ;
        RECT 5.155 5.535 5.325 5.705 ;
        RECT 5.615 5.535 5.785 5.705 ;
        RECT 6.075 5.535 6.245 5.705 ;
        RECT 6.535 5.535 6.705 5.705 ;
        RECT 6.995 5.535 7.165 5.705 ;
        RECT 7.455 5.535 7.625 5.705 ;
        RECT 7.915 5.535 8.085 5.705 ;
        RECT 15.075 5.535 15.245 5.705 ;
        RECT 15.535 5.535 15.705 5.705 ;
        RECT 15.995 5.535 16.165 5.705 ;
        RECT 16.455 5.535 16.625 5.705 ;
        RECT 16.915 5.535 17.085 5.705 ;
        RECT 17.375 5.535 17.545 5.705 ;
        RECT 17.835 5.535 18.005 5.705 ;
        RECT -287.485 2.815 -287.315 2.985 ;
        RECT -287.025 2.815 -286.855 2.985 ;
        RECT -286.565 2.815 -286.395 2.985 ;
        RECT -286.105 2.815 -285.935 2.985 ;
        RECT -285.645 2.815 -285.475 2.985 ;
        RECT -285.185 2.815 -285.015 2.985 ;
        RECT -284.725 2.815 -284.555 2.985 ;
        RECT -277.565 2.815 -277.395 2.985 ;
        RECT -277.105 2.815 -276.935 2.985 ;
        RECT -276.645 2.815 -276.475 2.985 ;
        RECT -276.185 2.815 -276.015 2.985 ;
        RECT -275.725 2.815 -275.555 2.985 ;
        RECT -275.265 2.815 -275.095 2.985 ;
        RECT -274.805 2.815 -274.635 2.985 ;
        RECT -267.645 2.815 -267.475 2.985 ;
        RECT -267.185 2.815 -267.015 2.985 ;
        RECT -266.725 2.815 -266.555 2.985 ;
        RECT -266.265 2.815 -266.095 2.985 ;
        RECT -265.805 2.815 -265.635 2.985 ;
        RECT -265.345 2.815 -265.175 2.985 ;
        RECT -264.885 2.815 -264.715 2.985 ;
        RECT -257.725 2.815 -257.555 2.985 ;
        RECT -257.265 2.815 -257.095 2.985 ;
        RECT -256.805 2.815 -256.635 2.985 ;
        RECT -256.345 2.815 -256.175 2.985 ;
        RECT -255.885 2.815 -255.715 2.985 ;
        RECT -255.425 2.815 -255.255 2.985 ;
        RECT -254.965 2.815 -254.795 2.985 ;
        RECT -247.805 2.815 -247.635 2.985 ;
        RECT -247.345 2.815 -247.175 2.985 ;
        RECT -246.885 2.815 -246.715 2.985 ;
        RECT -246.425 2.815 -246.255 2.985 ;
        RECT -245.965 2.815 -245.795 2.985 ;
        RECT -245.505 2.815 -245.335 2.985 ;
        RECT -245.045 2.815 -244.875 2.985 ;
        RECT -237.885 2.815 -237.715 2.985 ;
        RECT -237.425 2.815 -237.255 2.985 ;
        RECT -236.965 2.815 -236.795 2.985 ;
        RECT -236.505 2.815 -236.335 2.985 ;
        RECT -236.045 2.815 -235.875 2.985 ;
        RECT -235.585 2.815 -235.415 2.985 ;
        RECT -235.125 2.815 -234.955 2.985 ;
        RECT -227.965 2.815 -227.795 2.985 ;
        RECT -227.505 2.815 -227.335 2.985 ;
        RECT -227.045 2.815 -226.875 2.985 ;
        RECT -226.585 2.815 -226.415 2.985 ;
        RECT -226.125 2.815 -225.955 2.985 ;
        RECT -225.665 2.815 -225.495 2.985 ;
        RECT -225.205 2.815 -225.035 2.985 ;
        RECT -218.045 2.815 -217.875 2.985 ;
        RECT -217.585 2.815 -217.415 2.985 ;
        RECT -217.125 2.815 -216.955 2.985 ;
        RECT -216.665 2.815 -216.495 2.985 ;
        RECT -216.205 2.815 -216.035 2.985 ;
        RECT -215.745 2.815 -215.575 2.985 ;
        RECT -215.285 2.815 -215.115 2.985 ;
        RECT -208.125 2.815 -207.955 2.985 ;
        RECT -207.665 2.815 -207.495 2.985 ;
        RECT -207.205 2.815 -207.035 2.985 ;
        RECT -206.745 2.815 -206.575 2.985 ;
        RECT -206.285 2.815 -206.115 2.985 ;
        RECT -205.825 2.815 -205.655 2.985 ;
        RECT -205.365 2.815 -205.195 2.985 ;
        RECT -198.205 2.815 -198.035 2.985 ;
        RECT -197.745 2.815 -197.575 2.985 ;
        RECT -197.285 2.815 -197.115 2.985 ;
        RECT -196.825 2.815 -196.655 2.985 ;
        RECT -196.365 2.815 -196.195 2.985 ;
        RECT -195.905 2.815 -195.735 2.985 ;
        RECT -195.445 2.815 -195.275 2.985 ;
        RECT -188.285 2.815 -188.115 2.985 ;
        RECT -187.825 2.815 -187.655 2.985 ;
        RECT -187.365 2.815 -187.195 2.985 ;
        RECT -186.905 2.815 -186.735 2.985 ;
        RECT -186.445 2.815 -186.275 2.985 ;
        RECT -185.985 2.815 -185.815 2.985 ;
        RECT -185.525 2.815 -185.355 2.985 ;
        RECT -178.365 2.815 -178.195 2.985 ;
        RECT -177.905 2.815 -177.735 2.985 ;
        RECT -177.445 2.815 -177.275 2.985 ;
        RECT -176.985 2.815 -176.815 2.985 ;
        RECT -176.525 2.815 -176.355 2.985 ;
        RECT -176.065 2.815 -175.895 2.985 ;
        RECT -175.605 2.815 -175.435 2.985 ;
        RECT -168.445 2.815 -168.275 2.985 ;
        RECT -167.985 2.815 -167.815 2.985 ;
        RECT -167.525 2.815 -167.355 2.985 ;
        RECT -167.065 2.815 -166.895 2.985 ;
        RECT -166.605 2.815 -166.435 2.985 ;
        RECT -166.145 2.815 -165.975 2.985 ;
        RECT -165.685 2.815 -165.515 2.985 ;
        RECT -158.525 2.815 -158.355 2.985 ;
        RECT -158.065 2.815 -157.895 2.985 ;
        RECT -157.605 2.815 -157.435 2.985 ;
        RECT -157.145 2.815 -156.975 2.985 ;
        RECT -156.685 2.815 -156.515 2.985 ;
        RECT -156.225 2.815 -156.055 2.985 ;
        RECT -155.765 2.815 -155.595 2.985 ;
        RECT -148.605 2.815 -148.435 2.985 ;
        RECT -148.145 2.815 -147.975 2.985 ;
        RECT -147.685 2.815 -147.515 2.985 ;
        RECT -147.225 2.815 -147.055 2.985 ;
        RECT -146.765 2.815 -146.595 2.985 ;
        RECT -146.305 2.815 -146.135 2.985 ;
        RECT -145.845 2.815 -145.675 2.985 ;
        RECT -138.685 2.815 -138.515 2.985 ;
        RECT -138.225 2.815 -138.055 2.985 ;
        RECT -137.765 2.815 -137.595 2.985 ;
        RECT -137.305 2.815 -137.135 2.985 ;
        RECT -136.845 2.815 -136.675 2.985 ;
        RECT -136.385 2.815 -136.215 2.985 ;
        RECT -135.925 2.815 -135.755 2.985 ;
        RECT -128.765 2.815 -128.595 2.985 ;
        RECT -128.305 2.815 -128.135 2.985 ;
        RECT -127.845 2.815 -127.675 2.985 ;
        RECT -127.385 2.815 -127.215 2.985 ;
        RECT -126.925 2.815 -126.755 2.985 ;
        RECT -126.465 2.815 -126.295 2.985 ;
        RECT -126.005 2.815 -125.835 2.985 ;
        RECT -118.845 2.815 -118.675 2.985 ;
        RECT -118.385 2.815 -118.215 2.985 ;
        RECT -117.925 2.815 -117.755 2.985 ;
        RECT -117.465 2.815 -117.295 2.985 ;
        RECT -117.005 2.815 -116.835 2.985 ;
        RECT -116.545 2.815 -116.375 2.985 ;
        RECT -116.085 2.815 -115.915 2.985 ;
        RECT -108.925 2.815 -108.755 2.985 ;
        RECT -108.465 2.815 -108.295 2.985 ;
        RECT -108.005 2.815 -107.835 2.985 ;
        RECT -107.545 2.815 -107.375 2.985 ;
        RECT -107.085 2.815 -106.915 2.985 ;
        RECT -106.625 2.815 -106.455 2.985 ;
        RECT -106.165 2.815 -105.995 2.985 ;
        RECT -99.005 2.815 -98.835 2.985 ;
        RECT -98.545 2.815 -98.375 2.985 ;
        RECT -98.085 2.815 -97.915 2.985 ;
        RECT -97.625 2.815 -97.455 2.985 ;
        RECT -97.165 2.815 -96.995 2.985 ;
        RECT -96.705 2.815 -96.535 2.985 ;
        RECT -96.245 2.815 -96.075 2.985 ;
        RECT -89.085 2.815 -88.915 2.985 ;
        RECT -88.625 2.815 -88.455 2.985 ;
        RECT -88.165 2.815 -87.995 2.985 ;
        RECT -87.705 2.815 -87.535 2.985 ;
        RECT -87.245 2.815 -87.075 2.985 ;
        RECT -86.785 2.815 -86.615 2.985 ;
        RECT -86.325 2.815 -86.155 2.985 ;
        RECT -79.165 2.815 -78.995 2.985 ;
        RECT -78.705 2.815 -78.535 2.985 ;
        RECT -78.245 2.815 -78.075 2.985 ;
        RECT -77.785 2.815 -77.615 2.985 ;
        RECT -77.325 2.815 -77.155 2.985 ;
        RECT -76.865 2.815 -76.695 2.985 ;
        RECT -76.405 2.815 -76.235 2.985 ;
        RECT -69.245 2.815 -69.075 2.985 ;
        RECT -68.785 2.815 -68.615 2.985 ;
        RECT -68.325 2.815 -68.155 2.985 ;
        RECT -67.865 2.815 -67.695 2.985 ;
        RECT -67.405 2.815 -67.235 2.985 ;
        RECT -66.945 2.815 -66.775 2.985 ;
        RECT -66.485 2.815 -66.315 2.985 ;
        RECT -59.325 2.815 -59.155 2.985 ;
        RECT -58.865 2.815 -58.695 2.985 ;
        RECT -58.405 2.815 -58.235 2.985 ;
        RECT -57.945 2.815 -57.775 2.985 ;
        RECT -57.485 2.815 -57.315 2.985 ;
        RECT -57.025 2.815 -56.855 2.985 ;
        RECT -56.565 2.815 -56.395 2.985 ;
        RECT -49.405 2.815 -49.235 2.985 ;
        RECT -48.945 2.815 -48.775 2.985 ;
        RECT -48.485 2.815 -48.315 2.985 ;
        RECT -48.025 2.815 -47.855 2.985 ;
        RECT -47.565 2.815 -47.395 2.985 ;
        RECT -47.105 2.815 -46.935 2.985 ;
        RECT -46.645 2.815 -46.475 2.985 ;
        RECT -39.485 2.815 -39.315 2.985 ;
        RECT -39.025 2.815 -38.855 2.985 ;
        RECT -38.565 2.815 -38.395 2.985 ;
        RECT -38.105 2.815 -37.935 2.985 ;
        RECT -37.645 2.815 -37.475 2.985 ;
        RECT -37.185 2.815 -37.015 2.985 ;
        RECT -36.725 2.815 -36.555 2.985 ;
        RECT -29.565 2.815 -29.395 2.985 ;
        RECT -29.105 2.815 -28.935 2.985 ;
        RECT -28.645 2.815 -28.475 2.985 ;
        RECT -28.185 2.815 -28.015 2.985 ;
        RECT -27.725 2.815 -27.555 2.985 ;
        RECT -27.265 2.815 -27.095 2.985 ;
        RECT -26.805 2.815 -26.635 2.985 ;
        RECT -19.645 2.815 -19.475 2.985 ;
        RECT -19.185 2.815 -19.015 2.985 ;
        RECT -18.725 2.815 -18.555 2.985 ;
        RECT -18.265 2.815 -18.095 2.985 ;
        RECT -17.805 2.815 -17.635 2.985 ;
        RECT -17.345 2.815 -17.175 2.985 ;
        RECT -16.885 2.815 -16.715 2.985 ;
        RECT -9.725 2.815 -9.555 2.985 ;
        RECT -9.265 2.815 -9.095 2.985 ;
        RECT -8.805 2.815 -8.635 2.985 ;
        RECT -8.345 2.815 -8.175 2.985 ;
        RECT -7.885 2.815 -7.715 2.985 ;
        RECT -7.425 2.815 -7.255 2.985 ;
        RECT -6.965 2.815 -6.795 2.985 ;
        RECT 0.195 2.815 0.365 2.985 ;
        RECT 0.655 2.815 0.825 2.985 ;
        RECT 1.115 2.815 1.285 2.985 ;
        RECT 1.575 2.815 1.745 2.985 ;
        RECT 2.035 2.815 2.205 2.985 ;
        RECT 2.495 2.815 2.665 2.985 ;
        RECT 2.955 2.815 3.125 2.985 ;
        RECT 10.115 2.815 10.285 2.985 ;
        RECT 10.575 2.815 10.745 2.985 ;
        RECT 11.035 2.815 11.205 2.985 ;
        RECT 11.495 2.815 11.665 2.985 ;
        RECT 11.955 2.815 12.125 2.985 ;
        RECT 12.415 2.815 12.585 2.985 ;
        RECT 12.875 2.815 13.045 2.985 ;
        RECT 20.035 2.815 20.205 2.985 ;
        RECT 20.495 2.815 20.665 2.985 ;
        RECT 20.955 2.815 21.125 2.985 ;
        RECT 21.415 2.815 21.585 2.985 ;
        RECT 21.875 2.815 22.045 2.985 ;
        RECT 22.335 2.815 22.505 2.985 ;
        RECT 22.795 2.815 22.965 2.985 ;
        RECT -282.915 2.155 -282.745 2.325 ;
        RECT -282.915 1.695 -282.745 1.865 ;
        RECT -279.375 2.155 -279.205 2.325 ;
        RECT -272.995 2.155 -272.825 2.325 ;
        RECT -279.375 1.695 -279.205 1.865 ;
        RECT -272.995 1.695 -272.825 1.865 ;
        RECT -281.145 1.425 -280.975 1.595 ;
        RECT -282.915 1.235 -282.745 1.405 ;
        RECT -279.375 1.235 -279.205 1.405 ;
        RECT -269.455 2.155 -269.285 2.325 ;
        RECT -263.075 2.155 -262.905 2.325 ;
        RECT -269.455 1.695 -269.285 1.865 ;
        RECT -263.075 1.695 -262.905 1.865 ;
        RECT -271.225 1.425 -271.055 1.595 ;
        RECT -272.995 1.235 -272.825 1.405 ;
        RECT -269.455 1.235 -269.285 1.405 ;
        RECT -259.535 2.155 -259.365 2.325 ;
        RECT -253.155 2.155 -252.985 2.325 ;
        RECT -259.535 1.695 -259.365 1.865 ;
        RECT -253.155 1.695 -252.985 1.865 ;
        RECT -261.305 1.425 -261.135 1.595 ;
        RECT -263.075 1.235 -262.905 1.405 ;
        RECT -259.535 1.235 -259.365 1.405 ;
        RECT -249.615 2.155 -249.445 2.325 ;
        RECT -243.235 2.155 -243.065 2.325 ;
        RECT -249.615 1.695 -249.445 1.865 ;
        RECT -243.235 1.695 -243.065 1.865 ;
        RECT -251.385 1.425 -251.215 1.595 ;
        RECT -253.155 1.235 -252.985 1.405 ;
        RECT -249.615 1.235 -249.445 1.405 ;
        RECT -239.695 2.155 -239.525 2.325 ;
        RECT -233.315 2.155 -233.145 2.325 ;
        RECT -239.695 1.695 -239.525 1.865 ;
        RECT -233.315 1.695 -233.145 1.865 ;
        RECT -241.465 1.425 -241.295 1.595 ;
        RECT -243.235 1.235 -243.065 1.405 ;
        RECT -239.695 1.235 -239.525 1.405 ;
        RECT -229.775 2.155 -229.605 2.325 ;
        RECT -223.395 2.155 -223.225 2.325 ;
        RECT -229.775 1.695 -229.605 1.865 ;
        RECT -223.395 1.695 -223.225 1.865 ;
        RECT -231.545 1.425 -231.375 1.595 ;
        RECT -233.315 1.235 -233.145 1.405 ;
        RECT -229.775 1.235 -229.605 1.405 ;
        RECT -219.855 2.155 -219.685 2.325 ;
        RECT -213.475 2.155 -213.305 2.325 ;
        RECT -219.855 1.695 -219.685 1.865 ;
        RECT -213.475 1.695 -213.305 1.865 ;
        RECT -221.625 1.425 -221.455 1.595 ;
        RECT -223.395 1.235 -223.225 1.405 ;
        RECT -219.855 1.235 -219.685 1.405 ;
        RECT -209.935 2.155 -209.765 2.325 ;
        RECT -203.555 2.155 -203.385 2.325 ;
        RECT -209.935 1.695 -209.765 1.865 ;
        RECT -203.555 1.695 -203.385 1.865 ;
        RECT -211.705 1.425 -211.535 1.595 ;
        RECT -213.475 1.235 -213.305 1.405 ;
        RECT -209.935 1.235 -209.765 1.405 ;
        RECT -200.015 2.155 -199.845 2.325 ;
        RECT -193.635 2.155 -193.465 2.325 ;
        RECT -200.015 1.695 -199.845 1.865 ;
        RECT -193.635 1.695 -193.465 1.865 ;
        RECT -201.785 1.425 -201.615 1.595 ;
        RECT -203.555 1.235 -203.385 1.405 ;
        RECT -200.015 1.235 -199.845 1.405 ;
        RECT -190.095 2.155 -189.925 2.325 ;
        RECT -183.715 2.155 -183.545 2.325 ;
        RECT -190.095 1.695 -189.925 1.865 ;
        RECT -183.715 1.695 -183.545 1.865 ;
        RECT -191.865 1.425 -191.695 1.595 ;
        RECT -193.635 1.235 -193.465 1.405 ;
        RECT -190.095 1.235 -189.925 1.405 ;
        RECT -180.175 2.155 -180.005 2.325 ;
        RECT -173.795 2.155 -173.625 2.325 ;
        RECT -180.175 1.695 -180.005 1.865 ;
        RECT -173.795 1.695 -173.625 1.865 ;
        RECT -181.945 1.425 -181.775 1.595 ;
        RECT -183.715 1.235 -183.545 1.405 ;
        RECT -180.175 1.235 -180.005 1.405 ;
        RECT -170.255 2.155 -170.085 2.325 ;
        RECT -163.875 2.155 -163.705 2.325 ;
        RECT -170.255 1.695 -170.085 1.865 ;
        RECT -163.875 1.695 -163.705 1.865 ;
        RECT -172.025 1.425 -171.855 1.595 ;
        RECT -173.795 1.235 -173.625 1.405 ;
        RECT -170.255 1.235 -170.085 1.405 ;
        RECT -160.335 2.155 -160.165 2.325 ;
        RECT -153.955 2.155 -153.785 2.325 ;
        RECT -160.335 1.695 -160.165 1.865 ;
        RECT -153.955 1.695 -153.785 1.865 ;
        RECT -162.105 1.425 -161.935 1.595 ;
        RECT -163.875 1.235 -163.705 1.405 ;
        RECT -160.335 1.235 -160.165 1.405 ;
        RECT -150.415 2.155 -150.245 2.325 ;
        RECT -144.035 2.155 -143.865 2.325 ;
        RECT -150.415 1.695 -150.245 1.865 ;
        RECT -144.035 1.695 -143.865 1.865 ;
        RECT -152.185 1.425 -152.015 1.595 ;
        RECT -153.955 1.235 -153.785 1.405 ;
        RECT -150.415 1.235 -150.245 1.405 ;
        RECT -140.495 2.155 -140.325 2.325 ;
        RECT -134.115 2.155 -133.945 2.325 ;
        RECT -140.495 1.695 -140.325 1.865 ;
        RECT -134.115 1.695 -133.945 1.865 ;
        RECT -142.265 1.425 -142.095 1.595 ;
        RECT -144.035 1.235 -143.865 1.405 ;
        RECT -140.495 1.235 -140.325 1.405 ;
        RECT -130.575 2.155 -130.405 2.325 ;
        RECT -124.195 2.155 -124.025 2.325 ;
        RECT -130.575 1.695 -130.405 1.865 ;
        RECT -124.195 1.695 -124.025 1.865 ;
        RECT -132.345 1.425 -132.175 1.595 ;
        RECT -134.115 1.235 -133.945 1.405 ;
        RECT -130.575 1.235 -130.405 1.405 ;
        RECT -120.655 2.155 -120.485 2.325 ;
        RECT -114.275 2.155 -114.105 2.325 ;
        RECT -120.655 1.695 -120.485 1.865 ;
        RECT -114.275 1.695 -114.105 1.865 ;
        RECT -122.425 1.425 -122.255 1.595 ;
        RECT -124.195 1.235 -124.025 1.405 ;
        RECT -120.655 1.235 -120.485 1.405 ;
        RECT -110.735 2.155 -110.565 2.325 ;
        RECT -104.355 2.155 -104.185 2.325 ;
        RECT -110.735 1.695 -110.565 1.865 ;
        RECT -104.355 1.695 -104.185 1.865 ;
        RECT -112.505 1.425 -112.335 1.595 ;
        RECT -114.275 1.235 -114.105 1.405 ;
        RECT -110.735 1.235 -110.565 1.405 ;
        RECT -100.815 2.155 -100.645 2.325 ;
        RECT -94.435 2.155 -94.265 2.325 ;
        RECT -100.815 1.695 -100.645 1.865 ;
        RECT -94.435 1.695 -94.265 1.865 ;
        RECT -102.585 1.425 -102.415 1.595 ;
        RECT -104.355 1.235 -104.185 1.405 ;
        RECT -100.815 1.235 -100.645 1.405 ;
        RECT -90.895 2.155 -90.725 2.325 ;
        RECT -84.515 2.155 -84.345 2.325 ;
        RECT -90.895 1.695 -90.725 1.865 ;
        RECT -84.515 1.695 -84.345 1.865 ;
        RECT -92.665 1.425 -92.495 1.595 ;
        RECT -94.435 1.235 -94.265 1.405 ;
        RECT -90.895 1.235 -90.725 1.405 ;
        RECT -80.975 2.155 -80.805 2.325 ;
        RECT -74.595 2.155 -74.425 2.325 ;
        RECT -80.975 1.695 -80.805 1.865 ;
        RECT -74.595 1.695 -74.425 1.865 ;
        RECT -82.745 1.425 -82.575 1.595 ;
        RECT -84.515 1.235 -84.345 1.405 ;
        RECT -80.975 1.235 -80.805 1.405 ;
        RECT -71.055 2.155 -70.885 2.325 ;
        RECT -64.675 2.155 -64.505 2.325 ;
        RECT -71.055 1.695 -70.885 1.865 ;
        RECT -64.675 1.695 -64.505 1.865 ;
        RECT -72.825 1.425 -72.655 1.595 ;
        RECT -74.595 1.235 -74.425 1.405 ;
        RECT -71.055 1.235 -70.885 1.405 ;
        RECT -61.135 2.155 -60.965 2.325 ;
        RECT -54.755 2.155 -54.585 2.325 ;
        RECT -61.135 1.695 -60.965 1.865 ;
        RECT -54.755 1.695 -54.585 1.865 ;
        RECT -62.905 1.425 -62.735 1.595 ;
        RECT -64.675 1.235 -64.505 1.405 ;
        RECT -61.135 1.235 -60.965 1.405 ;
        RECT -51.215 2.155 -51.045 2.325 ;
        RECT -44.835 2.155 -44.665 2.325 ;
        RECT -51.215 1.695 -51.045 1.865 ;
        RECT -44.835 1.695 -44.665 1.865 ;
        RECT -52.985 1.425 -52.815 1.595 ;
        RECT -54.755 1.235 -54.585 1.405 ;
        RECT -51.215 1.235 -51.045 1.405 ;
        RECT -41.295 2.155 -41.125 2.325 ;
        RECT -34.915 2.155 -34.745 2.325 ;
        RECT -41.295 1.695 -41.125 1.865 ;
        RECT -34.915 1.695 -34.745 1.865 ;
        RECT -43.065 1.425 -42.895 1.595 ;
        RECT -44.835 1.235 -44.665 1.405 ;
        RECT -41.295 1.235 -41.125 1.405 ;
        RECT -31.375 2.155 -31.205 2.325 ;
        RECT -24.995 2.155 -24.825 2.325 ;
        RECT -31.375 1.695 -31.205 1.865 ;
        RECT -24.995 1.695 -24.825 1.865 ;
        RECT -33.145 1.425 -32.975 1.595 ;
        RECT -34.915 1.235 -34.745 1.405 ;
        RECT -31.375 1.235 -31.205 1.405 ;
        RECT -21.455 2.155 -21.285 2.325 ;
        RECT -15.075 2.155 -14.905 2.325 ;
        RECT -21.455 1.695 -21.285 1.865 ;
        RECT -15.075 1.695 -14.905 1.865 ;
        RECT -23.225 1.425 -23.055 1.595 ;
        RECT -24.995 1.235 -24.825 1.405 ;
        RECT -21.455 1.235 -21.285 1.405 ;
        RECT -11.535 2.155 -11.365 2.325 ;
        RECT -5.155 2.155 -4.985 2.325 ;
        RECT -11.535 1.695 -11.365 1.865 ;
        RECT -5.155 1.695 -4.985 1.865 ;
        RECT -13.305 1.425 -13.135 1.595 ;
        RECT -15.075 1.235 -14.905 1.405 ;
        RECT -11.535 1.235 -11.365 1.405 ;
        RECT -1.615 2.155 -1.445 2.325 ;
        RECT 4.765 2.155 4.935 2.325 ;
        RECT -1.615 1.695 -1.445 1.865 ;
        RECT 4.765 1.695 4.935 1.865 ;
        RECT -3.385 1.425 -3.215 1.595 ;
        RECT -5.155 1.235 -4.985 1.405 ;
        RECT -1.615 1.235 -1.445 1.405 ;
        RECT 8.305 2.155 8.475 2.325 ;
        RECT 14.685 2.155 14.855 2.325 ;
        RECT 8.305 1.695 8.475 1.865 ;
        RECT 14.685 1.695 14.855 1.865 ;
        RECT 6.535 1.425 6.705 1.595 ;
        RECT 4.765 1.235 4.935 1.405 ;
        RECT 8.305 1.235 8.475 1.405 ;
        RECT 18.225 2.155 18.395 2.325 ;
        RECT 18.225 1.695 18.395 1.865 ;
        RECT 16.455 1.425 16.625 1.595 ;
        RECT 14.685 1.235 14.855 1.405 ;
        RECT 18.225 1.235 18.395 1.405 ;
        RECT -286.115 -86.235 -285.945 -86.065 ;
        RECT -284.345 -86.335 -284.175 -86.165 ;
        RECT -282.575 -86.235 -282.405 -86.065 ;
        RECT -286.115 -86.695 -285.945 -86.525 ;
        RECT -286.115 -87.155 -285.945 -86.985 ;
        RECT -276.195 -86.235 -276.025 -86.065 ;
        RECT -274.425 -86.335 -274.255 -86.165 ;
        RECT -272.655 -86.235 -272.485 -86.065 ;
        RECT -282.575 -86.695 -282.405 -86.525 ;
        RECT -276.195 -86.695 -276.025 -86.525 ;
        RECT -282.575 -87.155 -282.405 -86.985 ;
        RECT -276.195 -87.155 -276.025 -86.985 ;
        RECT -266.275 -86.235 -266.105 -86.065 ;
        RECT -264.505 -86.335 -264.335 -86.165 ;
        RECT -262.735 -86.235 -262.565 -86.065 ;
        RECT -272.655 -86.695 -272.485 -86.525 ;
        RECT -266.275 -86.695 -266.105 -86.525 ;
        RECT -272.655 -87.155 -272.485 -86.985 ;
        RECT -266.275 -87.155 -266.105 -86.985 ;
        RECT -256.355 -86.235 -256.185 -86.065 ;
        RECT -254.585 -86.335 -254.415 -86.165 ;
        RECT -252.815 -86.235 -252.645 -86.065 ;
        RECT -262.735 -86.695 -262.565 -86.525 ;
        RECT -256.355 -86.695 -256.185 -86.525 ;
        RECT -262.735 -87.155 -262.565 -86.985 ;
        RECT -256.355 -87.155 -256.185 -86.985 ;
        RECT -246.435 -86.235 -246.265 -86.065 ;
        RECT -244.665 -86.335 -244.495 -86.165 ;
        RECT -242.895 -86.235 -242.725 -86.065 ;
        RECT -252.815 -86.695 -252.645 -86.525 ;
        RECT -246.435 -86.695 -246.265 -86.525 ;
        RECT -252.815 -87.155 -252.645 -86.985 ;
        RECT -246.435 -87.155 -246.265 -86.985 ;
        RECT -236.515 -86.235 -236.345 -86.065 ;
        RECT -234.745 -86.335 -234.575 -86.165 ;
        RECT -232.975 -86.235 -232.805 -86.065 ;
        RECT -242.895 -86.695 -242.725 -86.525 ;
        RECT -236.515 -86.695 -236.345 -86.525 ;
        RECT -242.895 -87.155 -242.725 -86.985 ;
        RECT -236.515 -87.155 -236.345 -86.985 ;
        RECT -226.595 -86.235 -226.425 -86.065 ;
        RECT -224.825 -86.335 -224.655 -86.165 ;
        RECT -223.055 -86.235 -222.885 -86.065 ;
        RECT -232.975 -86.695 -232.805 -86.525 ;
        RECT -226.595 -86.695 -226.425 -86.525 ;
        RECT -232.975 -87.155 -232.805 -86.985 ;
        RECT -226.595 -87.155 -226.425 -86.985 ;
        RECT -216.675 -86.235 -216.505 -86.065 ;
        RECT -214.905 -86.335 -214.735 -86.165 ;
        RECT -213.135 -86.235 -212.965 -86.065 ;
        RECT -223.055 -86.695 -222.885 -86.525 ;
        RECT -216.675 -86.695 -216.505 -86.525 ;
        RECT -223.055 -87.155 -222.885 -86.985 ;
        RECT -216.675 -87.155 -216.505 -86.985 ;
        RECT -206.755 -86.235 -206.585 -86.065 ;
        RECT -204.985 -86.335 -204.815 -86.165 ;
        RECT -203.215 -86.235 -203.045 -86.065 ;
        RECT -213.135 -86.695 -212.965 -86.525 ;
        RECT -206.755 -86.695 -206.585 -86.525 ;
        RECT -213.135 -87.155 -212.965 -86.985 ;
        RECT -206.755 -87.155 -206.585 -86.985 ;
        RECT -196.835 -86.235 -196.665 -86.065 ;
        RECT -195.065 -86.335 -194.895 -86.165 ;
        RECT -193.295 -86.235 -193.125 -86.065 ;
        RECT -203.215 -86.695 -203.045 -86.525 ;
        RECT -196.835 -86.695 -196.665 -86.525 ;
        RECT -203.215 -87.155 -203.045 -86.985 ;
        RECT -196.835 -87.155 -196.665 -86.985 ;
        RECT -186.915 -86.235 -186.745 -86.065 ;
        RECT -185.145 -86.335 -184.975 -86.165 ;
        RECT -183.375 -86.235 -183.205 -86.065 ;
        RECT -193.295 -86.695 -193.125 -86.525 ;
        RECT -186.915 -86.695 -186.745 -86.525 ;
        RECT -193.295 -87.155 -193.125 -86.985 ;
        RECT -186.915 -87.155 -186.745 -86.985 ;
        RECT -176.995 -86.235 -176.825 -86.065 ;
        RECT -175.225 -86.335 -175.055 -86.165 ;
        RECT -173.455 -86.235 -173.285 -86.065 ;
        RECT -183.375 -86.695 -183.205 -86.525 ;
        RECT -176.995 -86.695 -176.825 -86.525 ;
        RECT -183.375 -87.155 -183.205 -86.985 ;
        RECT -176.995 -87.155 -176.825 -86.985 ;
        RECT -167.075 -86.235 -166.905 -86.065 ;
        RECT -165.305 -86.335 -165.135 -86.165 ;
        RECT -163.535 -86.235 -163.365 -86.065 ;
        RECT -173.455 -86.695 -173.285 -86.525 ;
        RECT -167.075 -86.695 -166.905 -86.525 ;
        RECT -173.455 -87.155 -173.285 -86.985 ;
        RECT -167.075 -87.155 -166.905 -86.985 ;
        RECT -157.155 -86.235 -156.985 -86.065 ;
        RECT -155.385 -86.335 -155.215 -86.165 ;
        RECT -153.615 -86.235 -153.445 -86.065 ;
        RECT -163.535 -86.695 -163.365 -86.525 ;
        RECT -157.155 -86.695 -156.985 -86.525 ;
        RECT -163.535 -87.155 -163.365 -86.985 ;
        RECT -157.155 -87.155 -156.985 -86.985 ;
        RECT -147.235 -86.235 -147.065 -86.065 ;
        RECT -145.465 -86.335 -145.295 -86.165 ;
        RECT -143.695 -86.235 -143.525 -86.065 ;
        RECT -153.615 -86.695 -153.445 -86.525 ;
        RECT -147.235 -86.695 -147.065 -86.525 ;
        RECT -153.615 -87.155 -153.445 -86.985 ;
        RECT -147.235 -87.155 -147.065 -86.985 ;
        RECT -137.315 -86.235 -137.145 -86.065 ;
        RECT -135.545 -86.335 -135.375 -86.165 ;
        RECT -133.775 -86.235 -133.605 -86.065 ;
        RECT -143.695 -86.695 -143.525 -86.525 ;
        RECT -137.315 -86.695 -137.145 -86.525 ;
        RECT -143.695 -87.155 -143.525 -86.985 ;
        RECT -137.315 -87.155 -137.145 -86.985 ;
        RECT -127.395 -86.235 -127.225 -86.065 ;
        RECT -125.625 -86.335 -125.455 -86.165 ;
        RECT -123.855 -86.235 -123.685 -86.065 ;
        RECT -133.775 -86.695 -133.605 -86.525 ;
        RECT -127.395 -86.695 -127.225 -86.525 ;
        RECT -133.775 -87.155 -133.605 -86.985 ;
        RECT -127.395 -87.155 -127.225 -86.985 ;
        RECT -117.475 -86.235 -117.305 -86.065 ;
        RECT -115.705 -86.335 -115.535 -86.165 ;
        RECT -113.935 -86.235 -113.765 -86.065 ;
        RECT -123.855 -86.695 -123.685 -86.525 ;
        RECT -117.475 -86.695 -117.305 -86.525 ;
        RECT -123.855 -87.155 -123.685 -86.985 ;
        RECT -117.475 -87.155 -117.305 -86.985 ;
        RECT -107.555 -86.235 -107.385 -86.065 ;
        RECT -105.785 -86.335 -105.615 -86.165 ;
        RECT -104.015 -86.235 -103.845 -86.065 ;
        RECT -113.935 -86.695 -113.765 -86.525 ;
        RECT -107.555 -86.695 -107.385 -86.525 ;
        RECT -113.935 -87.155 -113.765 -86.985 ;
        RECT -107.555 -87.155 -107.385 -86.985 ;
        RECT -97.635 -86.235 -97.465 -86.065 ;
        RECT -95.865 -86.335 -95.695 -86.165 ;
        RECT -94.095 -86.235 -93.925 -86.065 ;
        RECT -104.015 -86.695 -103.845 -86.525 ;
        RECT -97.635 -86.695 -97.465 -86.525 ;
        RECT -104.015 -87.155 -103.845 -86.985 ;
        RECT -97.635 -87.155 -97.465 -86.985 ;
        RECT -87.715 -86.235 -87.545 -86.065 ;
        RECT -85.945 -86.335 -85.775 -86.165 ;
        RECT -84.175 -86.235 -84.005 -86.065 ;
        RECT -94.095 -86.695 -93.925 -86.525 ;
        RECT -87.715 -86.695 -87.545 -86.525 ;
        RECT -94.095 -87.155 -93.925 -86.985 ;
        RECT -87.715 -87.155 -87.545 -86.985 ;
        RECT -77.795 -86.235 -77.625 -86.065 ;
        RECT -76.025 -86.335 -75.855 -86.165 ;
        RECT -74.255 -86.235 -74.085 -86.065 ;
        RECT -84.175 -86.695 -84.005 -86.525 ;
        RECT -77.795 -86.695 -77.625 -86.525 ;
        RECT -84.175 -87.155 -84.005 -86.985 ;
        RECT -77.795 -87.155 -77.625 -86.985 ;
        RECT -67.875 -86.235 -67.705 -86.065 ;
        RECT -66.105 -86.335 -65.935 -86.165 ;
        RECT -64.335 -86.235 -64.165 -86.065 ;
        RECT -74.255 -86.695 -74.085 -86.525 ;
        RECT -67.875 -86.695 -67.705 -86.525 ;
        RECT -74.255 -87.155 -74.085 -86.985 ;
        RECT -67.875 -87.155 -67.705 -86.985 ;
        RECT -57.955 -86.235 -57.785 -86.065 ;
        RECT -56.185 -86.335 -56.015 -86.165 ;
        RECT -54.415 -86.235 -54.245 -86.065 ;
        RECT -64.335 -86.695 -64.165 -86.525 ;
        RECT -57.955 -86.695 -57.785 -86.525 ;
        RECT -64.335 -87.155 -64.165 -86.985 ;
        RECT -57.955 -87.155 -57.785 -86.985 ;
        RECT -48.035 -86.235 -47.865 -86.065 ;
        RECT -46.265 -86.335 -46.095 -86.165 ;
        RECT -44.495 -86.235 -44.325 -86.065 ;
        RECT -54.415 -86.695 -54.245 -86.525 ;
        RECT -48.035 -86.695 -47.865 -86.525 ;
        RECT -54.415 -87.155 -54.245 -86.985 ;
        RECT -48.035 -87.155 -47.865 -86.985 ;
        RECT -38.115 -86.235 -37.945 -86.065 ;
        RECT -36.345 -86.335 -36.175 -86.165 ;
        RECT -34.575 -86.235 -34.405 -86.065 ;
        RECT -44.495 -86.695 -44.325 -86.525 ;
        RECT -38.115 -86.695 -37.945 -86.525 ;
        RECT -44.495 -87.155 -44.325 -86.985 ;
        RECT -38.115 -87.155 -37.945 -86.985 ;
        RECT -28.195 -86.235 -28.025 -86.065 ;
        RECT -26.425 -86.335 -26.255 -86.165 ;
        RECT -24.655 -86.235 -24.485 -86.065 ;
        RECT -34.575 -86.695 -34.405 -86.525 ;
        RECT -28.195 -86.695 -28.025 -86.525 ;
        RECT -34.575 -87.155 -34.405 -86.985 ;
        RECT -28.195 -87.155 -28.025 -86.985 ;
        RECT -18.275 -86.235 -18.105 -86.065 ;
        RECT -16.505 -86.335 -16.335 -86.165 ;
        RECT -14.735 -86.235 -14.565 -86.065 ;
        RECT -24.655 -86.695 -24.485 -86.525 ;
        RECT -18.275 -86.695 -18.105 -86.525 ;
        RECT -24.655 -87.155 -24.485 -86.985 ;
        RECT -18.275 -87.155 -18.105 -86.985 ;
        RECT -8.355 -86.235 -8.185 -86.065 ;
        RECT -6.585 -86.335 -6.415 -86.165 ;
        RECT -4.815 -86.235 -4.645 -86.065 ;
        RECT -14.735 -86.695 -14.565 -86.525 ;
        RECT -8.355 -86.695 -8.185 -86.525 ;
        RECT -14.735 -87.155 -14.565 -86.985 ;
        RECT -8.355 -87.155 -8.185 -86.985 ;
        RECT 1.565 -86.235 1.735 -86.065 ;
        RECT 3.335 -86.335 3.505 -86.165 ;
        RECT 5.105 -86.235 5.275 -86.065 ;
        RECT -4.815 -86.695 -4.645 -86.525 ;
        RECT 1.565 -86.695 1.735 -86.525 ;
        RECT -4.815 -87.155 -4.645 -86.985 ;
        RECT 1.565 -87.155 1.735 -86.985 ;
        RECT 11.485 -86.235 11.655 -86.065 ;
        RECT 13.255 -86.335 13.425 -86.165 ;
        RECT 15.025 -86.235 15.195 -86.065 ;
        RECT 5.105 -86.695 5.275 -86.525 ;
        RECT 11.485 -86.695 11.655 -86.525 ;
        RECT 5.105 -87.155 5.275 -86.985 ;
        RECT 11.485 -87.155 11.655 -86.985 ;
        RECT 21.405 -86.235 21.575 -86.065 ;
        RECT 23.175 -86.335 23.345 -86.165 ;
        RECT 24.945 -86.235 25.115 -86.065 ;
        RECT 15.025 -86.695 15.195 -86.525 ;
        RECT 21.405 -86.695 21.575 -86.525 ;
        RECT 15.025 -87.155 15.195 -86.985 ;
        RECT 21.405 -87.155 21.575 -86.985 ;
        RECT 24.945 -86.695 25.115 -86.525 ;
        RECT 24.945 -87.155 25.115 -86.985 ;
        RECT -280.765 -87.815 -280.595 -87.645 ;
        RECT -280.305 -87.815 -280.135 -87.645 ;
        RECT -279.845 -87.815 -279.675 -87.645 ;
        RECT -279.385 -87.815 -279.215 -87.645 ;
        RECT -278.925 -87.815 -278.755 -87.645 ;
        RECT -278.465 -87.815 -278.295 -87.645 ;
        RECT -278.005 -87.815 -277.835 -87.645 ;
        RECT -270.845 -87.815 -270.675 -87.645 ;
        RECT -270.385 -87.815 -270.215 -87.645 ;
        RECT -269.925 -87.815 -269.755 -87.645 ;
        RECT -269.465 -87.815 -269.295 -87.645 ;
        RECT -269.005 -87.815 -268.835 -87.645 ;
        RECT -268.545 -87.815 -268.375 -87.645 ;
        RECT -268.085 -87.815 -267.915 -87.645 ;
        RECT -260.925 -87.815 -260.755 -87.645 ;
        RECT -260.465 -87.815 -260.295 -87.645 ;
        RECT -260.005 -87.815 -259.835 -87.645 ;
        RECT -259.545 -87.815 -259.375 -87.645 ;
        RECT -259.085 -87.815 -258.915 -87.645 ;
        RECT -258.625 -87.815 -258.455 -87.645 ;
        RECT -258.165 -87.815 -257.995 -87.645 ;
        RECT -251.005 -87.815 -250.835 -87.645 ;
        RECT -250.545 -87.815 -250.375 -87.645 ;
        RECT -250.085 -87.815 -249.915 -87.645 ;
        RECT -249.625 -87.815 -249.455 -87.645 ;
        RECT -249.165 -87.815 -248.995 -87.645 ;
        RECT -248.705 -87.815 -248.535 -87.645 ;
        RECT -248.245 -87.815 -248.075 -87.645 ;
        RECT -241.085 -87.815 -240.915 -87.645 ;
        RECT -240.625 -87.815 -240.455 -87.645 ;
        RECT -240.165 -87.815 -239.995 -87.645 ;
        RECT -239.705 -87.815 -239.535 -87.645 ;
        RECT -239.245 -87.815 -239.075 -87.645 ;
        RECT -238.785 -87.815 -238.615 -87.645 ;
        RECT -238.325 -87.815 -238.155 -87.645 ;
        RECT -231.165 -87.815 -230.995 -87.645 ;
        RECT -230.705 -87.815 -230.535 -87.645 ;
        RECT -230.245 -87.815 -230.075 -87.645 ;
        RECT -229.785 -87.815 -229.615 -87.645 ;
        RECT -229.325 -87.815 -229.155 -87.645 ;
        RECT -228.865 -87.815 -228.695 -87.645 ;
        RECT -228.405 -87.815 -228.235 -87.645 ;
        RECT -221.245 -87.815 -221.075 -87.645 ;
        RECT -220.785 -87.815 -220.615 -87.645 ;
        RECT -220.325 -87.815 -220.155 -87.645 ;
        RECT -219.865 -87.815 -219.695 -87.645 ;
        RECT -219.405 -87.815 -219.235 -87.645 ;
        RECT -218.945 -87.815 -218.775 -87.645 ;
        RECT -218.485 -87.815 -218.315 -87.645 ;
        RECT -211.325 -87.815 -211.155 -87.645 ;
        RECT -210.865 -87.815 -210.695 -87.645 ;
        RECT -210.405 -87.815 -210.235 -87.645 ;
        RECT -209.945 -87.815 -209.775 -87.645 ;
        RECT -209.485 -87.815 -209.315 -87.645 ;
        RECT -209.025 -87.815 -208.855 -87.645 ;
        RECT -208.565 -87.815 -208.395 -87.645 ;
        RECT -201.405 -87.815 -201.235 -87.645 ;
        RECT -200.945 -87.815 -200.775 -87.645 ;
        RECT -200.485 -87.815 -200.315 -87.645 ;
        RECT -200.025 -87.815 -199.855 -87.645 ;
        RECT -199.565 -87.815 -199.395 -87.645 ;
        RECT -199.105 -87.815 -198.935 -87.645 ;
        RECT -198.645 -87.815 -198.475 -87.645 ;
        RECT -191.485 -87.815 -191.315 -87.645 ;
        RECT -191.025 -87.815 -190.855 -87.645 ;
        RECT -190.565 -87.815 -190.395 -87.645 ;
        RECT -190.105 -87.815 -189.935 -87.645 ;
        RECT -189.645 -87.815 -189.475 -87.645 ;
        RECT -189.185 -87.815 -189.015 -87.645 ;
        RECT -188.725 -87.815 -188.555 -87.645 ;
        RECT -181.565 -87.815 -181.395 -87.645 ;
        RECT -181.105 -87.815 -180.935 -87.645 ;
        RECT -180.645 -87.815 -180.475 -87.645 ;
        RECT -180.185 -87.815 -180.015 -87.645 ;
        RECT -179.725 -87.815 -179.555 -87.645 ;
        RECT -179.265 -87.815 -179.095 -87.645 ;
        RECT -178.805 -87.815 -178.635 -87.645 ;
        RECT -171.645 -87.815 -171.475 -87.645 ;
        RECT -171.185 -87.815 -171.015 -87.645 ;
        RECT -170.725 -87.815 -170.555 -87.645 ;
        RECT -170.265 -87.815 -170.095 -87.645 ;
        RECT -169.805 -87.815 -169.635 -87.645 ;
        RECT -169.345 -87.815 -169.175 -87.645 ;
        RECT -168.885 -87.815 -168.715 -87.645 ;
        RECT -161.725 -87.815 -161.555 -87.645 ;
        RECT -161.265 -87.815 -161.095 -87.645 ;
        RECT -160.805 -87.815 -160.635 -87.645 ;
        RECT -160.345 -87.815 -160.175 -87.645 ;
        RECT -159.885 -87.815 -159.715 -87.645 ;
        RECT -159.425 -87.815 -159.255 -87.645 ;
        RECT -158.965 -87.815 -158.795 -87.645 ;
        RECT -151.805 -87.815 -151.635 -87.645 ;
        RECT -151.345 -87.815 -151.175 -87.645 ;
        RECT -150.885 -87.815 -150.715 -87.645 ;
        RECT -150.425 -87.815 -150.255 -87.645 ;
        RECT -149.965 -87.815 -149.795 -87.645 ;
        RECT -149.505 -87.815 -149.335 -87.645 ;
        RECT -149.045 -87.815 -148.875 -87.645 ;
        RECT -141.885 -87.815 -141.715 -87.645 ;
        RECT -141.425 -87.815 -141.255 -87.645 ;
        RECT -140.965 -87.815 -140.795 -87.645 ;
        RECT -140.505 -87.815 -140.335 -87.645 ;
        RECT -140.045 -87.815 -139.875 -87.645 ;
        RECT -139.585 -87.815 -139.415 -87.645 ;
        RECT -139.125 -87.815 -138.955 -87.645 ;
        RECT -131.965 -87.815 -131.795 -87.645 ;
        RECT -131.505 -87.815 -131.335 -87.645 ;
        RECT -131.045 -87.815 -130.875 -87.645 ;
        RECT -130.585 -87.815 -130.415 -87.645 ;
        RECT -130.125 -87.815 -129.955 -87.645 ;
        RECT -129.665 -87.815 -129.495 -87.645 ;
        RECT -129.205 -87.815 -129.035 -87.645 ;
        RECT -122.045 -87.815 -121.875 -87.645 ;
        RECT -121.585 -87.815 -121.415 -87.645 ;
        RECT -121.125 -87.815 -120.955 -87.645 ;
        RECT -120.665 -87.815 -120.495 -87.645 ;
        RECT -120.205 -87.815 -120.035 -87.645 ;
        RECT -119.745 -87.815 -119.575 -87.645 ;
        RECT -119.285 -87.815 -119.115 -87.645 ;
        RECT -112.125 -87.815 -111.955 -87.645 ;
        RECT -111.665 -87.815 -111.495 -87.645 ;
        RECT -111.205 -87.815 -111.035 -87.645 ;
        RECT -110.745 -87.815 -110.575 -87.645 ;
        RECT -110.285 -87.815 -110.115 -87.645 ;
        RECT -109.825 -87.815 -109.655 -87.645 ;
        RECT -109.365 -87.815 -109.195 -87.645 ;
        RECT -102.205 -87.815 -102.035 -87.645 ;
        RECT -101.745 -87.815 -101.575 -87.645 ;
        RECT -101.285 -87.815 -101.115 -87.645 ;
        RECT -100.825 -87.815 -100.655 -87.645 ;
        RECT -100.365 -87.815 -100.195 -87.645 ;
        RECT -99.905 -87.815 -99.735 -87.645 ;
        RECT -99.445 -87.815 -99.275 -87.645 ;
        RECT -92.285 -87.815 -92.115 -87.645 ;
        RECT -91.825 -87.815 -91.655 -87.645 ;
        RECT -91.365 -87.815 -91.195 -87.645 ;
        RECT -90.905 -87.815 -90.735 -87.645 ;
        RECT -90.445 -87.815 -90.275 -87.645 ;
        RECT -89.985 -87.815 -89.815 -87.645 ;
        RECT -89.525 -87.815 -89.355 -87.645 ;
        RECT -82.365 -87.815 -82.195 -87.645 ;
        RECT -81.905 -87.815 -81.735 -87.645 ;
        RECT -81.445 -87.815 -81.275 -87.645 ;
        RECT -80.985 -87.815 -80.815 -87.645 ;
        RECT -80.525 -87.815 -80.355 -87.645 ;
        RECT -80.065 -87.815 -79.895 -87.645 ;
        RECT -79.605 -87.815 -79.435 -87.645 ;
        RECT -72.445 -87.815 -72.275 -87.645 ;
        RECT -71.985 -87.815 -71.815 -87.645 ;
        RECT -71.525 -87.815 -71.355 -87.645 ;
        RECT -71.065 -87.815 -70.895 -87.645 ;
        RECT -70.605 -87.815 -70.435 -87.645 ;
        RECT -70.145 -87.815 -69.975 -87.645 ;
        RECT -69.685 -87.815 -69.515 -87.645 ;
        RECT -62.525 -87.815 -62.355 -87.645 ;
        RECT -62.065 -87.815 -61.895 -87.645 ;
        RECT -61.605 -87.815 -61.435 -87.645 ;
        RECT -61.145 -87.815 -60.975 -87.645 ;
        RECT -60.685 -87.815 -60.515 -87.645 ;
        RECT -60.225 -87.815 -60.055 -87.645 ;
        RECT -59.765 -87.815 -59.595 -87.645 ;
        RECT -52.605 -87.815 -52.435 -87.645 ;
        RECT -52.145 -87.815 -51.975 -87.645 ;
        RECT -51.685 -87.815 -51.515 -87.645 ;
        RECT -51.225 -87.815 -51.055 -87.645 ;
        RECT -50.765 -87.815 -50.595 -87.645 ;
        RECT -50.305 -87.815 -50.135 -87.645 ;
        RECT -49.845 -87.815 -49.675 -87.645 ;
        RECT -42.685 -87.815 -42.515 -87.645 ;
        RECT -42.225 -87.815 -42.055 -87.645 ;
        RECT -41.765 -87.815 -41.595 -87.645 ;
        RECT -41.305 -87.815 -41.135 -87.645 ;
        RECT -40.845 -87.815 -40.675 -87.645 ;
        RECT -40.385 -87.815 -40.215 -87.645 ;
        RECT -39.925 -87.815 -39.755 -87.645 ;
        RECT -32.765 -87.815 -32.595 -87.645 ;
        RECT -32.305 -87.815 -32.135 -87.645 ;
        RECT -31.845 -87.815 -31.675 -87.645 ;
        RECT -31.385 -87.815 -31.215 -87.645 ;
        RECT -30.925 -87.815 -30.755 -87.645 ;
        RECT -30.465 -87.815 -30.295 -87.645 ;
        RECT -30.005 -87.815 -29.835 -87.645 ;
        RECT -22.845 -87.815 -22.675 -87.645 ;
        RECT -22.385 -87.815 -22.215 -87.645 ;
        RECT -21.925 -87.815 -21.755 -87.645 ;
        RECT -21.465 -87.815 -21.295 -87.645 ;
        RECT -21.005 -87.815 -20.835 -87.645 ;
        RECT -20.545 -87.815 -20.375 -87.645 ;
        RECT -20.085 -87.815 -19.915 -87.645 ;
        RECT -12.925 -87.815 -12.755 -87.645 ;
        RECT -12.465 -87.815 -12.295 -87.645 ;
        RECT -12.005 -87.815 -11.835 -87.645 ;
        RECT -11.545 -87.815 -11.375 -87.645 ;
        RECT -11.085 -87.815 -10.915 -87.645 ;
        RECT -10.625 -87.815 -10.455 -87.645 ;
        RECT -10.165 -87.815 -9.995 -87.645 ;
        RECT -3.005 -87.815 -2.835 -87.645 ;
        RECT -2.545 -87.815 -2.375 -87.645 ;
        RECT -2.085 -87.815 -1.915 -87.645 ;
        RECT -1.625 -87.815 -1.455 -87.645 ;
        RECT -1.165 -87.815 -0.995 -87.645 ;
        RECT -0.705 -87.815 -0.535 -87.645 ;
        RECT -0.245 -87.815 -0.075 -87.645 ;
        RECT 6.915 -87.815 7.085 -87.645 ;
        RECT 7.375 -87.815 7.545 -87.645 ;
        RECT 7.835 -87.815 8.005 -87.645 ;
        RECT 8.295 -87.815 8.465 -87.645 ;
        RECT 8.755 -87.815 8.925 -87.645 ;
        RECT 9.215 -87.815 9.385 -87.645 ;
        RECT 9.675 -87.815 9.845 -87.645 ;
        RECT 16.835 -87.815 17.005 -87.645 ;
        RECT 17.295 -87.815 17.465 -87.645 ;
        RECT 17.755 -87.815 17.925 -87.645 ;
        RECT 18.215 -87.815 18.385 -87.645 ;
        RECT 18.675 -87.815 18.845 -87.645 ;
        RECT 19.135 -87.815 19.305 -87.645 ;
        RECT 19.595 -87.815 19.765 -87.645 ;
        RECT -285.725 -90.535 -285.555 -90.365 ;
        RECT -285.265 -90.535 -285.095 -90.365 ;
        RECT -284.805 -90.535 -284.635 -90.365 ;
        RECT -284.345 -90.535 -284.175 -90.365 ;
        RECT -283.885 -90.535 -283.715 -90.365 ;
        RECT -283.425 -90.535 -283.255 -90.365 ;
        RECT -282.965 -90.535 -282.795 -90.365 ;
        RECT -275.805 -90.535 -275.635 -90.365 ;
        RECT -275.345 -90.535 -275.175 -90.365 ;
        RECT -274.885 -90.535 -274.715 -90.365 ;
        RECT -274.425 -90.535 -274.255 -90.365 ;
        RECT -273.965 -90.535 -273.795 -90.365 ;
        RECT -273.505 -90.535 -273.335 -90.365 ;
        RECT -273.045 -90.535 -272.875 -90.365 ;
        RECT -265.885 -90.535 -265.715 -90.365 ;
        RECT -265.425 -90.535 -265.255 -90.365 ;
        RECT -264.965 -90.535 -264.795 -90.365 ;
        RECT -264.505 -90.535 -264.335 -90.365 ;
        RECT -264.045 -90.535 -263.875 -90.365 ;
        RECT -263.585 -90.535 -263.415 -90.365 ;
        RECT -263.125 -90.535 -262.955 -90.365 ;
        RECT -255.965 -90.535 -255.795 -90.365 ;
        RECT -255.505 -90.535 -255.335 -90.365 ;
        RECT -255.045 -90.535 -254.875 -90.365 ;
        RECT -254.585 -90.535 -254.415 -90.365 ;
        RECT -254.125 -90.535 -253.955 -90.365 ;
        RECT -253.665 -90.535 -253.495 -90.365 ;
        RECT -253.205 -90.535 -253.035 -90.365 ;
        RECT -246.045 -90.535 -245.875 -90.365 ;
        RECT -245.585 -90.535 -245.415 -90.365 ;
        RECT -245.125 -90.535 -244.955 -90.365 ;
        RECT -244.665 -90.535 -244.495 -90.365 ;
        RECT -244.205 -90.535 -244.035 -90.365 ;
        RECT -243.745 -90.535 -243.575 -90.365 ;
        RECT -243.285 -90.535 -243.115 -90.365 ;
        RECT -236.125 -90.535 -235.955 -90.365 ;
        RECT -235.665 -90.535 -235.495 -90.365 ;
        RECT -235.205 -90.535 -235.035 -90.365 ;
        RECT -234.745 -90.535 -234.575 -90.365 ;
        RECT -234.285 -90.535 -234.115 -90.365 ;
        RECT -233.825 -90.535 -233.655 -90.365 ;
        RECT -233.365 -90.535 -233.195 -90.365 ;
        RECT -226.205 -90.535 -226.035 -90.365 ;
        RECT -225.745 -90.535 -225.575 -90.365 ;
        RECT -225.285 -90.535 -225.115 -90.365 ;
        RECT -224.825 -90.535 -224.655 -90.365 ;
        RECT -224.365 -90.535 -224.195 -90.365 ;
        RECT -223.905 -90.535 -223.735 -90.365 ;
        RECT -223.445 -90.535 -223.275 -90.365 ;
        RECT -216.285 -90.535 -216.115 -90.365 ;
        RECT -215.825 -90.535 -215.655 -90.365 ;
        RECT -215.365 -90.535 -215.195 -90.365 ;
        RECT -214.905 -90.535 -214.735 -90.365 ;
        RECT -214.445 -90.535 -214.275 -90.365 ;
        RECT -213.985 -90.535 -213.815 -90.365 ;
        RECT -213.525 -90.535 -213.355 -90.365 ;
        RECT -206.365 -90.535 -206.195 -90.365 ;
        RECT -205.905 -90.535 -205.735 -90.365 ;
        RECT -205.445 -90.535 -205.275 -90.365 ;
        RECT -204.985 -90.535 -204.815 -90.365 ;
        RECT -204.525 -90.535 -204.355 -90.365 ;
        RECT -204.065 -90.535 -203.895 -90.365 ;
        RECT -203.605 -90.535 -203.435 -90.365 ;
        RECT -196.445 -90.535 -196.275 -90.365 ;
        RECT -195.985 -90.535 -195.815 -90.365 ;
        RECT -195.525 -90.535 -195.355 -90.365 ;
        RECT -195.065 -90.535 -194.895 -90.365 ;
        RECT -194.605 -90.535 -194.435 -90.365 ;
        RECT -194.145 -90.535 -193.975 -90.365 ;
        RECT -193.685 -90.535 -193.515 -90.365 ;
        RECT -186.525 -90.535 -186.355 -90.365 ;
        RECT -186.065 -90.535 -185.895 -90.365 ;
        RECT -185.605 -90.535 -185.435 -90.365 ;
        RECT -185.145 -90.535 -184.975 -90.365 ;
        RECT -184.685 -90.535 -184.515 -90.365 ;
        RECT -184.225 -90.535 -184.055 -90.365 ;
        RECT -183.765 -90.535 -183.595 -90.365 ;
        RECT -176.605 -90.535 -176.435 -90.365 ;
        RECT -176.145 -90.535 -175.975 -90.365 ;
        RECT -175.685 -90.535 -175.515 -90.365 ;
        RECT -175.225 -90.535 -175.055 -90.365 ;
        RECT -174.765 -90.535 -174.595 -90.365 ;
        RECT -174.305 -90.535 -174.135 -90.365 ;
        RECT -173.845 -90.535 -173.675 -90.365 ;
        RECT -166.685 -90.535 -166.515 -90.365 ;
        RECT -166.225 -90.535 -166.055 -90.365 ;
        RECT -165.765 -90.535 -165.595 -90.365 ;
        RECT -165.305 -90.535 -165.135 -90.365 ;
        RECT -164.845 -90.535 -164.675 -90.365 ;
        RECT -164.385 -90.535 -164.215 -90.365 ;
        RECT -163.925 -90.535 -163.755 -90.365 ;
        RECT -156.765 -90.535 -156.595 -90.365 ;
        RECT -156.305 -90.535 -156.135 -90.365 ;
        RECT -155.845 -90.535 -155.675 -90.365 ;
        RECT -155.385 -90.535 -155.215 -90.365 ;
        RECT -154.925 -90.535 -154.755 -90.365 ;
        RECT -154.465 -90.535 -154.295 -90.365 ;
        RECT -154.005 -90.535 -153.835 -90.365 ;
        RECT -146.845 -90.535 -146.675 -90.365 ;
        RECT -146.385 -90.535 -146.215 -90.365 ;
        RECT -145.925 -90.535 -145.755 -90.365 ;
        RECT -145.465 -90.535 -145.295 -90.365 ;
        RECT -145.005 -90.535 -144.835 -90.365 ;
        RECT -144.545 -90.535 -144.375 -90.365 ;
        RECT -144.085 -90.535 -143.915 -90.365 ;
        RECT -136.925 -90.535 -136.755 -90.365 ;
        RECT -136.465 -90.535 -136.295 -90.365 ;
        RECT -136.005 -90.535 -135.835 -90.365 ;
        RECT -135.545 -90.535 -135.375 -90.365 ;
        RECT -135.085 -90.535 -134.915 -90.365 ;
        RECT -134.625 -90.535 -134.455 -90.365 ;
        RECT -134.165 -90.535 -133.995 -90.365 ;
        RECT -127.005 -90.535 -126.835 -90.365 ;
        RECT -126.545 -90.535 -126.375 -90.365 ;
        RECT -126.085 -90.535 -125.915 -90.365 ;
        RECT -125.625 -90.535 -125.455 -90.365 ;
        RECT -125.165 -90.535 -124.995 -90.365 ;
        RECT -124.705 -90.535 -124.535 -90.365 ;
        RECT -124.245 -90.535 -124.075 -90.365 ;
        RECT -117.085 -90.535 -116.915 -90.365 ;
        RECT -116.625 -90.535 -116.455 -90.365 ;
        RECT -116.165 -90.535 -115.995 -90.365 ;
        RECT -115.705 -90.535 -115.535 -90.365 ;
        RECT -115.245 -90.535 -115.075 -90.365 ;
        RECT -114.785 -90.535 -114.615 -90.365 ;
        RECT -114.325 -90.535 -114.155 -90.365 ;
        RECT -107.165 -90.535 -106.995 -90.365 ;
        RECT -106.705 -90.535 -106.535 -90.365 ;
        RECT -106.245 -90.535 -106.075 -90.365 ;
        RECT -105.785 -90.535 -105.615 -90.365 ;
        RECT -105.325 -90.535 -105.155 -90.365 ;
        RECT -104.865 -90.535 -104.695 -90.365 ;
        RECT -104.405 -90.535 -104.235 -90.365 ;
        RECT -97.245 -90.535 -97.075 -90.365 ;
        RECT -96.785 -90.535 -96.615 -90.365 ;
        RECT -96.325 -90.535 -96.155 -90.365 ;
        RECT -95.865 -90.535 -95.695 -90.365 ;
        RECT -95.405 -90.535 -95.235 -90.365 ;
        RECT -94.945 -90.535 -94.775 -90.365 ;
        RECT -94.485 -90.535 -94.315 -90.365 ;
        RECT -87.325 -90.535 -87.155 -90.365 ;
        RECT -86.865 -90.535 -86.695 -90.365 ;
        RECT -86.405 -90.535 -86.235 -90.365 ;
        RECT -85.945 -90.535 -85.775 -90.365 ;
        RECT -85.485 -90.535 -85.315 -90.365 ;
        RECT -85.025 -90.535 -84.855 -90.365 ;
        RECT -84.565 -90.535 -84.395 -90.365 ;
        RECT -77.405 -90.535 -77.235 -90.365 ;
        RECT -76.945 -90.535 -76.775 -90.365 ;
        RECT -76.485 -90.535 -76.315 -90.365 ;
        RECT -76.025 -90.535 -75.855 -90.365 ;
        RECT -75.565 -90.535 -75.395 -90.365 ;
        RECT -75.105 -90.535 -74.935 -90.365 ;
        RECT -74.645 -90.535 -74.475 -90.365 ;
        RECT -67.485 -90.535 -67.315 -90.365 ;
        RECT -67.025 -90.535 -66.855 -90.365 ;
        RECT -66.565 -90.535 -66.395 -90.365 ;
        RECT -66.105 -90.535 -65.935 -90.365 ;
        RECT -65.645 -90.535 -65.475 -90.365 ;
        RECT -65.185 -90.535 -65.015 -90.365 ;
        RECT -64.725 -90.535 -64.555 -90.365 ;
        RECT -57.565 -90.535 -57.395 -90.365 ;
        RECT -57.105 -90.535 -56.935 -90.365 ;
        RECT -56.645 -90.535 -56.475 -90.365 ;
        RECT -56.185 -90.535 -56.015 -90.365 ;
        RECT -55.725 -90.535 -55.555 -90.365 ;
        RECT -55.265 -90.535 -55.095 -90.365 ;
        RECT -54.805 -90.535 -54.635 -90.365 ;
        RECT -47.645 -90.535 -47.475 -90.365 ;
        RECT -47.185 -90.535 -47.015 -90.365 ;
        RECT -46.725 -90.535 -46.555 -90.365 ;
        RECT -46.265 -90.535 -46.095 -90.365 ;
        RECT -45.805 -90.535 -45.635 -90.365 ;
        RECT -45.345 -90.535 -45.175 -90.365 ;
        RECT -44.885 -90.535 -44.715 -90.365 ;
        RECT -37.725 -90.535 -37.555 -90.365 ;
        RECT -37.265 -90.535 -37.095 -90.365 ;
        RECT -36.805 -90.535 -36.635 -90.365 ;
        RECT -36.345 -90.535 -36.175 -90.365 ;
        RECT -35.885 -90.535 -35.715 -90.365 ;
        RECT -35.425 -90.535 -35.255 -90.365 ;
        RECT -34.965 -90.535 -34.795 -90.365 ;
        RECT -27.805 -90.535 -27.635 -90.365 ;
        RECT -27.345 -90.535 -27.175 -90.365 ;
        RECT -26.885 -90.535 -26.715 -90.365 ;
        RECT -26.425 -90.535 -26.255 -90.365 ;
        RECT -25.965 -90.535 -25.795 -90.365 ;
        RECT -25.505 -90.535 -25.335 -90.365 ;
        RECT -25.045 -90.535 -24.875 -90.365 ;
        RECT -17.885 -90.535 -17.715 -90.365 ;
        RECT -17.425 -90.535 -17.255 -90.365 ;
        RECT -16.965 -90.535 -16.795 -90.365 ;
        RECT -16.505 -90.535 -16.335 -90.365 ;
        RECT -16.045 -90.535 -15.875 -90.365 ;
        RECT -15.585 -90.535 -15.415 -90.365 ;
        RECT -15.125 -90.535 -14.955 -90.365 ;
        RECT -7.965 -90.535 -7.795 -90.365 ;
        RECT -7.505 -90.535 -7.335 -90.365 ;
        RECT -7.045 -90.535 -6.875 -90.365 ;
        RECT -6.585 -90.535 -6.415 -90.365 ;
        RECT -6.125 -90.535 -5.955 -90.365 ;
        RECT -5.665 -90.535 -5.495 -90.365 ;
        RECT -5.205 -90.535 -5.035 -90.365 ;
        RECT 1.955 -90.535 2.125 -90.365 ;
        RECT 2.415 -90.535 2.585 -90.365 ;
        RECT 2.875 -90.535 3.045 -90.365 ;
        RECT 3.335 -90.535 3.505 -90.365 ;
        RECT 3.795 -90.535 3.965 -90.365 ;
        RECT 4.255 -90.535 4.425 -90.365 ;
        RECT 4.715 -90.535 4.885 -90.365 ;
        RECT 11.875 -90.535 12.045 -90.365 ;
        RECT 12.335 -90.535 12.505 -90.365 ;
        RECT 12.795 -90.535 12.965 -90.365 ;
        RECT 13.255 -90.535 13.425 -90.365 ;
        RECT 13.715 -90.535 13.885 -90.365 ;
        RECT 14.175 -90.535 14.345 -90.365 ;
        RECT 14.635 -90.535 14.805 -90.365 ;
        RECT 21.795 -90.535 21.965 -90.365 ;
        RECT 22.255 -90.535 22.425 -90.365 ;
        RECT 22.715 -90.535 22.885 -90.365 ;
        RECT 23.175 -90.535 23.345 -90.365 ;
        RECT 23.635 -90.535 23.805 -90.365 ;
        RECT 24.095 -90.535 24.265 -90.365 ;
        RECT 24.555 -90.535 24.725 -90.365 ;
        RECT -281.155 -91.195 -280.985 -91.025 ;
        RECT -281.155 -91.655 -280.985 -91.485 ;
        RECT -277.615 -91.195 -277.445 -91.025 ;
        RECT -271.235 -91.195 -271.065 -91.025 ;
        RECT -277.615 -91.655 -277.445 -91.485 ;
        RECT -271.235 -91.655 -271.065 -91.485 ;
        RECT -279.385 -91.925 -279.215 -91.755 ;
        RECT -281.155 -92.115 -280.985 -91.945 ;
        RECT -277.615 -92.115 -277.445 -91.945 ;
        RECT -267.695 -91.195 -267.525 -91.025 ;
        RECT -261.315 -91.195 -261.145 -91.025 ;
        RECT -267.695 -91.655 -267.525 -91.485 ;
        RECT -261.315 -91.655 -261.145 -91.485 ;
        RECT -269.465 -91.925 -269.295 -91.755 ;
        RECT -271.235 -92.115 -271.065 -91.945 ;
        RECT -267.695 -92.115 -267.525 -91.945 ;
        RECT -257.775 -91.195 -257.605 -91.025 ;
        RECT -251.395 -91.195 -251.225 -91.025 ;
        RECT -257.775 -91.655 -257.605 -91.485 ;
        RECT -251.395 -91.655 -251.225 -91.485 ;
        RECT -259.545 -91.925 -259.375 -91.755 ;
        RECT -261.315 -92.115 -261.145 -91.945 ;
        RECT -257.775 -92.115 -257.605 -91.945 ;
        RECT -247.855 -91.195 -247.685 -91.025 ;
        RECT -241.475 -91.195 -241.305 -91.025 ;
        RECT -247.855 -91.655 -247.685 -91.485 ;
        RECT -241.475 -91.655 -241.305 -91.485 ;
        RECT -249.625 -91.925 -249.455 -91.755 ;
        RECT -251.395 -92.115 -251.225 -91.945 ;
        RECT -247.855 -92.115 -247.685 -91.945 ;
        RECT -237.935 -91.195 -237.765 -91.025 ;
        RECT -231.555 -91.195 -231.385 -91.025 ;
        RECT -237.935 -91.655 -237.765 -91.485 ;
        RECT -231.555 -91.655 -231.385 -91.485 ;
        RECT -239.705 -91.925 -239.535 -91.755 ;
        RECT -241.475 -92.115 -241.305 -91.945 ;
        RECT -237.935 -92.115 -237.765 -91.945 ;
        RECT -228.015 -91.195 -227.845 -91.025 ;
        RECT -221.635 -91.195 -221.465 -91.025 ;
        RECT -228.015 -91.655 -227.845 -91.485 ;
        RECT -221.635 -91.655 -221.465 -91.485 ;
        RECT -229.785 -91.925 -229.615 -91.755 ;
        RECT -231.555 -92.115 -231.385 -91.945 ;
        RECT -228.015 -92.115 -227.845 -91.945 ;
        RECT -218.095 -91.195 -217.925 -91.025 ;
        RECT -211.715 -91.195 -211.545 -91.025 ;
        RECT -218.095 -91.655 -217.925 -91.485 ;
        RECT -211.715 -91.655 -211.545 -91.485 ;
        RECT -219.865 -91.925 -219.695 -91.755 ;
        RECT -221.635 -92.115 -221.465 -91.945 ;
        RECT -218.095 -92.115 -217.925 -91.945 ;
        RECT -208.175 -91.195 -208.005 -91.025 ;
        RECT -201.795 -91.195 -201.625 -91.025 ;
        RECT -208.175 -91.655 -208.005 -91.485 ;
        RECT -201.795 -91.655 -201.625 -91.485 ;
        RECT -209.945 -91.925 -209.775 -91.755 ;
        RECT -211.715 -92.115 -211.545 -91.945 ;
        RECT -208.175 -92.115 -208.005 -91.945 ;
        RECT -198.255 -91.195 -198.085 -91.025 ;
        RECT -191.875 -91.195 -191.705 -91.025 ;
        RECT -198.255 -91.655 -198.085 -91.485 ;
        RECT -191.875 -91.655 -191.705 -91.485 ;
        RECT -200.025 -91.925 -199.855 -91.755 ;
        RECT -201.795 -92.115 -201.625 -91.945 ;
        RECT -198.255 -92.115 -198.085 -91.945 ;
        RECT -188.335 -91.195 -188.165 -91.025 ;
        RECT -181.955 -91.195 -181.785 -91.025 ;
        RECT -188.335 -91.655 -188.165 -91.485 ;
        RECT -181.955 -91.655 -181.785 -91.485 ;
        RECT -190.105 -91.925 -189.935 -91.755 ;
        RECT -191.875 -92.115 -191.705 -91.945 ;
        RECT -188.335 -92.115 -188.165 -91.945 ;
        RECT -178.415 -91.195 -178.245 -91.025 ;
        RECT -172.035 -91.195 -171.865 -91.025 ;
        RECT -178.415 -91.655 -178.245 -91.485 ;
        RECT -172.035 -91.655 -171.865 -91.485 ;
        RECT -180.185 -91.925 -180.015 -91.755 ;
        RECT -181.955 -92.115 -181.785 -91.945 ;
        RECT -178.415 -92.115 -178.245 -91.945 ;
        RECT -168.495 -91.195 -168.325 -91.025 ;
        RECT -162.115 -91.195 -161.945 -91.025 ;
        RECT -168.495 -91.655 -168.325 -91.485 ;
        RECT -162.115 -91.655 -161.945 -91.485 ;
        RECT -170.265 -91.925 -170.095 -91.755 ;
        RECT -172.035 -92.115 -171.865 -91.945 ;
        RECT -168.495 -92.115 -168.325 -91.945 ;
        RECT -158.575 -91.195 -158.405 -91.025 ;
        RECT -152.195 -91.195 -152.025 -91.025 ;
        RECT -158.575 -91.655 -158.405 -91.485 ;
        RECT -152.195 -91.655 -152.025 -91.485 ;
        RECT -160.345 -91.925 -160.175 -91.755 ;
        RECT -162.115 -92.115 -161.945 -91.945 ;
        RECT -158.575 -92.115 -158.405 -91.945 ;
        RECT -148.655 -91.195 -148.485 -91.025 ;
        RECT -142.275 -91.195 -142.105 -91.025 ;
        RECT -148.655 -91.655 -148.485 -91.485 ;
        RECT -142.275 -91.655 -142.105 -91.485 ;
        RECT -150.425 -91.925 -150.255 -91.755 ;
        RECT -152.195 -92.115 -152.025 -91.945 ;
        RECT -148.655 -92.115 -148.485 -91.945 ;
        RECT -138.735 -91.195 -138.565 -91.025 ;
        RECT -132.355 -91.195 -132.185 -91.025 ;
        RECT -138.735 -91.655 -138.565 -91.485 ;
        RECT -132.355 -91.655 -132.185 -91.485 ;
        RECT -140.505 -91.925 -140.335 -91.755 ;
        RECT -142.275 -92.115 -142.105 -91.945 ;
        RECT -138.735 -92.115 -138.565 -91.945 ;
        RECT -128.815 -91.195 -128.645 -91.025 ;
        RECT -122.435 -91.195 -122.265 -91.025 ;
        RECT -128.815 -91.655 -128.645 -91.485 ;
        RECT -122.435 -91.655 -122.265 -91.485 ;
        RECT -130.585 -91.925 -130.415 -91.755 ;
        RECT -132.355 -92.115 -132.185 -91.945 ;
        RECT -128.815 -92.115 -128.645 -91.945 ;
        RECT -118.895 -91.195 -118.725 -91.025 ;
        RECT -112.515 -91.195 -112.345 -91.025 ;
        RECT -118.895 -91.655 -118.725 -91.485 ;
        RECT -112.515 -91.655 -112.345 -91.485 ;
        RECT -120.665 -91.925 -120.495 -91.755 ;
        RECT -122.435 -92.115 -122.265 -91.945 ;
        RECT -118.895 -92.115 -118.725 -91.945 ;
        RECT -108.975 -91.195 -108.805 -91.025 ;
        RECT -102.595 -91.195 -102.425 -91.025 ;
        RECT -108.975 -91.655 -108.805 -91.485 ;
        RECT -102.595 -91.655 -102.425 -91.485 ;
        RECT -110.745 -91.925 -110.575 -91.755 ;
        RECT -112.515 -92.115 -112.345 -91.945 ;
        RECT -108.975 -92.115 -108.805 -91.945 ;
        RECT -99.055 -91.195 -98.885 -91.025 ;
        RECT -92.675 -91.195 -92.505 -91.025 ;
        RECT -99.055 -91.655 -98.885 -91.485 ;
        RECT -92.675 -91.655 -92.505 -91.485 ;
        RECT -100.825 -91.925 -100.655 -91.755 ;
        RECT -102.595 -92.115 -102.425 -91.945 ;
        RECT -99.055 -92.115 -98.885 -91.945 ;
        RECT -89.135 -91.195 -88.965 -91.025 ;
        RECT -82.755 -91.195 -82.585 -91.025 ;
        RECT -89.135 -91.655 -88.965 -91.485 ;
        RECT -82.755 -91.655 -82.585 -91.485 ;
        RECT -90.905 -91.925 -90.735 -91.755 ;
        RECT -92.675 -92.115 -92.505 -91.945 ;
        RECT -89.135 -92.115 -88.965 -91.945 ;
        RECT -79.215 -91.195 -79.045 -91.025 ;
        RECT -72.835 -91.195 -72.665 -91.025 ;
        RECT -79.215 -91.655 -79.045 -91.485 ;
        RECT -72.835 -91.655 -72.665 -91.485 ;
        RECT -80.985 -91.925 -80.815 -91.755 ;
        RECT -82.755 -92.115 -82.585 -91.945 ;
        RECT -79.215 -92.115 -79.045 -91.945 ;
        RECT -69.295 -91.195 -69.125 -91.025 ;
        RECT -62.915 -91.195 -62.745 -91.025 ;
        RECT -69.295 -91.655 -69.125 -91.485 ;
        RECT -62.915 -91.655 -62.745 -91.485 ;
        RECT -71.065 -91.925 -70.895 -91.755 ;
        RECT -72.835 -92.115 -72.665 -91.945 ;
        RECT -69.295 -92.115 -69.125 -91.945 ;
        RECT -59.375 -91.195 -59.205 -91.025 ;
        RECT -52.995 -91.195 -52.825 -91.025 ;
        RECT -59.375 -91.655 -59.205 -91.485 ;
        RECT -52.995 -91.655 -52.825 -91.485 ;
        RECT -61.145 -91.925 -60.975 -91.755 ;
        RECT -62.915 -92.115 -62.745 -91.945 ;
        RECT -59.375 -92.115 -59.205 -91.945 ;
        RECT -49.455 -91.195 -49.285 -91.025 ;
        RECT -43.075 -91.195 -42.905 -91.025 ;
        RECT -49.455 -91.655 -49.285 -91.485 ;
        RECT -43.075 -91.655 -42.905 -91.485 ;
        RECT -51.225 -91.925 -51.055 -91.755 ;
        RECT -52.995 -92.115 -52.825 -91.945 ;
        RECT -49.455 -92.115 -49.285 -91.945 ;
        RECT -39.535 -91.195 -39.365 -91.025 ;
        RECT -33.155 -91.195 -32.985 -91.025 ;
        RECT -39.535 -91.655 -39.365 -91.485 ;
        RECT -33.155 -91.655 -32.985 -91.485 ;
        RECT -41.305 -91.925 -41.135 -91.755 ;
        RECT -43.075 -92.115 -42.905 -91.945 ;
        RECT -39.535 -92.115 -39.365 -91.945 ;
        RECT -29.615 -91.195 -29.445 -91.025 ;
        RECT -23.235 -91.195 -23.065 -91.025 ;
        RECT -29.615 -91.655 -29.445 -91.485 ;
        RECT -23.235 -91.655 -23.065 -91.485 ;
        RECT -31.385 -91.925 -31.215 -91.755 ;
        RECT -33.155 -92.115 -32.985 -91.945 ;
        RECT -29.615 -92.115 -29.445 -91.945 ;
        RECT -19.695 -91.195 -19.525 -91.025 ;
        RECT -13.315 -91.195 -13.145 -91.025 ;
        RECT -19.695 -91.655 -19.525 -91.485 ;
        RECT -13.315 -91.655 -13.145 -91.485 ;
        RECT -21.465 -91.925 -21.295 -91.755 ;
        RECT -23.235 -92.115 -23.065 -91.945 ;
        RECT -19.695 -92.115 -19.525 -91.945 ;
        RECT -9.775 -91.195 -9.605 -91.025 ;
        RECT -3.395 -91.195 -3.225 -91.025 ;
        RECT -9.775 -91.655 -9.605 -91.485 ;
        RECT -3.395 -91.655 -3.225 -91.485 ;
        RECT -11.545 -91.925 -11.375 -91.755 ;
        RECT -13.315 -92.115 -13.145 -91.945 ;
        RECT -9.775 -92.115 -9.605 -91.945 ;
        RECT 0.145 -91.195 0.315 -91.025 ;
        RECT 6.525 -91.195 6.695 -91.025 ;
        RECT 0.145 -91.655 0.315 -91.485 ;
        RECT 6.525 -91.655 6.695 -91.485 ;
        RECT -1.625 -91.925 -1.455 -91.755 ;
        RECT -3.395 -92.115 -3.225 -91.945 ;
        RECT 0.145 -92.115 0.315 -91.945 ;
        RECT 10.065 -91.195 10.235 -91.025 ;
        RECT 16.445 -91.195 16.615 -91.025 ;
        RECT 10.065 -91.655 10.235 -91.485 ;
        RECT 16.445 -91.655 16.615 -91.485 ;
        RECT 8.295 -91.925 8.465 -91.755 ;
        RECT 6.525 -92.115 6.695 -91.945 ;
        RECT 10.065 -92.115 10.235 -91.945 ;
        RECT 19.985 -91.195 20.155 -91.025 ;
        RECT 19.985 -91.655 20.155 -91.485 ;
        RECT 18.215 -91.925 18.385 -91.755 ;
        RECT 16.445 -92.115 16.615 -91.945 ;
        RECT 19.985 -92.115 20.155 -91.945 ;
        RECT -285.865 -173.945 -285.695 -173.775 ;
        RECT -284.095 -174.045 -283.925 -173.875 ;
        RECT -282.325 -173.945 -282.155 -173.775 ;
        RECT -285.865 -174.405 -285.695 -174.235 ;
        RECT -285.865 -174.865 -285.695 -174.695 ;
        RECT -275.945 -173.945 -275.775 -173.775 ;
        RECT -274.175 -174.045 -274.005 -173.875 ;
        RECT -272.405 -173.945 -272.235 -173.775 ;
        RECT -282.325 -174.405 -282.155 -174.235 ;
        RECT -275.945 -174.405 -275.775 -174.235 ;
        RECT -282.325 -174.865 -282.155 -174.695 ;
        RECT -275.945 -174.865 -275.775 -174.695 ;
        RECT -266.025 -173.945 -265.855 -173.775 ;
        RECT -264.255 -174.045 -264.085 -173.875 ;
        RECT -262.485 -173.945 -262.315 -173.775 ;
        RECT -272.405 -174.405 -272.235 -174.235 ;
        RECT -266.025 -174.405 -265.855 -174.235 ;
        RECT -272.405 -174.865 -272.235 -174.695 ;
        RECT -266.025 -174.865 -265.855 -174.695 ;
        RECT -256.105 -173.945 -255.935 -173.775 ;
        RECT -254.335 -174.045 -254.165 -173.875 ;
        RECT -252.565 -173.945 -252.395 -173.775 ;
        RECT -262.485 -174.405 -262.315 -174.235 ;
        RECT -256.105 -174.405 -255.935 -174.235 ;
        RECT -262.485 -174.865 -262.315 -174.695 ;
        RECT -256.105 -174.865 -255.935 -174.695 ;
        RECT -246.185 -173.945 -246.015 -173.775 ;
        RECT -244.415 -174.045 -244.245 -173.875 ;
        RECT -242.645 -173.945 -242.475 -173.775 ;
        RECT -252.565 -174.405 -252.395 -174.235 ;
        RECT -246.185 -174.405 -246.015 -174.235 ;
        RECT -252.565 -174.865 -252.395 -174.695 ;
        RECT -246.185 -174.865 -246.015 -174.695 ;
        RECT -236.265 -173.945 -236.095 -173.775 ;
        RECT -234.495 -174.045 -234.325 -173.875 ;
        RECT -232.725 -173.945 -232.555 -173.775 ;
        RECT -242.645 -174.405 -242.475 -174.235 ;
        RECT -236.265 -174.405 -236.095 -174.235 ;
        RECT -242.645 -174.865 -242.475 -174.695 ;
        RECT -236.265 -174.865 -236.095 -174.695 ;
        RECT -226.345 -173.945 -226.175 -173.775 ;
        RECT -224.575 -174.045 -224.405 -173.875 ;
        RECT -222.805 -173.945 -222.635 -173.775 ;
        RECT -232.725 -174.405 -232.555 -174.235 ;
        RECT -226.345 -174.405 -226.175 -174.235 ;
        RECT -232.725 -174.865 -232.555 -174.695 ;
        RECT -226.345 -174.865 -226.175 -174.695 ;
        RECT -216.425 -173.945 -216.255 -173.775 ;
        RECT -214.655 -174.045 -214.485 -173.875 ;
        RECT -212.885 -173.945 -212.715 -173.775 ;
        RECT -222.805 -174.405 -222.635 -174.235 ;
        RECT -216.425 -174.405 -216.255 -174.235 ;
        RECT -222.805 -174.865 -222.635 -174.695 ;
        RECT -216.425 -174.865 -216.255 -174.695 ;
        RECT -206.505 -173.945 -206.335 -173.775 ;
        RECT -204.735 -174.045 -204.565 -173.875 ;
        RECT -202.965 -173.945 -202.795 -173.775 ;
        RECT -212.885 -174.405 -212.715 -174.235 ;
        RECT -206.505 -174.405 -206.335 -174.235 ;
        RECT -212.885 -174.865 -212.715 -174.695 ;
        RECT -206.505 -174.865 -206.335 -174.695 ;
        RECT -196.585 -173.945 -196.415 -173.775 ;
        RECT -194.815 -174.045 -194.645 -173.875 ;
        RECT -193.045 -173.945 -192.875 -173.775 ;
        RECT -202.965 -174.405 -202.795 -174.235 ;
        RECT -196.585 -174.405 -196.415 -174.235 ;
        RECT -202.965 -174.865 -202.795 -174.695 ;
        RECT -196.585 -174.865 -196.415 -174.695 ;
        RECT -186.665 -173.945 -186.495 -173.775 ;
        RECT -184.895 -174.045 -184.725 -173.875 ;
        RECT -183.125 -173.945 -182.955 -173.775 ;
        RECT -193.045 -174.405 -192.875 -174.235 ;
        RECT -186.665 -174.405 -186.495 -174.235 ;
        RECT -193.045 -174.865 -192.875 -174.695 ;
        RECT -186.665 -174.865 -186.495 -174.695 ;
        RECT -176.745 -173.945 -176.575 -173.775 ;
        RECT -174.975 -174.045 -174.805 -173.875 ;
        RECT -173.205 -173.945 -173.035 -173.775 ;
        RECT -183.125 -174.405 -182.955 -174.235 ;
        RECT -176.745 -174.405 -176.575 -174.235 ;
        RECT -183.125 -174.865 -182.955 -174.695 ;
        RECT -176.745 -174.865 -176.575 -174.695 ;
        RECT -166.825 -173.945 -166.655 -173.775 ;
        RECT -165.055 -174.045 -164.885 -173.875 ;
        RECT -163.285 -173.945 -163.115 -173.775 ;
        RECT -173.205 -174.405 -173.035 -174.235 ;
        RECT -166.825 -174.405 -166.655 -174.235 ;
        RECT -173.205 -174.865 -173.035 -174.695 ;
        RECT -166.825 -174.865 -166.655 -174.695 ;
        RECT -156.905 -173.945 -156.735 -173.775 ;
        RECT -155.135 -174.045 -154.965 -173.875 ;
        RECT -153.365 -173.945 -153.195 -173.775 ;
        RECT -163.285 -174.405 -163.115 -174.235 ;
        RECT -156.905 -174.405 -156.735 -174.235 ;
        RECT -163.285 -174.865 -163.115 -174.695 ;
        RECT -156.905 -174.865 -156.735 -174.695 ;
        RECT -146.985 -173.945 -146.815 -173.775 ;
        RECT -145.215 -174.045 -145.045 -173.875 ;
        RECT -143.445 -173.945 -143.275 -173.775 ;
        RECT -153.365 -174.405 -153.195 -174.235 ;
        RECT -146.985 -174.405 -146.815 -174.235 ;
        RECT -153.365 -174.865 -153.195 -174.695 ;
        RECT -146.985 -174.865 -146.815 -174.695 ;
        RECT -137.065 -173.945 -136.895 -173.775 ;
        RECT -135.295 -174.045 -135.125 -173.875 ;
        RECT -133.525 -173.945 -133.355 -173.775 ;
        RECT -143.445 -174.405 -143.275 -174.235 ;
        RECT -137.065 -174.405 -136.895 -174.235 ;
        RECT -143.445 -174.865 -143.275 -174.695 ;
        RECT -137.065 -174.865 -136.895 -174.695 ;
        RECT -127.145 -173.945 -126.975 -173.775 ;
        RECT -125.375 -174.045 -125.205 -173.875 ;
        RECT -123.605 -173.945 -123.435 -173.775 ;
        RECT -133.525 -174.405 -133.355 -174.235 ;
        RECT -127.145 -174.405 -126.975 -174.235 ;
        RECT -133.525 -174.865 -133.355 -174.695 ;
        RECT -127.145 -174.865 -126.975 -174.695 ;
        RECT -117.225 -173.945 -117.055 -173.775 ;
        RECT -115.455 -174.045 -115.285 -173.875 ;
        RECT -113.685 -173.945 -113.515 -173.775 ;
        RECT -123.605 -174.405 -123.435 -174.235 ;
        RECT -117.225 -174.405 -117.055 -174.235 ;
        RECT -123.605 -174.865 -123.435 -174.695 ;
        RECT -117.225 -174.865 -117.055 -174.695 ;
        RECT -107.305 -173.945 -107.135 -173.775 ;
        RECT -105.535 -174.045 -105.365 -173.875 ;
        RECT -103.765 -173.945 -103.595 -173.775 ;
        RECT -113.685 -174.405 -113.515 -174.235 ;
        RECT -107.305 -174.405 -107.135 -174.235 ;
        RECT -113.685 -174.865 -113.515 -174.695 ;
        RECT -107.305 -174.865 -107.135 -174.695 ;
        RECT -97.385 -173.945 -97.215 -173.775 ;
        RECT -95.615 -174.045 -95.445 -173.875 ;
        RECT -93.845 -173.945 -93.675 -173.775 ;
        RECT -103.765 -174.405 -103.595 -174.235 ;
        RECT -97.385 -174.405 -97.215 -174.235 ;
        RECT -103.765 -174.865 -103.595 -174.695 ;
        RECT -97.385 -174.865 -97.215 -174.695 ;
        RECT -87.465 -173.945 -87.295 -173.775 ;
        RECT -85.695 -174.045 -85.525 -173.875 ;
        RECT -83.925 -173.945 -83.755 -173.775 ;
        RECT -93.845 -174.405 -93.675 -174.235 ;
        RECT -87.465 -174.405 -87.295 -174.235 ;
        RECT -93.845 -174.865 -93.675 -174.695 ;
        RECT -87.465 -174.865 -87.295 -174.695 ;
        RECT -77.545 -173.945 -77.375 -173.775 ;
        RECT -75.775 -174.045 -75.605 -173.875 ;
        RECT -74.005 -173.945 -73.835 -173.775 ;
        RECT -83.925 -174.405 -83.755 -174.235 ;
        RECT -77.545 -174.405 -77.375 -174.235 ;
        RECT -83.925 -174.865 -83.755 -174.695 ;
        RECT -77.545 -174.865 -77.375 -174.695 ;
        RECT -67.625 -173.945 -67.455 -173.775 ;
        RECT -65.855 -174.045 -65.685 -173.875 ;
        RECT -64.085 -173.945 -63.915 -173.775 ;
        RECT -74.005 -174.405 -73.835 -174.235 ;
        RECT -67.625 -174.405 -67.455 -174.235 ;
        RECT -74.005 -174.865 -73.835 -174.695 ;
        RECT -67.625 -174.865 -67.455 -174.695 ;
        RECT -57.705 -173.945 -57.535 -173.775 ;
        RECT -55.935 -174.045 -55.765 -173.875 ;
        RECT -54.165 -173.945 -53.995 -173.775 ;
        RECT -64.085 -174.405 -63.915 -174.235 ;
        RECT -57.705 -174.405 -57.535 -174.235 ;
        RECT -64.085 -174.865 -63.915 -174.695 ;
        RECT -57.705 -174.865 -57.535 -174.695 ;
        RECT -47.785 -173.945 -47.615 -173.775 ;
        RECT -46.015 -174.045 -45.845 -173.875 ;
        RECT -44.245 -173.945 -44.075 -173.775 ;
        RECT -54.165 -174.405 -53.995 -174.235 ;
        RECT -47.785 -174.405 -47.615 -174.235 ;
        RECT -54.165 -174.865 -53.995 -174.695 ;
        RECT -47.785 -174.865 -47.615 -174.695 ;
        RECT -37.865 -173.945 -37.695 -173.775 ;
        RECT -36.095 -174.045 -35.925 -173.875 ;
        RECT -34.325 -173.945 -34.155 -173.775 ;
        RECT -44.245 -174.405 -44.075 -174.235 ;
        RECT -37.865 -174.405 -37.695 -174.235 ;
        RECT -44.245 -174.865 -44.075 -174.695 ;
        RECT -37.865 -174.865 -37.695 -174.695 ;
        RECT -27.945 -173.945 -27.775 -173.775 ;
        RECT -26.175 -174.045 -26.005 -173.875 ;
        RECT -24.405 -173.945 -24.235 -173.775 ;
        RECT -34.325 -174.405 -34.155 -174.235 ;
        RECT -27.945 -174.405 -27.775 -174.235 ;
        RECT -34.325 -174.865 -34.155 -174.695 ;
        RECT -27.945 -174.865 -27.775 -174.695 ;
        RECT -18.025 -173.945 -17.855 -173.775 ;
        RECT -16.255 -174.045 -16.085 -173.875 ;
        RECT -14.485 -173.945 -14.315 -173.775 ;
        RECT -24.405 -174.405 -24.235 -174.235 ;
        RECT -18.025 -174.405 -17.855 -174.235 ;
        RECT -24.405 -174.865 -24.235 -174.695 ;
        RECT -18.025 -174.865 -17.855 -174.695 ;
        RECT -8.105 -173.945 -7.935 -173.775 ;
        RECT -6.335 -174.045 -6.165 -173.875 ;
        RECT -4.565 -173.945 -4.395 -173.775 ;
        RECT -14.485 -174.405 -14.315 -174.235 ;
        RECT -8.105 -174.405 -7.935 -174.235 ;
        RECT -14.485 -174.865 -14.315 -174.695 ;
        RECT -8.105 -174.865 -7.935 -174.695 ;
        RECT 1.815 -173.945 1.985 -173.775 ;
        RECT 3.585 -174.045 3.755 -173.875 ;
        RECT 5.355 -173.945 5.525 -173.775 ;
        RECT -4.565 -174.405 -4.395 -174.235 ;
        RECT 1.815 -174.405 1.985 -174.235 ;
        RECT -4.565 -174.865 -4.395 -174.695 ;
        RECT 1.815 -174.865 1.985 -174.695 ;
        RECT 11.735 -173.945 11.905 -173.775 ;
        RECT 13.505 -174.045 13.675 -173.875 ;
        RECT 15.275 -173.945 15.445 -173.775 ;
        RECT 5.355 -174.405 5.525 -174.235 ;
        RECT 11.735 -174.405 11.905 -174.235 ;
        RECT 5.355 -174.865 5.525 -174.695 ;
        RECT 11.735 -174.865 11.905 -174.695 ;
        RECT 21.655 -173.945 21.825 -173.775 ;
        RECT 23.425 -174.045 23.595 -173.875 ;
        RECT 25.195 -173.945 25.365 -173.775 ;
        RECT 15.275 -174.405 15.445 -174.235 ;
        RECT 21.655 -174.405 21.825 -174.235 ;
        RECT 15.275 -174.865 15.445 -174.695 ;
        RECT 21.655 -174.865 21.825 -174.695 ;
        RECT 25.195 -174.405 25.365 -174.235 ;
        RECT 25.195 -174.865 25.365 -174.695 ;
        RECT -280.515 -175.525 -280.345 -175.355 ;
        RECT -280.055 -175.525 -279.885 -175.355 ;
        RECT -279.595 -175.525 -279.425 -175.355 ;
        RECT -279.135 -175.525 -278.965 -175.355 ;
        RECT -278.675 -175.525 -278.505 -175.355 ;
        RECT -278.215 -175.525 -278.045 -175.355 ;
        RECT -277.755 -175.525 -277.585 -175.355 ;
        RECT -270.595 -175.525 -270.425 -175.355 ;
        RECT -270.135 -175.525 -269.965 -175.355 ;
        RECT -269.675 -175.525 -269.505 -175.355 ;
        RECT -269.215 -175.525 -269.045 -175.355 ;
        RECT -268.755 -175.525 -268.585 -175.355 ;
        RECT -268.295 -175.525 -268.125 -175.355 ;
        RECT -267.835 -175.525 -267.665 -175.355 ;
        RECT -260.675 -175.525 -260.505 -175.355 ;
        RECT -260.215 -175.525 -260.045 -175.355 ;
        RECT -259.755 -175.525 -259.585 -175.355 ;
        RECT -259.295 -175.525 -259.125 -175.355 ;
        RECT -258.835 -175.525 -258.665 -175.355 ;
        RECT -258.375 -175.525 -258.205 -175.355 ;
        RECT -257.915 -175.525 -257.745 -175.355 ;
        RECT -250.755 -175.525 -250.585 -175.355 ;
        RECT -250.295 -175.525 -250.125 -175.355 ;
        RECT -249.835 -175.525 -249.665 -175.355 ;
        RECT -249.375 -175.525 -249.205 -175.355 ;
        RECT -248.915 -175.525 -248.745 -175.355 ;
        RECT -248.455 -175.525 -248.285 -175.355 ;
        RECT -247.995 -175.525 -247.825 -175.355 ;
        RECT -240.835 -175.525 -240.665 -175.355 ;
        RECT -240.375 -175.525 -240.205 -175.355 ;
        RECT -239.915 -175.525 -239.745 -175.355 ;
        RECT -239.455 -175.525 -239.285 -175.355 ;
        RECT -238.995 -175.525 -238.825 -175.355 ;
        RECT -238.535 -175.525 -238.365 -175.355 ;
        RECT -238.075 -175.525 -237.905 -175.355 ;
        RECT -230.915 -175.525 -230.745 -175.355 ;
        RECT -230.455 -175.525 -230.285 -175.355 ;
        RECT -229.995 -175.525 -229.825 -175.355 ;
        RECT -229.535 -175.525 -229.365 -175.355 ;
        RECT -229.075 -175.525 -228.905 -175.355 ;
        RECT -228.615 -175.525 -228.445 -175.355 ;
        RECT -228.155 -175.525 -227.985 -175.355 ;
        RECT -220.995 -175.525 -220.825 -175.355 ;
        RECT -220.535 -175.525 -220.365 -175.355 ;
        RECT -220.075 -175.525 -219.905 -175.355 ;
        RECT -219.615 -175.525 -219.445 -175.355 ;
        RECT -219.155 -175.525 -218.985 -175.355 ;
        RECT -218.695 -175.525 -218.525 -175.355 ;
        RECT -218.235 -175.525 -218.065 -175.355 ;
        RECT -211.075 -175.525 -210.905 -175.355 ;
        RECT -210.615 -175.525 -210.445 -175.355 ;
        RECT -210.155 -175.525 -209.985 -175.355 ;
        RECT -209.695 -175.525 -209.525 -175.355 ;
        RECT -209.235 -175.525 -209.065 -175.355 ;
        RECT -208.775 -175.525 -208.605 -175.355 ;
        RECT -208.315 -175.525 -208.145 -175.355 ;
        RECT -201.155 -175.525 -200.985 -175.355 ;
        RECT -200.695 -175.525 -200.525 -175.355 ;
        RECT -200.235 -175.525 -200.065 -175.355 ;
        RECT -199.775 -175.525 -199.605 -175.355 ;
        RECT -199.315 -175.525 -199.145 -175.355 ;
        RECT -198.855 -175.525 -198.685 -175.355 ;
        RECT -198.395 -175.525 -198.225 -175.355 ;
        RECT -191.235 -175.525 -191.065 -175.355 ;
        RECT -190.775 -175.525 -190.605 -175.355 ;
        RECT -190.315 -175.525 -190.145 -175.355 ;
        RECT -189.855 -175.525 -189.685 -175.355 ;
        RECT -189.395 -175.525 -189.225 -175.355 ;
        RECT -188.935 -175.525 -188.765 -175.355 ;
        RECT -188.475 -175.525 -188.305 -175.355 ;
        RECT -181.315 -175.525 -181.145 -175.355 ;
        RECT -180.855 -175.525 -180.685 -175.355 ;
        RECT -180.395 -175.525 -180.225 -175.355 ;
        RECT -179.935 -175.525 -179.765 -175.355 ;
        RECT -179.475 -175.525 -179.305 -175.355 ;
        RECT -179.015 -175.525 -178.845 -175.355 ;
        RECT -178.555 -175.525 -178.385 -175.355 ;
        RECT -171.395 -175.525 -171.225 -175.355 ;
        RECT -170.935 -175.525 -170.765 -175.355 ;
        RECT -170.475 -175.525 -170.305 -175.355 ;
        RECT -170.015 -175.525 -169.845 -175.355 ;
        RECT -169.555 -175.525 -169.385 -175.355 ;
        RECT -169.095 -175.525 -168.925 -175.355 ;
        RECT -168.635 -175.525 -168.465 -175.355 ;
        RECT -161.475 -175.525 -161.305 -175.355 ;
        RECT -161.015 -175.525 -160.845 -175.355 ;
        RECT -160.555 -175.525 -160.385 -175.355 ;
        RECT -160.095 -175.525 -159.925 -175.355 ;
        RECT -159.635 -175.525 -159.465 -175.355 ;
        RECT -159.175 -175.525 -159.005 -175.355 ;
        RECT -158.715 -175.525 -158.545 -175.355 ;
        RECT -151.555 -175.525 -151.385 -175.355 ;
        RECT -151.095 -175.525 -150.925 -175.355 ;
        RECT -150.635 -175.525 -150.465 -175.355 ;
        RECT -150.175 -175.525 -150.005 -175.355 ;
        RECT -149.715 -175.525 -149.545 -175.355 ;
        RECT -149.255 -175.525 -149.085 -175.355 ;
        RECT -148.795 -175.525 -148.625 -175.355 ;
        RECT -141.635 -175.525 -141.465 -175.355 ;
        RECT -141.175 -175.525 -141.005 -175.355 ;
        RECT -140.715 -175.525 -140.545 -175.355 ;
        RECT -140.255 -175.525 -140.085 -175.355 ;
        RECT -139.795 -175.525 -139.625 -175.355 ;
        RECT -139.335 -175.525 -139.165 -175.355 ;
        RECT -138.875 -175.525 -138.705 -175.355 ;
        RECT -131.715 -175.525 -131.545 -175.355 ;
        RECT -131.255 -175.525 -131.085 -175.355 ;
        RECT -130.795 -175.525 -130.625 -175.355 ;
        RECT -130.335 -175.525 -130.165 -175.355 ;
        RECT -129.875 -175.525 -129.705 -175.355 ;
        RECT -129.415 -175.525 -129.245 -175.355 ;
        RECT -128.955 -175.525 -128.785 -175.355 ;
        RECT -121.795 -175.525 -121.625 -175.355 ;
        RECT -121.335 -175.525 -121.165 -175.355 ;
        RECT -120.875 -175.525 -120.705 -175.355 ;
        RECT -120.415 -175.525 -120.245 -175.355 ;
        RECT -119.955 -175.525 -119.785 -175.355 ;
        RECT -119.495 -175.525 -119.325 -175.355 ;
        RECT -119.035 -175.525 -118.865 -175.355 ;
        RECT -111.875 -175.525 -111.705 -175.355 ;
        RECT -111.415 -175.525 -111.245 -175.355 ;
        RECT -110.955 -175.525 -110.785 -175.355 ;
        RECT -110.495 -175.525 -110.325 -175.355 ;
        RECT -110.035 -175.525 -109.865 -175.355 ;
        RECT -109.575 -175.525 -109.405 -175.355 ;
        RECT -109.115 -175.525 -108.945 -175.355 ;
        RECT -101.955 -175.525 -101.785 -175.355 ;
        RECT -101.495 -175.525 -101.325 -175.355 ;
        RECT -101.035 -175.525 -100.865 -175.355 ;
        RECT -100.575 -175.525 -100.405 -175.355 ;
        RECT -100.115 -175.525 -99.945 -175.355 ;
        RECT -99.655 -175.525 -99.485 -175.355 ;
        RECT -99.195 -175.525 -99.025 -175.355 ;
        RECT -92.035 -175.525 -91.865 -175.355 ;
        RECT -91.575 -175.525 -91.405 -175.355 ;
        RECT -91.115 -175.525 -90.945 -175.355 ;
        RECT -90.655 -175.525 -90.485 -175.355 ;
        RECT -90.195 -175.525 -90.025 -175.355 ;
        RECT -89.735 -175.525 -89.565 -175.355 ;
        RECT -89.275 -175.525 -89.105 -175.355 ;
        RECT -82.115 -175.525 -81.945 -175.355 ;
        RECT -81.655 -175.525 -81.485 -175.355 ;
        RECT -81.195 -175.525 -81.025 -175.355 ;
        RECT -80.735 -175.525 -80.565 -175.355 ;
        RECT -80.275 -175.525 -80.105 -175.355 ;
        RECT -79.815 -175.525 -79.645 -175.355 ;
        RECT -79.355 -175.525 -79.185 -175.355 ;
        RECT -72.195 -175.525 -72.025 -175.355 ;
        RECT -71.735 -175.525 -71.565 -175.355 ;
        RECT -71.275 -175.525 -71.105 -175.355 ;
        RECT -70.815 -175.525 -70.645 -175.355 ;
        RECT -70.355 -175.525 -70.185 -175.355 ;
        RECT -69.895 -175.525 -69.725 -175.355 ;
        RECT -69.435 -175.525 -69.265 -175.355 ;
        RECT -62.275 -175.525 -62.105 -175.355 ;
        RECT -61.815 -175.525 -61.645 -175.355 ;
        RECT -61.355 -175.525 -61.185 -175.355 ;
        RECT -60.895 -175.525 -60.725 -175.355 ;
        RECT -60.435 -175.525 -60.265 -175.355 ;
        RECT -59.975 -175.525 -59.805 -175.355 ;
        RECT -59.515 -175.525 -59.345 -175.355 ;
        RECT -52.355 -175.525 -52.185 -175.355 ;
        RECT -51.895 -175.525 -51.725 -175.355 ;
        RECT -51.435 -175.525 -51.265 -175.355 ;
        RECT -50.975 -175.525 -50.805 -175.355 ;
        RECT -50.515 -175.525 -50.345 -175.355 ;
        RECT -50.055 -175.525 -49.885 -175.355 ;
        RECT -49.595 -175.525 -49.425 -175.355 ;
        RECT -42.435 -175.525 -42.265 -175.355 ;
        RECT -41.975 -175.525 -41.805 -175.355 ;
        RECT -41.515 -175.525 -41.345 -175.355 ;
        RECT -41.055 -175.525 -40.885 -175.355 ;
        RECT -40.595 -175.525 -40.425 -175.355 ;
        RECT -40.135 -175.525 -39.965 -175.355 ;
        RECT -39.675 -175.525 -39.505 -175.355 ;
        RECT -32.515 -175.525 -32.345 -175.355 ;
        RECT -32.055 -175.525 -31.885 -175.355 ;
        RECT -31.595 -175.525 -31.425 -175.355 ;
        RECT -31.135 -175.525 -30.965 -175.355 ;
        RECT -30.675 -175.525 -30.505 -175.355 ;
        RECT -30.215 -175.525 -30.045 -175.355 ;
        RECT -29.755 -175.525 -29.585 -175.355 ;
        RECT -22.595 -175.525 -22.425 -175.355 ;
        RECT -22.135 -175.525 -21.965 -175.355 ;
        RECT -21.675 -175.525 -21.505 -175.355 ;
        RECT -21.215 -175.525 -21.045 -175.355 ;
        RECT -20.755 -175.525 -20.585 -175.355 ;
        RECT -20.295 -175.525 -20.125 -175.355 ;
        RECT -19.835 -175.525 -19.665 -175.355 ;
        RECT -12.675 -175.525 -12.505 -175.355 ;
        RECT -12.215 -175.525 -12.045 -175.355 ;
        RECT -11.755 -175.525 -11.585 -175.355 ;
        RECT -11.295 -175.525 -11.125 -175.355 ;
        RECT -10.835 -175.525 -10.665 -175.355 ;
        RECT -10.375 -175.525 -10.205 -175.355 ;
        RECT -9.915 -175.525 -9.745 -175.355 ;
        RECT -2.755 -175.525 -2.585 -175.355 ;
        RECT -2.295 -175.525 -2.125 -175.355 ;
        RECT -1.835 -175.525 -1.665 -175.355 ;
        RECT -1.375 -175.525 -1.205 -175.355 ;
        RECT -0.915 -175.525 -0.745 -175.355 ;
        RECT -0.455 -175.525 -0.285 -175.355 ;
        RECT 0.005 -175.525 0.175 -175.355 ;
        RECT 7.165 -175.525 7.335 -175.355 ;
        RECT 7.625 -175.525 7.795 -175.355 ;
        RECT 8.085 -175.525 8.255 -175.355 ;
        RECT 8.545 -175.525 8.715 -175.355 ;
        RECT 9.005 -175.525 9.175 -175.355 ;
        RECT 9.465 -175.525 9.635 -175.355 ;
        RECT 9.925 -175.525 10.095 -175.355 ;
        RECT 17.085 -175.525 17.255 -175.355 ;
        RECT 17.545 -175.525 17.715 -175.355 ;
        RECT 18.005 -175.525 18.175 -175.355 ;
        RECT 18.465 -175.525 18.635 -175.355 ;
        RECT 18.925 -175.525 19.095 -175.355 ;
        RECT 19.385 -175.525 19.555 -175.355 ;
        RECT 19.845 -175.525 20.015 -175.355 ;
        RECT -285.475 -178.245 -285.305 -178.075 ;
        RECT -285.015 -178.245 -284.845 -178.075 ;
        RECT -284.555 -178.245 -284.385 -178.075 ;
        RECT -284.095 -178.245 -283.925 -178.075 ;
        RECT -283.635 -178.245 -283.465 -178.075 ;
        RECT -283.175 -178.245 -283.005 -178.075 ;
        RECT -282.715 -178.245 -282.545 -178.075 ;
        RECT -275.555 -178.245 -275.385 -178.075 ;
        RECT -275.095 -178.245 -274.925 -178.075 ;
        RECT -274.635 -178.245 -274.465 -178.075 ;
        RECT -274.175 -178.245 -274.005 -178.075 ;
        RECT -273.715 -178.245 -273.545 -178.075 ;
        RECT -273.255 -178.245 -273.085 -178.075 ;
        RECT -272.795 -178.245 -272.625 -178.075 ;
        RECT -265.635 -178.245 -265.465 -178.075 ;
        RECT -265.175 -178.245 -265.005 -178.075 ;
        RECT -264.715 -178.245 -264.545 -178.075 ;
        RECT -264.255 -178.245 -264.085 -178.075 ;
        RECT -263.795 -178.245 -263.625 -178.075 ;
        RECT -263.335 -178.245 -263.165 -178.075 ;
        RECT -262.875 -178.245 -262.705 -178.075 ;
        RECT -255.715 -178.245 -255.545 -178.075 ;
        RECT -255.255 -178.245 -255.085 -178.075 ;
        RECT -254.795 -178.245 -254.625 -178.075 ;
        RECT -254.335 -178.245 -254.165 -178.075 ;
        RECT -253.875 -178.245 -253.705 -178.075 ;
        RECT -253.415 -178.245 -253.245 -178.075 ;
        RECT -252.955 -178.245 -252.785 -178.075 ;
        RECT -245.795 -178.245 -245.625 -178.075 ;
        RECT -245.335 -178.245 -245.165 -178.075 ;
        RECT -244.875 -178.245 -244.705 -178.075 ;
        RECT -244.415 -178.245 -244.245 -178.075 ;
        RECT -243.955 -178.245 -243.785 -178.075 ;
        RECT -243.495 -178.245 -243.325 -178.075 ;
        RECT -243.035 -178.245 -242.865 -178.075 ;
        RECT -235.875 -178.245 -235.705 -178.075 ;
        RECT -235.415 -178.245 -235.245 -178.075 ;
        RECT -234.955 -178.245 -234.785 -178.075 ;
        RECT -234.495 -178.245 -234.325 -178.075 ;
        RECT -234.035 -178.245 -233.865 -178.075 ;
        RECT -233.575 -178.245 -233.405 -178.075 ;
        RECT -233.115 -178.245 -232.945 -178.075 ;
        RECT -225.955 -178.245 -225.785 -178.075 ;
        RECT -225.495 -178.245 -225.325 -178.075 ;
        RECT -225.035 -178.245 -224.865 -178.075 ;
        RECT -224.575 -178.245 -224.405 -178.075 ;
        RECT -224.115 -178.245 -223.945 -178.075 ;
        RECT -223.655 -178.245 -223.485 -178.075 ;
        RECT -223.195 -178.245 -223.025 -178.075 ;
        RECT -216.035 -178.245 -215.865 -178.075 ;
        RECT -215.575 -178.245 -215.405 -178.075 ;
        RECT -215.115 -178.245 -214.945 -178.075 ;
        RECT -214.655 -178.245 -214.485 -178.075 ;
        RECT -214.195 -178.245 -214.025 -178.075 ;
        RECT -213.735 -178.245 -213.565 -178.075 ;
        RECT -213.275 -178.245 -213.105 -178.075 ;
        RECT -206.115 -178.245 -205.945 -178.075 ;
        RECT -205.655 -178.245 -205.485 -178.075 ;
        RECT -205.195 -178.245 -205.025 -178.075 ;
        RECT -204.735 -178.245 -204.565 -178.075 ;
        RECT -204.275 -178.245 -204.105 -178.075 ;
        RECT -203.815 -178.245 -203.645 -178.075 ;
        RECT -203.355 -178.245 -203.185 -178.075 ;
        RECT -196.195 -178.245 -196.025 -178.075 ;
        RECT -195.735 -178.245 -195.565 -178.075 ;
        RECT -195.275 -178.245 -195.105 -178.075 ;
        RECT -194.815 -178.245 -194.645 -178.075 ;
        RECT -194.355 -178.245 -194.185 -178.075 ;
        RECT -193.895 -178.245 -193.725 -178.075 ;
        RECT -193.435 -178.245 -193.265 -178.075 ;
        RECT -186.275 -178.245 -186.105 -178.075 ;
        RECT -185.815 -178.245 -185.645 -178.075 ;
        RECT -185.355 -178.245 -185.185 -178.075 ;
        RECT -184.895 -178.245 -184.725 -178.075 ;
        RECT -184.435 -178.245 -184.265 -178.075 ;
        RECT -183.975 -178.245 -183.805 -178.075 ;
        RECT -183.515 -178.245 -183.345 -178.075 ;
        RECT -176.355 -178.245 -176.185 -178.075 ;
        RECT -175.895 -178.245 -175.725 -178.075 ;
        RECT -175.435 -178.245 -175.265 -178.075 ;
        RECT -174.975 -178.245 -174.805 -178.075 ;
        RECT -174.515 -178.245 -174.345 -178.075 ;
        RECT -174.055 -178.245 -173.885 -178.075 ;
        RECT -173.595 -178.245 -173.425 -178.075 ;
        RECT -166.435 -178.245 -166.265 -178.075 ;
        RECT -165.975 -178.245 -165.805 -178.075 ;
        RECT -165.515 -178.245 -165.345 -178.075 ;
        RECT -165.055 -178.245 -164.885 -178.075 ;
        RECT -164.595 -178.245 -164.425 -178.075 ;
        RECT -164.135 -178.245 -163.965 -178.075 ;
        RECT -163.675 -178.245 -163.505 -178.075 ;
        RECT -156.515 -178.245 -156.345 -178.075 ;
        RECT -156.055 -178.245 -155.885 -178.075 ;
        RECT -155.595 -178.245 -155.425 -178.075 ;
        RECT -155.135 -178.245 -154.965 -178.075 ;
        RECT -154.675 -178.245 -154.505 -178.075 ;
        RECT -154.215 -178.245 -154.045 -178.075 ;
        RECT -153.755 -178.245 -153.585 -178.075 ;
        RECT -146.595 -178.245 -146.425 -178.075 ;
        RECT -146.135 -178.245 -145.965 -178.075 ;
        RECT -145.675 -178.245 -145.505 -178.075 ;
        RECT -145.215 -178.245 -145.045 -178.075 ;
        RECT -144.755 -178.245 -144.585 -178.075 ;
        RECT -144.295 -178.245 -144.125 -178.075 ;
        RECT -143.835 -178.245 -143.665 -178.075 ;
        RECT -136.675 -178.245 -136.505 -178.075 ;
        RECT -136.215 -178.245 -136.045 -178.075 ;
        RECT -135.755 -178.245 -135.585 -178.075 ;
        RECT -135.295 -178.245 -135.125 -178.075 ;
        RECT -134.835 -178.245 -134.665 -178.075 ;
        RECT -134.375 -178.245 -134.205 -178.075 ;
        RECT -133.915 -178.245 -133.745 -178.075 ;
        RECT -126.755 -178.245 -126.585 -178.075 ;
        RECT -126.295 -178.245 -126.125 -178.075 ;
        RECT -125.835 -178.245 -125.665 -178.075 ;
        RECT -125.375 -178.245 -125.205 -178.075 ;
        RECT -124.915 -178.245 -124.745 -178.075 ;
        RECT -124.455 -178.245 -124.285 -178.075 ;
        RECT -123.995 -178.245 -123.825 -178.075 ;
        RECT -116.835 -178.245 -116.665 -178.075 ;
        RECT -116.375 -178.245 -116.205 -178.075 ;
        RECT -115.915 -178.245 -115.745 -178.075 ;
        RECT -115.455 -178.245 -115.285 -178.075 ;
        RECT -114.995 -178.245 -114.825 -178.075 ;
        RECT -114.535 -178.245 -114.365 -178.075 ;
        RECT -114.075 -178.245 -113.905 -178.075 ;
        RECT -106.915 -178.245 -106.745 -178.075 ;
        RECT -106.455 -178.245 -106.285 -178.075 ;
        RECT -105.995 -178.245 -105.825 -178.075 ;
        RECT -105.535 -178.245 -105.365 -178.075 ;
        RECT -105.075 -178.245 -104.905 -178.075 ;
        RECT -104.615 -178.245 -104.445 -178.075 ;
        RECT -104.155 -178.245 -103.985 -178.075 ;
        RECT -96.995 -178.245 -96.825 -178.075 ;
        RECT -96.535 -178.245 -96.365 -178.075 ;
        RECT -96.075 -178.245 -95.905 -178.075 ;
        RECT -95.615 -178.245 -95.445 -178.075 ;
        RECT -95.155 -178.245 -94.985 -178.075 ;
        RECT -94.695 -178.245 -94.525 -178.075 ;
        RECT -94.235 -178.245 -94.065 -178.075 ;
        RECT -87.075 -178.245 -86.905 -178.075 ;
        RECT -86.615 -178.245 -86.445 -178.075 ;
        RECT -86.155 -178.245 -85.985 -178.075 ;
        RECT -85.695 -178.245 -85.525 -178.075 ;
        RECT -85.235 -178.245 -85.065 -178.075 ;
        RECT -84.775 -178.245 -84.605 -178.075 ;
        RECT -84.315 -178.245 -84.145 -178.075 ;
        RECT -77.155 -178.245 -76.985 -178.075 ;
        RECT -76.695 -178.245 -76.525 -178.075 ;
        RECT -76.235 -178.245 -76.065 -178.075 ;
        RECT -75.775 -178.245 -75.605 -178.075 ;
        RECT -75.315 -178.245 -75.145 -178.075 ;
        RECT -74.855 -178.245 -74.685 -178.075 ;
        RECT -74.395 -178.245 -74.225 -178.075 ;
        RECT -67.235 -178.245 -67.065 -178.075 ;
        RECT -66.775 -178.245 -66.605 -178.075 ;
        RECT -66.315 -178.245 -66.145 -178.075 ;
        RECT -65.855 -178.245 -65.685 -178.075 ;
        RECT -65.395 -178.245 -65.225 -178.075 ;
        RECT -64.935 -178.245 -64.765 -178.075 ;
        RECT -64.475 -178.245 -64.305 -178.075 ;
        RECT -57.315 -178.245 -57.145 -178.075 ;
        RECT -56.855 -178.245 -56.685 -178.075 ;
        RECT -56.395 -178.245 -56.225 -178.075 ;
        RECT -55.935 -178.245 -55.765 -178.075 ;
        RECT -55.475 -178.245 -55.305 -178.075 ;
        RECT -55.015 -178.245 -54.845 -178.075 ;
        RECT -54.555 -178.245 -54.385 -178.075 ;
        RECT -47.395 -178.245 -47.225 -178.075 ;
        RECT -46.935 -178.245 -46.765 -178.075 ;
        RECT -46.475 -178.245 -46.305 -178.075 ;
        RECT -46.015 -178.245 -45.845 -178.075 ;
        RECT -45.555 -178.245 -45.385 -178.075 ;
        RECT -45.095 -178.245 -44.925 -178.075 ;
        RECT -44.635 -178.245 -44.465 -178.075 ;
        RECT -37.475 -178.245 -37.305 -178.075 ;
        RECT -37.015 -178.245 -36.845 -178.075 ;
        RECT -36.555 -178.245 -36.385 -178.075 ;
        RECT -36.095 -178.245 -35.925 -178.075 ;
        RECT -35.635 -178.245 -35.465 -178.075 ;
        RECT -35.175 -178.245 -35.005 -178.075 ;
        RECT -34.715 -178.245 -34.545 -178.075 ;
        RECT -27.555 -178.245 -27.385 -178.075 ;
        RECT -27.095 -178.245 -26.925 -178.075 ;
        RECT -26.635 -178.245 -26.465 -178.075 ;
        RECT -26.175 -178.245 -26.005 -178.075 ;
        RECT -25.715 -178.245 -25.545 -178.075 ;
        RECT -25.255 -178.245 -25.085 -178.075 ;
        RECT -24.795 -178.245 -24.625 -178.075 ;
        RECT -17.635 -178.245 -17.465 -178.075 ;
        RECT -17.175 -178.245 -17.005 -178.075 ;
        RECT -16.715 -178.245 -16.545 -178.075 ;
        RECT -16.255 -178.245 -16.085 -178.075 ;
        RECT -15.795 -178.245 -15.625 -178.075 ;
        RECT -15.335 -178.245 -15.165 -178.075 ;
        RECT -14.875 -178.245 -14.705 -178.075 ;
        RECT -7.715 -178.245 -7.545 -178.075 ;
        RECT -7.255 -178.245 -7.085 -178.075 ;
        RECT -6.795 -178.245 -6.625 -178.075 ;
        RECT -6.335 -178.245 -6.165 -178.075 ;
        RECT -5.875 -178.245 -5.705 -178.075 ;
        RECT -5.415 -178.245 -5.245 -178.075 ;
        RECT -4.955 -178.245 -4.785 -178.075 ;
        RECT 2.205 -178.245 2.375 -178.075 ;
        RECT 2.665 -178.245 2.835 -178.075 ;
        RECT 3.125 -178.245 3.295 -178.075 ;
        RECT 3.585 -178.245 3.755 -178.075 ;
        RECT 4.045 -178.245 4.215 -178.075 ;
        RECT 4.505 -178.245 4.675 -178.075 ;
        RECT 4.965 -178.245 5.135 -178.075 ;
        RECT 12.125 -178.245 12.295 -178.075 ;
        RECT 12.585 -178.245 12.755 -178.075 ;
        RECT 13.045 -178.245 13.215 -178.075 ;
        RECT 13.505 -178.245 13.675 -178.075 ;
        RECT 13.965 -178.245 14.135 -178.075 ;
        RECT 14.425 -178.245 14.595 -178.075 ;
        RECT 14.885 -178.245 15.055 -178.075 ;
        RECT 22.045 -178.245 22.215 -178.075 ;
        RECT 22.505 -178.245 22.675 -178.075 ;
        RECT 22.965 -178.245 23.135 -178.075 ;
        RECT 23.425 -178.245 23.595 -178.075 ;
        RECT 23.885 -178.245 24.055 -178.075 ;
        RECT 24.345 -178.245 24.515 -178.075 ;
        RECT 24.805 -178.245 24.975 -178.075 ;
        RECT -280.905 -178.905 -280.735 -178.735 ;
        RECT -280.905 -179.365 -280.735 -179.195 ;
        RECT -277.365 -178.905 -277.195 -178.735 ;
        RECT -270.985 -178.905 -270.815 -178.735 ;
        RECT -277.365 -179.365 -277.195 -179.195 ;
        RECT -270.985 -179.365 -270.815 -179.195 ;
        RECT -279.135 -179.635 -278.965 -179.465 ;
        RECT -280.905 -179.825 -280.735 -179.655 ;
        RECT -277.365 -179.825 -277.195 -179.655 ;
        RECT -267.445 -178.905 -267.275 -178.735 ;
        RECT -261.065 -178.905 -260.895 -178.735 ;
        RECT -267.445 -179.365 -267.275 -179.195 ;
        RECT -261.065 -179.365 -260.895 -179.195 ;
        RECT -269.215 -179.635 -269.045 -179.465 ;
        RECT -270.985 -179.825 -270.815 -179.655 ;
        RECT -267.445 -179.825 -267.275 -179.655 ;
        RECT -257.525 -178.905 -257.355 -178.735 ;
        RECT -251.145 -178.905 -250.975 -178.735 ;
        RECT -257.525 -179.365 -257.355 -179.195 ;
        RECT -251.145 -179.365 -250.975 -179.195 ;
        RECT -259.295 -179.635 -259.125 -179.465 ;
        RECT -261.065 -179.825 -260.895 -179.655 ;
        RECT -257.525 -179.825 -257.355 -179.655 ;
        RECT -247.605 -178.905 -247.435 -178.735 ;
        RECT -241.225 -178.905 -241.055 -178.735 ;
        RECT -247.605 -179.365 -247.435 -179.195 ;
        RECT -241.225 -179.365 -241.055 -179.195 ;
        RECT -249.375 -179.635 -249.205 -179.465 ;
        RECT -251.145 -179.825 -250.975 -179.655 ;
        RECT -247.605 -179.825 -247.435 -179.655 ;
        RECT -237.685 -178.905 -237.515 -178.735 ;
        RECT -231.305 -178.905 -231.135 -178.735 ;
        RECT -237.685 -179.365 -237.515 -179.195 ;
        RECT -231.305 -179.365 -231.135 -179.195 ;
        RECT -239.455 -179.635 -239.285 -179.465 ;
        RECT -241.225 -179.825 -241.055 -179.655 ;
        RECT -237.685 -179.825 -237.515 -179.655 ;
        RECT -227.765 -178.905 -227.595 -178.735 ;
        RECT -221.385 -178.905 -221.215 -178.735 ;
        RECT -227.765 -179.365 -227.595 -179.195 ;
        RECT -221.385 -179.365 -221.215 -179.195 ;
        RECT -229.535 -179.635 -229.365 -179.465 ;
        RECT -231.305 -179.825 -231.135 -179.655 ;
        RECT -227.765 -179.825 -227.595 -179.655 ;
        RECT -217.845 -178.905 -217.675 -178.735 ;
        RECT -211.465 -178.905 -211.295 -178.735 ;
        RECT -217.845 -179.365 -217.675 -179.195 ;
        RECT -211.465 -179.365 -211.295 -179.195 ;
        RECT -219.615 -179.635 -219.445 -179.465 ;
        RECT -221.385 -179.825 -221.215 -179.655 ;
        RECT -217.845 -179.825 -217.675 -179.655 ;
        RECT -207.925 -178.905 -207.755 -178.735 ;
        RECT -201.545 -178.905 -201.375 -178.735 ;
        RECT -207.925 -179.365 -207.755 -179.195 ;
        RECT -201.545 -179.365 -201.375 -179.195 ;
        RECT -209.695 -179.635 -209.525 -179.465 ;
        RECT -211.465 -179.825 -211.295 -179.655 ;
        RECT -207.925 -179.825 -207.755 -179.655 ;
        RECT -198.005 -178.905 -197.835 -178.735 ;
        RECT -191.625 -178.905 -191.455 -178.735 ;
        RECT -198.005 -179.365 -197.835 -179.195 ;
        RECT -191.625 -179.365 -191.455 -179.195 ;
        RECT -199.775 -179.635 -199.605 -179.465 ;
        RECT -201.545 -179.825 -201.375 -179.655 ;
        RECT -198.005 -179.825 -197.835 -179.655 ;
        RECT -188.085 -178.905 -187.915 -178.735 ;
        RECT -181.705 -178.905 -181.535 -178.735 ;
        RECT -188.085 -179.365 -187.915 -179.195 ;
        RECT -181.705 -179.365 -181.535 -179.195 ;
        RECT -189.855 -179.635 -189.685 -179.465 ;
        RECT -191.625 -179.825 -191.455 -179.655 ;
        RECT -188.085 -179.825 -187.915 -179.655 ;
        RECT -178.165 -178.905 -177.995 -178.735 ;
        RECT -171.785 -178.905 -171.615 -178.735 ;
        RECT -178.165 -179.365 -177.995 -179.195 ;
        RECT -171.785 -179.365 -171.615 -179.195 ;
        RECT -179.935 -179.635 -179.765 -179.465 ;
        RECT -181.705 -179.825 -181.535 -179.655 ;
        RECT -178.165 -179.825 -177.995 -179.655 ;
        RECT -168.245 -178.905 -168.075 -178.735 ;
        RECT -161.865 -178.905 -161.695 -178.735 ;
        RECT -168.245 -179.365 -168.075 -179.195 ;
        RECT -161.865 -179.365 -161.695 -179.195 ;
        RECT -170.015 -179.635 -169.845 -179.465 ;
        RECT -171.785 -179.825 -171.615 -179.655 ;
        RECT -168.245 -179.825 -168.075 -179.655 ;
        RECT -158.325 -178.905 -158.155 -178.735 ;
        RECT -151.945 -178.905 -151.775 -178.735 ;
        RECT -158.325 -179.365 -158.155 -179.195 ;
        RECT -151.945 -179.365 -151.775 -179.195 ;
        RECT -160.095 -179.635 -159.925 -179.465 ;
        RECT -161.865 -179.825 -161.695 -179.655 ;
        RECT -158.325 -179.825 -158.155 -179.655 ;
        RECT -148.405 -178.905 -148.235 -178.735 ;
        RECT -142.025 -178.905 -141.855 -178.735 ;
        RECT -148.405 -179.365 -148.235 -179.195 ;
        RECT -142.025 -179.365 -141.855 -179.195 ;
        RECT -150.175 -179.635 -150.005 -179.465 ;
        RECT -151.945 -179.825 -151.775 -179.655 ;
        RECT -148.405 -179.825 -148.235 -179.655 ;
        RECT -138.485 -178.905 -138.315 -178.735 ;
        RECT -132.105 -178.905 -131.935 -178.735 ;
        RECT -138.485 -179.365 -138.315 -179.195 ;
        RECT -132.105 -179.365 -131.935 -179.195 ;
        RECT -140.255 -179.635 -140.085 -179.465 ;
        RECT -142.025 -179.825 -141.855 -179.655 ;
        RECT -138.485 -179.825 -138.315 -179.655 ;
        RECT -128.565 -178.905 -128.395 -178.735 ;
        RECT -122.185 -178.905 -122.015 -178.735 ;
        RECT -128.565 -179.365 -128.395 -179.195 ;
        RECT -122.185 -179.365 -122.015 -179.195 ;
        RECT -130.335 -179.635 -130.165 -179.465 ;
        RECT -132.105 -179.825 -131.935 -179.655 ;
        RECT -128.565 -179.825 -128.395 -179.655 ;
        RECT -118.645 -178.905 -118.475 -178.735 ;
        RECT -112.265 -178.905 -112.095 -178.735 ;
        RECT -118.645 -179.365 -118.475 -179.195 ;
        RECT -112.265 -179.365 -112.095 -179.195 ;
        RECT -120.415 -179.635 -120.245 -179.465 ;
        RECT -122.185 -179.825 -122.015 -179.655 ;
        RECT -118.645 -179.825 -118.475 -179.655 ;
        RECT -108.725 -178.905 -108.555 -178.735 ;
        RECT -102.345 -178.905 -102.175 -178.735 ;
        RECT -108.725 -179.365 -108.555 -179.195 ;
        RECT -102.345 -179.365 -102.175 -179.195 ;
        RECT -110.495 -179.635 -110.325 -179.465 ;
        RECT -112.265 -179.825 -112.095 -179.655 ;
        RECT -108.725 -179.825 -108.555 -179.655 ;
        RECT -98.805 -178.905 -98.635 -178.735 ;
        RECT -92.425 -178.905 -92.255 -178.735 ;
        RECT -98.805 -179.365 -98.635 -179.195 ;
        RECT -92.425 -179.365 -92.255 -179.195 ;
        RECT -100.575 -179.635 -100.405 -179.465 ;
        RECT -102.345 -179.825 -102.175 -179.655 ;
        RECT -98.805 -179.825 -98.635 -179.655 ;
        RECT -88.885 -178.905 -88.715 -178.735 ;
        RECT -82.505 -178.905 -82.335 -178.735 ;
        RECT -88.885 -179.365 -88.715 -179.195 ;
        RECT -82.505 -179.365 -82.335 -179.195 ;
        RECT -90.655 -179.635 -90.485 -179.465 ;
        RECT -92.425 -179.825 -92.255 -179.655 ;
        RECT -88.885 -179.825 -88.715 -179.655 ;
        RECT -78.965 -178.905 -78.795 -178.735 ;
        RECT -72.585 -178.905 -72.415 -178.735 ;
        RECT -78.965 -179.365 -78.795 -179.195 ;
        RECT -72.585 -179.365 -72.415 -179.195 ;
        RECT -80.735 -179.635 -80.565 -179.465 ;
        RECT -82.505 -179.825 -82.335 -179.655 ;
        RECT -78.965 -179.825 -78.795 -179.655 ;
        RECT -69.045 -178.905 -68.875 -178.735 ;
        RECT -62.665 -178.905 -62.495 -178.735 ;
        RECT -69.045 -179.365 -68.875 -179.195 ;
        RECT -62.665 -179.365 -62.495 -179.195 ;
        RECT -70.815 -179.635 -70.645 -179.465 ;
        RECT -72.585 -179.825 -72.415 -179.655 ;
        RECT -69.045 -179.825 -68.875 -179.655 ;
        RECT -59.125 -178.905 -58.955 -178.735 ;
        RECT -52.745 -178.905 -52.575 -178.735 ;
        RECT -59.125 -179.365 -58.955 -179.195 ;
        RECT -52.745 -179.365 -52.575 -179.195 ;
        RECT -60.895 -179.635 -60.725 -179.465 ;
        RECT -62.665 -179.825 -62.495 -179.655 ;
        RECT -59.125 -179.825 -58.955 -179.655 ;
        RECT -49.205 -178.905 -49.035 -178.735 ;
        RECT -42.825 -178.905 -42.655 -178.735 ;
        RECT -49.205 -179.365 -49.035 -179.195 ;
        RECT -42.825 -179.365 -42.655 -179.195 ;
        RECT -50.975 -179.635 -50.805 -179.465 ;
        RECT -52.745 -179.825 -52.575 -179.655 ;
        RECT -49.205 -179.825 -49.035 -179.655 ;
        RECT -39.285 -178.905 -39.115 -178.735 ;
        RECT -32.905 -178.905 -32.735 -178.735 ;
        RECT -39.285 -179.365 -39.115 -179.195 ;
        RECT -32.905 -179.365 -32.735 -179.195 ;
        RECT -41.055 -179.635 -40.885 -179.465 ;
        RECT -42.825 -179.825 -42.655 -179.655 ;
        RECT -39.285 -179.825 -39.115 -179.655 ;
        RECT -29.365 -178.905 -29.195 -178.735 ;
        RECT -22.985 -178.905 -22.815 -178.735 ;
        RECT -29.365 -179.365 -29.195 -179.195 ;
        RECT -22.985 -179.365 -22.815 -179.195 ;
        RECT -31.135 -179.635 -30.965 -179.465 ;
        RECT -32.905 -179.825 -32.735 -179.655 ;
        RECT -29.365 -179.825 -29.195 -179.655 ;
        RECT -19.445 -178.905 -19.275 -178.735 ;
        RECT -13.065 -178.905 -12.895 -178.735 ;
        RECT -19.445 -179.365 -19.275 -179.195 ;
        RECT -13.065 -179.365 -12.895 -179.195 ;
        RECT -21.215 -179.635 -21.045 -179.465 ;
        RECT -22.985 -179.825 -22.815 -179.655 ;
        RECT -19.445 -179.825 -19.275 -179.655 ;
        RECT -9.525 -178.905 -9.355 -178.735 ;
        RECT -3.145 -178.905 -2.975 -178.735 ;
        RECT -9.525 -179.365 -9.355 -179.195 ;
        RECT -3.145 -179.365 -2.975 -179.195 ;
        RECT -11.295 -179.635 -11.125 -179.465 ;
        RECT -13.065 -179.825 -12.895 -179.655 ;
        RECT -9.525 -179.825 -9.355 -179.655 ;
        RECT 0.395 -178.905 0.565 -178.735 ;
        RECT 6.775 -178.905 6.945 -178.735 ;
        RECT 0.395 -179.365 0.565 -179.195 ;
        RECT 6.775 -179.365 6.945 -179.195 ;
        RECT -1.375 -179.635 -1.205 -179.465 ;
        RECT -3.145 -179.825 -2.975 -179.655 ;
        RECT 0.395 -179.825 0.565 -179.655 ;
        RECT 10.315 -178.905 10.485 -178.735 ;
        RECT 16.695 -178.905 16.865 -178.735 ;
        RECT 10.315 -179.365 10.485 -179.195 ;
        RECT 16.695 -179.365 16.865 -179.195 ;
        RECT 8.545 -179.635 8.715 -179.465 ;
        RECT 6.775 -179.825 6.945 -179.655 ;
        RECT 10.315 -179.825 10.485 -179.655 ;
        RECT 20.235 -178.905 20.405 -178.735 ;
        RECT 20.235 -179.365 20.405 -179.195 ;
        RECT 18.465 -179.635 18.635 -179.465 ;
        RECT 16.695 -179.825 16.865 -179.655 ;
        RECT 20.235 -179.825 20.405 -179.655 ;
      LAYER met1 ;
        RECT -288.280 93.760 -284.260 95.140 ;
        RECT -278.360 93.760 -274.340 95.140 ;
        RECT -268.440 93.760 -264.420 95.140 ;
        RECT -258.520 93.760 -254.500 95.140 ;
        RECT -248.600 93.760 -244.580 95.140 ;
        RECT -238.680 93.760 -234.660 95.140 ;
        RECT -228.760 93.760 -224.740 95.140 ;
        RECT -218.840 93.760 -214.820 95.140 ;
        RECT -208.920 93.760 -204.900 95.140 ;
        RECT -199.000 93.760 -194.980 95.140 ;
        RECT -189.080 93.760 -185.060 95.140 ;
        RECT -179.160 93.760 -175.140 95.140 ;
        RECT -169.240 93.760 -165.220 95.140 ;
        RECT -159.320 93.760 -155.300 95.140 ;
        RECT -149.400 93.760 -145.380 95.140 ;
        RECT -139.480 93.760 -135.460 95.140 ;
        RECT -129.560 93.760 -125.540 95.140 ;
        RECT -119.640 93.760 -115.620 95.140 ;
        RECT -109.720 93.760 -105.700 95.140 ;
        RECT -99.800 93.760 -95.780 95.140 ;
        RECT -89.880 93.760 -85.860 95.140 ;
        RECT -79.960 93.760 -75.940 95.140 ;
        RECT -70.040 93.760 -66.020 95.140 ;
        RECT -60.120 93.760 -56.100 95.140 ;
        RECT -50.200 93.760 -46.180 95.140 ;
        RECT -40.280 93.760 -36.260 95.140 ;
        RECT -30.360 93.760 -26.340 95.140 ;
        RECT -20.440 93.760 -16.420 95.140 ;
        RECT -10.520 93.760 -6.500 95.140 ;
        RECT -0.600 93.760 3.420 95.140 ;
        RECT 9.320 93.760 13.340 95.140 ;
        RECT 19.240 93.760 23.260 95.140 ;
        RECT -282.920 93.090 -279.700 93.570 ;
        RECT -273.000 93.090 -269.780 93.570 ;
        RECT -263.080 93.090 -259.860 93.570 ;
        RECT -253.160 93.090 -249.940 93.570 ;
        RECT -243.240 93.090 -240.020 93.570 ;
        RECT -233.320 93.090 -230.100 93.570 ;
        RECT -223.400 93.090 -220.180 93.570 ;
        RECT -213.480 93.090 -210.260 93.570 ;
        RECT -203.560 93.090 -200.340 93.570 ;
        RECT -193.640 93.090 -190.420 93.570 ;
        RECT -183.720 93.090 -180.500 93.570 ;
        RECT -173.800 93.090 -170.580 93.570 ;
        RECT -163.880 93.090 -160.660 93.570 ;
        RECT -153.960 93.090 -150.740 93.570 ;
        RECT -144.040 93.090 -140.820 93.570 ;
        RECT -134.120 93.090 -130.900 93.570 ;
        RECT -124.200 93.090 -120.980 93.570 ;
        RECT -114.280 93.090 -111.060 93.570 ;
        RECT -104.360 93.090 -101.140 93.570 ;
        RECT -94.440 93.090 -91.220 93.570 ;
        RECT -84.520 93.090 -81.300 93.570 ;
        RECT -74.600 93.090 -71.380 93.570 ;
        RECT -64.680 93.090 -61.460 93.570 ;
        RECT -54.760 93.090 -51.540 93.570 ;
        RECT -44.840 93.090 -41.620 93.570 ;
        RECT -34.920 93.090 -31.700 93.570 ;
        RECT -25.000 93.090 -21.780 93.570 ;
        RECT -15.080 93.090 -11.860 93.570 ;
        RECT -5.160 93.090 -1.940 93.570 ;
        RECT 4.760 93.090 7.980 93.570 ;
        RECT 14.680 93.090 17.900 93.570 ;
        RECT -287.880 90.370 -284.660 90.850 ;
        RECT -277.960 90.370 -274.740 90.850 ;
        RECT -268.040 90.370 -264.820 90.850 ;
        RECT -258.120 90.370 -254.900 90.850 ;
        RECT -248.200 90.370 -244.980 90.850 ;
        RECT -238.280 90.370 -235.060 90.850 ;
        RECT -228.360 90.370 -225.140 90.850 ;
        RECT -218.440 90.370 -215.220 90.850 ;
        RECT -208.520 90.370 -205.300 90.850 ;
        RECT -198.600 90.370 -195.380 90.850 ;
        RECT -188.680 90.370 -185.460 90.850 ;
        RECT -178.760 90.370 -175.540 90.850 ;
        RECT -168.840 90.370 -165.620 90.850 ;
        RECT -158.920 90.370 -155.700 90.850 ;
        RECT -149.000 90.370 -145.780 90.850 ;
        RECT -139.080 90.370 -135.860 90.850 ;
        RECT -129.160 90.370 -125.940 90.850 ;
        RECT -119.240 90.370 -116.020 90.850 ;
        RECT -109.320 90.370 -106.100 90.850 ;
        RECT -99.400 90.370 -96.180 90.850 ;
        RECT -89.480 90.370 -86.260 90.850 ;
        RECT -79.560 90.370 -76.340 90.850 ;
        RECT -69.640 90.370 -66.420 90.850 ;
        RECT -59.720 90.370 -56.500 90.850 ;
        RECT -49.800 90.370 -46.580 90.850 ;
        RECT -39.880 90.370 -36.660 90.850 ;
        RECT -29.960 90.370 -26.740 90.850 ;
        RECT -20.040 90.370 -16.820 90.850 ;
        RECT -10.120 90.370 -6.900 90.850 ;
        RECT -0.200 90.370 3.020 90.850 ;
        RECT 9.720 90.370 12.940 90.850 ;
        RECT 19.640 90.370 22.860 90.850 ;
        RECT -283.320 88.800 -279.300 90.180 ;
        RECT -273.400 88.800 -269.380 90.180 ;
        RECT -263.480 88.800 -259.460 90.180 ;
        RECT -253.560 88.800 -249.540 90.180 ;
        RECT -243.640 88.800 -239.620 90.180 ;
        RECT -233.720 88.800 -229.700 90.180 ;
        RECT -223.800 88.800 -219.780 90.180 ;
        RECT -213.880 88.800 -209.860 90.180 ;
        RECT -203.960 88.800 -199.940 90.180 ;
        RECT -194.040 88.800 -190.020 90.180 ;
        RECT -184.120 88.800 -180.100 90.180 ;
        RECT -174.200 88.800 -170.180 90.180 ;
        RECT -164.280 88.800 -160.260 90.180 ;
        RECT -154.360 88.800 -150.340 90.180 ;
        RECT -144.440 88.800 -140.420 90.180 ;
        RECT -134.520 88.800 -130.500 90.180 ;
        RECT -124.600 88.800 -120.580 90.180 ;
        RECT -114.680 88.800 -110.660 90.180 ;
        RECT -104.760 88.800 -100.740 90.180 ;
        RECT -94.840 88.800 -90.820 90.180 ;
        RECT -84.920 88.800 -80.900 90.180 ;
        RECT -75.000 88.800 -70.980 90.180 ;
        RECT -65.080 88.800 -61.060 90.180 ;
        RECT -55.160 88.800 -51.140 90.180 ;
        RECT -45.240 88.800 -41.220 90.180 ;
        RECT -35.320 88.800 -31.300 90.180 ;
        RECT -25.400 88.800 -21.380 90.180 ;
        RECT -15.480 88.800 -11.460 90.180 ;
        RECT -5.560 88.800 -1.540 90.180 ;
        RECT 4.360 88.800 8.380 90.180 ;
        RECT 14.280 88.800 18.300 90.180 ;
        RECT -288.030 6.050 -284.010 7.430 ;
        RECT -278.110 6.050 -274.090 7.430 ;
        RECT -268.190 6.050 -264.170 7.430 ;
        RECT -258.270 6.050 -254.250 7.430 ;
        RECT -248.350 6.050 -244.330 7.430 ;
        RECT -238.430 6.050 -234.410 7.430 ;
        RECT -228.510 6.050 -224.490 7.430 ;
        RECT -218.590 6.050 -214.570 7.430 ;
        RECT -208.670 6.050 -204.650 7.430 ;
        RECT -198.750 6.050 -194.730 7.430 ;
        RECT -188.830 6.050 -184.810 7.430 ;
        RECT -178.910 6.050 -174.890 7.430 ;
        RECT -168.990 6.050 -164.970 7.430 ;
        RECT -159.070 6.050 -155.050 7.430 ;
        RECT -149.150 6.050 -145.130 7.430 ;
        RECT -139.230 6.050 -135.210 7.430 ;
        RECT -129.310 6.050 -125.290 7.430 ;
        RECT -119.390 6.050 -115.370 7.430 ;
        RECT -109.470 6.050 -105.450 7.430 ;
        RECT -99.550 6.050 -95.530 7.430 ;
        RECT -89.630 6.050 -85.610 7.430 ;
        RECT -79.710 6.050 -75.690 7.430 ;
        RECT -69.790 6.050 -65.770 7.430 ;
        RECT -59.870 6.050 -55.850 7.430 ;
        RECT -49.950 6.050 -45.930 7.430 ;
        RECT -40.030 6.050 -36.010 7.430 ;
        RECT -30.110 6.050 -26.090 7.430 ;
        RECT -20.190 6.050 -16.170 7.430 ;
        RECT -10.270 6.050 -6.250 7.430 ;
        RECT -0.350 6.050 3.670 7.430 ;
        RECT 9.570 6.050 13.590 7.430 ;
        RECT 19.490 6.050 23.510 7.430 ;
        RECT -282.670 5.380 -279.450 5.860 ;
        RECT -272.750 5.380 -269.530 5.860 ;
        RECT -262.830 5.380 -259.610 5.860 ;
        RECT -252.910 5.380 -249.690 5.860 ;
        RECT -242.990 5.380 -239.770 5.860 ;
        RECT -233.070 5.380 -229.850 5.860 ;
        RECT -223.150 5.380 -219.930 5.860 ;
        RECT -213.230 5.380 -210.010 5.860 ;
        RECT -203.310 5.380 -200.090 5.860 ;
        RECT -193.390 5.380 -190.170 5.860 ;
        RECT -183.470 5.380 -180.250 5.860 ;
        RECT -173.550 5.380 -170.330 5.860 ;
        RECT -163.630 5.380 -160.410 5.860 ;
        RECT -153.710 5.380 -150.490 5.860 ;
        RECT -143.790 5.380 -140.570 5.860 ;
        RECT -133.870 5.380 -130.650 5.860 ;
        RECT -123.950 5.380 -120.730 5.860 ;
        RECT -114.030 5.380 -110.810 5.860 ;
        RECT -104.110 5.380 -100.890 5.860 ;
        RECT -94.190 5.380 -90.970 5.860 ;
        RECT -84.270 5.380 -81.050 5.860 ;
        RECT -74.350 5.380 -71.130 5.860 ;
        RECT -64.430 5.380 -61.210 5.860 ;
        RECT -54.510 5.380 -51.290 5.860 ;
        RECT -44.590 5.380 -41.370 5.860 ;
        RECT -34.670 5.380 -31.450 5.860 ;
        RECT -24.750 5.380 -21.530 5.860 ;
        RECT -14.830 5.380 -11.610 5.860 ;
        RECT -4.910 5.380 -1.690 5.860 ;
        RECT 5.010 5.380 8.230 5.860 ;
        RECT 14.930 5.380 18.150 5.860 ;
        RECT -287.630 2.660 -284.410 3.140 ;
        RECT -277.710 2.660 -274.490 3.140 ;
        RECT -267.790 2.660 -264.570 3.140 ;
        RECT -257.870 2.660 -254.650 3.140 ;
        RECT -247.950 2.660 -244.730 3.140 ;
        RECT -238.030 2.660 -234.810 3.140 ;
        RECT -228.110 2.660 -224.890 3.140 ;
        RECT -218.190 2.660 -214.970 3.140 ;
        RECT -208.270 2.660 -205.050 3.140 ;
        RECT -198.350 2.660 -195.130 3.140 ;
        RECT -188.430 2.660 -185.210 3.140 ;
        RECT -178.510 2.660 -175.290 3.140 ;
        RECT -168.590 2.660 -165.370 3.140 ;
        RECT -158.670 2.660 -155.450 3.140 ;
        RECT -148.750 2.660 -145.530 3.140 ;
        RECT -138.830 2.660 -135.610 3.140 ;
        RECT -128.910 2.660 -125.690 3.140 ;
        RECT -118.990 2.660 -115.770 3.140 ;
        RECT -109.070 2.660 -105.850 3.140 ;
        RECT -99.150 2.660 -95.930 3.140 ;
        RECT -89.230 2.660 -86.010 3.140 ;
        RECT -79.310 2.660 -76.090 3.140 ;
        RECT -69.390 2.660 -66.170 3.140 ;
        RECT -59.470 2.660 -56.250 3.140 ;
        RECT -49.550 2.660 -46.330 3.140 ;
        RECT -39.630 2.660 -36.410 3.140 ;
        RECT -29.710 2.660 -26.490 3.140 ;
        RECT -19.790 2.660 -16.570 3.140 ;
        RECT -9.870 2.660 -6.650 3.140 ;
        RECT 0.050 2.660 3.270 3.140 ;
        RECT 9.970 2.660 13.190 3.140 ;
        RECT 19.890 2.660 23.110 3.140 ;
        RECT -283.070 1.090 -279.050 2.470 ;
        RECT -273.150 1.090 -269.130 2.470 ;
        RECT -263.230 1.090 -259.210 2.470 ;
        RECT -253.310 1.090 -249.290 2.470 ;
        RECT -243.390 1.090 -239.370 2.470 ;
        RECT -233.470 1.090 -229.450 2.470 ;
        RECT -223.550 1.090 -219.530 2.470 ;
        RECT -213.630 1.090 -209.610 2.470 ;
        RECT -203.710 1.090 -199.690 2.470 ;
        RECT -193.790 1.090 -189.770 2.470 ;
        RECT -183.870 1.090 -179.850 2.470 ;
        RECT -173.950 1.090 -169.930 2.470 ;
        RECT -164.030 1.090 -160.010 2.470 ;
        RECT -154.110 1.090 -150.090 2.470 ;
        RECT -144.190 1.090 -140.170 2.470 ;
        RECT -134.270 1.090 -130.250 2.470 ;
        RECT -124.350 1.090 -120.330 2.470 ;
        RECT -114.430 1.090 -110.410 2.470 ;
        RECT -104.510 1.090 -100.490 2.470 ;
        RECT -94.590 1.090 -90.570 2.470 ;
        RECT -84.670 1.090 -80.650 2.470 ;
        RECT -74.750 1.090 -70.730 2.470 ;
        RECT -64.830 1.090 -60.810 2.470 ;
        RECT -54.910 1.090 -50.890 2.470 ;
        RECT -44.990 1.090 -40.970 2.470 ;
        RECT -35.070 1.090 -31.050 2.470 ;
        RECT -25.150 1.090 -21.130 2.470 ;
        RECT -15.230 1.090 -11.210 2.470 ;
        RECT -5.310 1.090 -1.290 2.470 ;
        RECT 4.610 1.090 8.630 2.470 ;
        RECT 14.530 1.090 18.550 2.470 ;
        RECT -286.270 -87.300 -282.250 -85.920 ;
        RECT -276.350 -87.300 -272.330 -85.920 ;
        RECT -266.430 -87.300 -262.410 -85.920 ;
        RECT -256.510 -87.300 -252.490 -85.920 ;
        RECT -246.590 -87.300 -242.570 -85.920 ;
        RECT -236.670 -87.300 -232.650 -85.920 ;
        RECT -226.750 -87.300 -222.730 -85.920 ;
        RECT -216.830 -87.300 -212.810 -85.920 ;
        RECT -206.910 -87.300 -202.890 -85.920 ;
        RECT -196.990 -87.300 -192.970 -85.920 ;
        RECT -187.070 -87.300 -183.050 -85.920 ;
        RECT -177.150 -87.300 -173.130 -85.920 ;
        RECT -167.230 -87.300 -163.210 -85.920 ;
        RECT -157.310 -87.300 -153.290 -85.920 ;
        RECT -147.390 -87.300 -143.370 -85.920 ;
        RECT -137.470 -87.300 -133.450 -85.920 ;
        RECT -127.550 -87.300 -123.530 -85.920 ;
        RECT -117.630 -87.300 -113.610 -85.920 ;
        RECT -107.710 -87.300 -103.690 -85.920 ;
        RECT -97.790 -87.300 -93.770 -85.920 ;
        RECT -87.870 -87.300 -83.850 -85.920 ;
        RECT -77.950 -87.300 -73.930 -85.920 ;
        RECT -68.030 -87.300 -64.010 -85.920 ;
        RECT -58.110 -87.300 -54.090 -85.920 ;
        RECT -48.190 -87.300 -44.170 -85.920 ;
        RECT -38.270 -87.300 -34.250 -85.920 ;
        RECT -28.350 -87.300 -24.330 -85.920 ;
        RECT -18.430 -87.300 -14.410 -85.920 ;
        RECT -8.510 -87.300 -4.490 -85.920 ;
        RECT 1.410 -87.300 5.430 -85.920 ;
        RECT 11.330 -87.300 15.350 -85.920 ;
        RECT 21.250 -87.300 25.270 -85.920 ;
        RECT -280.910 -87.970 -277.690 -87.490 ;
        RECT -270.990 -87.970 -267.770 -87.490 ;
        RECT -261.070 -87.970 -257.850 -87.490 ;
        RECT -251.150 -87.970 -247.930 -87.490 ;
        RECT -241.230 -87.970 -238.010 -87.490 ;
        RECT -231.310 -87.970 -228.090 -87.490 ;
        RECT -221.390 -87.970 -218.170 -87.490 ;
        RECT -211.470 -87.970 -208.250 -87.490 ;
        RECT -201.550 -87.970 -198.330 -87.490 ;
        RECT -191.630 -87.970 -188.410 -87.490 ;
        RECT -181.710 -87.970 -178.490 -87.490 ;
        RECT -171.790 -87.970 -168.570 -87.490 ;
        RECT -161.870 -87.970 -158.650 -87.490 ;
        RECT -151.950 -87.970 -148.730 -87.490 ;
        RECT -142.030 -87.970 -138.810 -87.490 ;
        RECT -132.110 -87.970 -128.890 -87.490 ;
        RECT -122.190 -87.970 -118.970 -87.490 ;
        RECT -112.270 -87.970 -109.050 -87.490 ;
        RECT -102.350 -87.970 -99.130 -87.490 ;
        RECT -92.430 -87.970 -89.210 -87.490 ;
        RECT -82.510 -87.970 -79.290 -87.490 ;
        RECT -72.590 -87.970 -69.370 -87.490 ;
        RECT -62.670 -87.970 -59.450 -87.490 ;
        RECT -52.750 -87.970 -49.530 -87.490 ;
        RECT -42.830 -87.970 -39.610 -87.490 ;
        RECT -32.910 -87.970 -29.690 -87.490 ;
        RECT -22.990 -87.970 -19.770 -87.490 ;
        RECT -13.070 -87.970 -9.850 -87.490 ;
        RECT -3.150 -87.970 0.070 -87.490 ;
        RECT 6.770 -87.970 9.990 -87.490 ;
        RECT 16.690 -87.970 19.910 -87.490 ;
        RECT -285.870 -90.690 -282.650 -90.210 ;
        RECT -275.950 -90.690 -272.730 -90.210 ;
        RECT -266.030 -90.690 -262.810 -90.210 ;
        RECT -256.110 -90.690 -252.890 -90.210 ;
        RECT -246.190 -90.690 -242.970 -90.210 ;
        RECT -236.270 -90.690 -233.050 -90.210 ;
        RECT -226.350 -90.690 -223.130 -90.210 ;
        RECT -216.430 -90.690 -213.210 -90.210 ;
        RECT -206.510 -90.690 -203.290 -90.210 ;
        RECT -196.590 -90.690 -193.370 -90.210 ;
        RECT -186.670 -90.690 -183.450 -90.210 ;
        RECT -176.750 -90.690 -173.530 -90.210 ;
        RECT -166.830 -90.690 -163.610 -90.210 ;
        RECT -156.910 -90.690 -153.690 -90.210 ;
        RECT -146.990 -90.690 -143.770 -90.210 ;
        RECT -137.070 -90.690 -133.850 -90.210 ;
        RECT -127.150 -90.690 -123.930 -90.210 ;
        RECT -117.230 -90.690 -114.010 -90.210 ;
        RECT -107.310 -90.690 -104.090 -90.210 ;
        RECT -97.390 -90.690 -94.170 -90.210 ;
        RECT -87.470 -90.690 -84.250 -90.210 ;
        RECT -77.550 -90.690 -74.330 -90.210 ;
        RECT -67.630 -90.690 -64.410 -90.210 ;
        RECT -57.710 -90.690 -54.490 -90.210 ;
        RECT -47.790 -90.690 -44.570 -90.210 ;
        RECT -37.870 -90.690 -34.650 -90.210 ;
        RECT -27.950 -90.690 -24.730 -90.210 ;
        RECT -18.030 -90.690 -14.810 -90.210 ;
        RECT -8.110 -90.690 -4.890 -90.210 ;
        RECT 1.810 -90.690 5.030 -90.210 ;
        RECT 11.730 -90.690 14.950 -90.210 ;
        RECT 21.650 -90.690 24.870 -90.210 ;
        RECT -281.310 -92.260 -277.290 -90.880 ;
        RECT -271.390 -92.260 -267.370 -90.880 ;
        RECT -261.470 -92.260 -257.450 -90.880 ;
        RECT -251.550 -92.260 -247.530 -90.880 ;
        RECT -241.630 -92.260 -237.610 -90.880 ;
        RECT -231.710 -92.260 -227.690 -90.880 ;
        RECT -221.790 -92.260 -217.770 -90.880 ;
        RECT -211.870 -92.260 -207.850 -90.880 ;
        RECT -201.950 -92.260 -197.930 -90.880 ;
        RECT -192.030 -92.260 -188.010 -90.880 ;
        RECT -182.110 -92.260 -178.090 -90.880 ;
        RECT -172.190 -92.260 -168.170 -90.880 ;
        RECT -162.270 -92.260 -158.250 -90.880 ;
        RECT -152.350 -92.260 -148.330 -90.880 ;
        RECT -142.430 -92.260 -138.410 -90.880 ;
        RECT -132.510 -92.260 -128.490 -90.880 ;
        RECT -122.590 -92.260 -118.570 -90.880 ;
        RECT -112.670 -92.260 -108.650 -90.880 ;
        RECT -102.750 -92.260 -98.730 -90.880 ;
        RECT -92.830 -92.260 -88.810 -90.880 ;
        RECT -82.910 -92.260 -78.890 -90.880 ;
        RECT -72.990 -92.260 -68.970 -90.880 ;
        RECT -63.070 -92.260 -59.050 -90.880 ;
        RECT -53.150 -92.260 -49.130 -90.880 ;
        RECT -43.230 -92.260 -39.210 -90.880 ;
        RECT -33.310 -92.260 -29.290 -90.880 ;
        RECT -23.390 -92.260 -19.370 -90.880 ;
        RECT -13.470 -92.260 -9.450 -90.880 ;
        RECT -3.550 -92.260 0.470 -90.880 ;
        RECT 6.370 -92.260 10.390 -90.880 ;
        RECT 16.290 -92.260 20.310 -90.880 ;
        RECT -286.020 -175.010 -282.000 -173.630 ;
        RECT -276.100 -175.010 -272.080 -173.630 ;
        RECT -266.180 -175.010 -262.160 -173.630 ;
        RECT -256.260 -175.010 -252.240 -173.630 ;
        RECT -246.340 -175.010 -242.320 -173.630 ;
        RECT -236.420 -175.010 -232.400 -173.630 ;
        RECT -226.500 -175.010 -222.480 -173.630 ;
        RECT -216.580 -175.010 -212.560 -173.630 ;
        RECT -206.660 -175.010 -202.640 -173.630 ;
        RECT -196.740 -175.010 -192.720 -173.630 ;
        RECT -186.820 -175.010 -182.800 -173.630 ;
        RECT -176.900 -175.010 -172.880 -173.630 ;
        RECT -166.980 -175.010 -162.960 -173.630 ;
        RECT -157.060 -175.010 -153.040 -173.630 ;
        RECT -147.140 -175.010 -143.120 -173.630 ;
        RECT -137.220 -175.010 -133.200 -173.630 ;
        RECT -127.300 -175.010 -123.280 -173.630 ;
        RECT -117.380 -175.010 -113.360 -173.630 ;
        RECT -107.460 -175.010 -103.440 -173.630 ;
        RECT -97.540 -175.010 -93.520 -173.630 ;
        RECT -87.620 -175.010 -83.600 -173.630 ;
        RECT -77.700 -175.010 -73.680 -173.630 ;
        RECT -67.780 -175.010 -63.760 -173.630 ;
        RECT -57.860 -175.010 -53.840 -173.630 ;
        RECT -47.940 -175.010 -43.920 -173.630 ;
        RECT -38.020 -175.010 -34.000 -173.630 ;
        RECT -28.100 -175.010 -24.080 -173.630 ;
        RECT -18.180 -175.010 -14.160 -173.630 ;
        RECT -8.260 -175.010 -4.240 -173.630 ;
        RECT 1.660 -175.010 5.680 -173.630 ;
        RECT 11.580 -175.010 15.600 -173.630 ;
        RECT 21.500 -175.010 25.520 -173.630 ;
        RECT -280.660 -175.680 -277.440 -175.200 ;
        RECT -270.740 -175.680 -267.520 -175.200 ;
        RECT -260.820 -175.680 -257.600 -175.200 ;
        RECT -250.900 -175.680 -247.680 -175.200 ;
        RECT -240.980 -175.680 -237.760 -175.200 ;
        RECT -231.060 -175.680 -227.840 -175.200 ;
        RECT -221.140 -175.680 -217.920 -175.200 ;
        RECT -211.220 -175.680 -208.000 -175.200 ;
        RECT -201.300 -175.680 -198.080 -175.200 ;
        RECT -191.380 -175.680 -188.160 -175.200 ;
        RECT -181.460 -175.680 -178.240 -175.200 ;
        RECT -171.540 -175.680 -168.320 -175.200 ;
        RECT -161.620 -175.680 -158.400 -175.200 ;
        RECT -151.700 -175.680 -148.480 -175.200 ;
        RECT -141.780 -175.680 -138.560 -175.200 ;
        RECT -131.860 -175.680 -128.640 -175.200 ;
        RECT -121.940 -175.680 -118.720 -175.200 ;
        RECT -112.020 -175.680 -108.800 -175.200 ;
        RECT -102.100 -175.680 -98.880 -175.200 ;
        RECT -92.180 -175.680 -88.960 -175.200 ;
        RECT -82.260 -175.680 -79.040 -175.200 ;
        RECT -72.340 -175.680 -69.120 -175.200 ;
        RECT -62.420 -175.680 -59.200 -175.200 ;
        RECT -52.500 -175.680 -49.280 -175.200 ;
        RECT -42.580 -175.680 -39.360 -175.200 ;
        RECT -32.660 -175.680 -29.440 -175.200 ;
        RECT -22.740 -175.680 -19.520 -175.200 ;
        RECT -12.820 -175.680 -9.600 -175.200 ;
        RECT -2.900 -175.680 0.320 -175.200 ;
        RECT 7.020 -175.680 10.240 -175.200 ;
        RECT 16.940 -175.680 20.160 -175.200 ;
        RECT -285.620 -178.400 -282.400 -177.920 ;
        RECT -275.700 -178.400 -272.480 -177.920 ;
        RECT -265.780 -178.400 -262.560 -177.920 ;
        RECT -255.860 -178.400 -252.640 -177.920 ;
        RECT -245.940 -178.400 -242.720 -177.920 ;
        RECT -236.020 -178.400 -232.800 -177.920 ;
        RECT -226.100 -178.400 -222.880 -177.920 ;
        RECT -216.180 -178.400 -212.960 -177.920 ;
        RECT -206.260 -178.400 -203.040 -177.920 ;
        RECT -196.340 -178.400 -193.120 -177.920 ;
        RECT -186.420 -178.400 -183.200 -177.920 ;
        RECT -176.500 -178.400 -173.280 -177.920 ;
        RECT -166.580 -178.400 -163.360 -177.920 ;
        RECT -156.660 -178.400 -153.440 -177.920 ;
        RECT -146.740 -178.400 -143.520 -177.920 ;
        RECT -136.820 -178.400 -133.600 -177.920 ;
        RECT -126.900 -178.400 -123.680 -177.920 ;
        RECT -116.980 -178.400 -113.760 -177.920 ;
        RECT -107.060 -178.400 -103.840 -177.920 ;
        RECT -97.140 -178.400 -93.920 -177.920 ;
        RECT -87.220 -178.400 -84.000 -177.920 ;
        RECT -77.300 -178.400 -74.080 -177.920 ;
        RECT -67.380 -178.400 -64.160 -177.920 ;
        RECT -57.460 -178.400 -54.240 -177.920 ;
        RECT -47.540 -178.400 -44.320 -177.920 ;
        RECT -37.620 -178.400 -34.400 -177.920 ;
        RECT -27.700 -178.400 -24.480 -177.920 ;
        RECT -17.780 -178.400 -14.560 -177.920 ;
        RECT -7.860 -178.400 -4.640 -177.920 ;
        RECT 2.060 -178.400 5.280 -177.920 ;
        RECT 11.980 -178.400 15.200 -177.920 ;
        RECT 21.900 -178.400 25.120 -177.920 ;
        RECT -281.060 -179.970 -277.040 -178.590 ;
        RECT -271.140 -179.970 -267.120 -178.590 ;
        RECT -261.220 -179.970 -257.200 -178.590 ;
        RECT -251.300 -179.970 -247.280 -178.590 ;
        RECT -241.380 -179.970 -237.360 -178.590 ;
        RECT -231.460 -179.970 -227.440 -178.590 ;
        RECT -221.540 -179.970 -217.520 -178.590 ;
        RECT -211.620 -179.970 -207.600 -178.590 ;
        RECT -201.700 -179.970 -197.680 -178.590 ;
        RECT -191.780 -179.970 -187.760 -178.590 ;
        RECT -181.860 -179.970 -177.840 -178.590 ;
        RECT -171.940 -179.970 -167.920 -178.590 ;
        RECT -162.020 -179.970 -158.000 -178.590 ;
        RECT -152.100 -179.970 -148.080 -178.590 ;
        RECT -142.180 -179.970 -138.160 -178.590 ;
        RECT -132.260 -179.970 -128.240 -178.590 ;
        RECT -122.340 -179.970 -118.320 -178.590 ;
        RECT -112.420 -179.970 -108.400 -178.590 ;
        RECT -102.500 -179.970 -98.480 -178.590 ;
        RECT -92.580 -179.970 -88.560 -178.590 ;
        RECT -82.660 -179.970 -78.640 -178.590 ;
        RECT -72.740 -179.970 -68.720 -178.590 ;
        RECT -62.820 -179.970 -58.800 -178.590 ;
        RECT -52.900 -179.970 -48.880 -178.590 ;
        RECT -42.980 -179.970 -38.960 -178.590 ;
        RECT -33.060 -179.970 -29.040 -178.590 ;
        RECT -23.140 -179.970 -19.120 -178.590 ;
        RECT -13.220 -179.970 -9.200 -178.590 ;
        RECT -3.300 -179.970 0.720 -178.590 ;
        RECT 6.620 -179.970 10.640 -178.590 ;
        RECT 16.540 -179.970 20.560 -178.590 ;
      LAYER via ;
        RECT -287.695 94.070 -287.435 94.330 ;
        RECT -277.775 94.070 -277.515 94.330 ;
        RECT -267.855 94.070 -267.595 94.330 ;
        RECT -257.935 94.070 -257.675 94.330 ;
        RECT -248.015 94.070 -247.755 94.330 ;
        RECT -238.095 94.070 -237.835 94.330 ;
        RECT -228.175 94.070 -227.915 94.330 ;
        RECT -218.255 94.070 -217.995 94.330 ;
        RECT -208.335 94.070 -208.075 94.330 ;
        RECT -198.415 94.070 -198.155 94.330 ;
        RECT -188.495 94.070 -188.235 94.330 ;
        RECT -178.575 94.070 -178.315 94.330 ;
        RECT -168.655 94.070 -168.395 94.330 ;
        RECT -158.735 94.070 -158.475 94.330 ;
        RECT -148.815 94.070 -148.555 94.330 ;
        RECT -138.895 94.070 -138.635 94.330 ;
        RECT -128.975 94.070 -128.715 94.330 ;
        RECT -119.055 94.070 -118.795 94.330 ;
        RECT -109.135 94.070 -108.875 94.330 ;
        RECT -99.215 94.070 -98.955 94.330 ;
        RECT -89.295 94.070 -89.035 94.330 ;
        RECT -79.375 94.070 -79.115 94.330 ;
        RECT -69.455 94.070 -69.195 94.330 ;
        RECT -59.535 94.070 -59.275 94.330 ;
        RECT -49.615 94.070 -49.355 94.330 ;
        RECT -39.695 94.070 -39.435 94.330 ;
        RECT -29.775 94.070 -29.515 94.330 ;
        RECT -19.855 94.070 -19.595 94.330 ;
        RECT -9.935 94.070 -9.675 94.330 ;
        RECT -0.015 94.070 0.245 94.330 ;
        RECT 9.905 94.070 10.165 94.330 ;
        RECT 19.825 94.070 20.085 94.330 ;
        RECT -280.525 93.200 -280.265 93.460 ;
        RECT -280.055 93.200 -279.795 93.460 ;
        RECT -270.605 93.200 -270.345 93.460 ;
        RECT -270.135 93.200 -269.875 93.460 ;
        RECT -260.685 93.200 -260.425 93.460 ;
        RECT -260.215 93.200 -259.955 93.460 ;
        RECT -250.765 93.200 -250.505 93.460 ;
        RECT -250.295 93.200 -250.035 93.460 ;
        RECT -240.845 93.200 -240.585 93.460 ;
        RECT -240.375 93.200 -240.115 93.460 ;
        RECT -230.925 93.200 -230.665 93.460 ;
        RECT -230.455 93.200 -230.195 93.460 ;
        RECT -221.005 93.200 -220.745 93.460 ;
        RECT -220.535 93.200 -220.275 93.460 ;
        RECT -211.085 93.200 -210.825 93.460 ;
        RECT -210.615 93.200 -210.355 93.460 ;
        RECT -201.165 93.200 -200.905 93.460 ;
        RECT -200.695 93.200 -200.435 93.460 ;
        RECT -191.245 93.200 -190.985 93.460 ;
        RECT -190.775 93.200 -190.515 93.460 ;
        RECT -181.325 93.200 -181.065 93.460 ;
        RECT -180.855 93.200 -180.595 93.460 ;
        RECT -171.405 93.200 -171.145 93.460 ;
        RECT -170.935 93.200 -170.675 93.460 ;
        RECT -161.485 93.200 -161.225 93.460 ;
        RECT -161.015 93.200 -160.755 93.460 ;
        RECT -151.565 93.200 -151.305 93.460 ;
        RECT -151.095 93.200 -150.835 93.460 ;
        RECT -141.645 93.200 -141.385 93.460 ;
        RECT -141.175 93.200 -140.915 93.460 ;
        RECT -131.725 93.200 -131.465 93.460 ;
        RECT -131.255 93.200 -130.995 93.460 ;
        RECT -121.805 93.200 -121.545 93.460 ;
        RECT -121.335 93.200 -121.075 93.460 ;
        RECT -111.885 93.200 -111.625 93.460 ;
        RECT -111.415 93.200 -111.155 93.460 ;
        RECT -101.965 93.200 -101.705 93.460 ;
        RECT -101.495 93.200 -101.235 93.460 ;
        RECT -92.045 93.200 -91.785 93.460 ;
        RECT -91.575 93.200 -91.315 93.460 ;
        RECT -82.125 93.200 -81.865 93.460 ;
        RECT -81.655 93.200 -81.395 93.460 ;
        RECT -72.205 93.200 -71.945 93.460 ;
        RECT -71.735 93.200 -71.475 93.460 ;
        RECT -62.285 93.200 -62.025 93.460 ;
        RECT -61.815 93.200 -61.555 93.460 ;
        RECT -52.365 93.200 -52.105 93.460 ;
        RECT -51.895 93.200 -51.635 93.460 ;
        RECT -42.445 93.200 -42.185 93.460 ;
        RECT -41.975 93.200 -41.715 93.460 ;
        RECT -32.525 93.200 -32.265 93.460 ;
        RECT -32.055 93.200 -31.795 93.460 ;
        RECT -22.605 93.200 -22.345 93.460 ;
        RECT -22.135 93.200 -21.875 93.460 ;
        RECT -12.685 93.200 -12.425 93.460 ;
        RECT -12.215 93.200 -11.955 93.460 ;
        RECT -2.765 93.200 -2.505 93.460 ;
        RECT -2.295 93.200 -2.035 93.460 ;
        RECT 7.155 93.200 7.415 93.460 ;
        RECT 7.625 93.200 7.885 93.460 ;
        RECT 17.075 93.200 17.335 93.460 ;
        RECT 17.545 93.200 17.805 93.460 ;
        RECT -287.785 90.470 -287.525 90.730 ;
        RECT -287.325 90.480 -287.065 90.740 ;
        RECT -277.865 90.470 -277.605 90.730 ;
        RECT -277.405 90.480 -277.145 90.740 ;
        RECT -267.945 90.470 -267.685 90.730 ;
        RECT -267.485 90.480 -267.225 90.740 ;
        RECT -258.025 90.470 -257.765 90.730 ;
        RECT -257.565 90.480 -257.305 90.740 ;
        RECT -248.105 90.470 -247.845 90.730 ;
        RECT -247.645 90.480 -247.385 90.740 ;
        RECT -238.185 90.470 -237.925 90.730 ;
        RECT -237.725 90.480 -237.465 90.740 ;
        RECT -228.265 90.470 -228.005 90.730 ;
        RECT -227.805 90.480 -227.545 90.740 ;
        RECT -218.345 90.470 -218.085 90.730 ;
        RECT -217.885 90.480 -217.625 90.740 ;
        RECT -208.425 90.470 -208.165 90.730 ;
        RECT -207.965 90.480 -207.705 90.740 ;
        RECT -198.505 90.470 -198.245 90.730 ;
        RECT -198.045 90.480 -197.785 90.740 ;
        RECT -188.585 90.470 -188.325 90.730 ;
        RECT -188.125 90.480 -187.865 90.740 ;
        RECT -178.665 90.470 -178.405 90.730 ;
        RECT -178.205 90.480 -177.945 90.740 ;
        RECT -168.745 90.470 -168.485 90.730 ;
        RECT -168.285 90.480 -168.025 90.740 ;
        RECT -158.825 90.470 -158.565 90.730 ;
        RECT -158.365 90.480 -158.105 90.740 ;
        RECT -148.905 90.470 -148.645 90.730 ;
        RECT -148.445 90.480 -148.185 90.740 ;
        RECT -138.985 90.470 -138.725 90.730 ;
        RECT -138.525 90.480 -138.265 90.740 ;
        RECT -129.065 90.470 -128.805 90.730 ;
        RECT -128.605 90.480 -128.345 90.740 ;
        RECT -119.145 90.470 -118.885 90.730 ;
        RECT -118.685 90.480 -118.425 90.740 ;
        RECT -109.225 90.470 -108.965 90.730 ;
        RECT -108.765 90.480 -108.505 90.740 ;
        RECT -99.305 90.470 -99.045 90.730 ;
        RECT -98.845 90.480 -98.585 90.740 ;
        RECT -89.385 90.470 -89.125 90.730 ;
        RECT -88.925 90.480 -88.665 90.740 ;
        RECT -79.465 90.470 -79.205 90.730 ;
        RECT -79.005 90.480 -78.745 90.740 ;
        RECT -69.545 90.470 -69.285 90.730 ;
        RECT -69.085 90.480 -68.825 90.740 ;
        RECT -59.625 90.470 -59.365 90.730 ;
        RECT -59.165 90.480 -58.905 90.740 ;
        RECT -49.705 90.470 -49.445 90.730 ;
        RECT -49.245 90.480 -48.985 90.740 ;
        RECT -39.785 90.470 -39.525 90.730 ;
        RECT -39.325 90.480 -39.065 90.740 ;
        RECT -29.865 90.470 -29.605 90.730 ;
        RECT -29.405 90.480 -29.145 90.740 ;
        RECT -19.945 90.470 -19.685 90.730 ;
        RECT -19.485 90.480 -19.225 90.740 ;
        RECT -10.025 90.470 -9.765 90.730 ;
        RECT -9.565 90.480 -9.305 90.740 ;
        RECT -0.105 90.470 0.155 90.730 ;
        RECT 0.355 90.480 0.615 90.740 ;
        RECT 9.815 90.470 10.075 90.730 ;
        RECT 10.275 90.480 10.535 90.740 ;
        RECT 19.735 90.470 19.995 90.730 ;
        RECT 20.195 90.480 20.455 90.740 ;
        RECT -280.135 89.710 -279.875 89.970 ;
        RECT -270.215 89.710 -269.955 89.970 ;
        RECT -260.295 89.710 -260.035 89.970 ;
        RECT -250.375 89.710 -250.115 89.970 ;
        RECT -240.455 89.710 -240.195 89.970 ;
        RECT -230.535 89.710 -230.275 89.970 ;
        RECT -220.615 89.710 -220.355 89.970 ;
        RECT -210.695 89.710 -210.435 89.970 ;
        RECT -200.775 89.710 -200.515 89.970 ;
        RECT -190.855 89.710 -190.595 89.970 ;
        RECT -180.935 89.710 -180.675 89.970 ;
        RECT -171.015 89.710 -170.755 89.970 ;
        RECT -161.095 89.710 -160.835 89.970 ;
        RECT -151.175 89.710 -150.915 89.970 ;
        RECT -141.255 89.710 -140.995 89.970 ;
        RECT -131.335 89.710 -131.075 89.970 ;
        RECT -121.415 89.710 -121.155 89.970 ;
        RECT -111.495 89.710 -111.235 89.970 ;
        RECT -101.575 89.710 -101.315 89.970 ;
        RECT -91.655 89.710 -91.395 89.970 ;
        RECT -81.735 89.710 -81.475 89.970 ;
        RECT -71.815 89.710 -71.555 89.970 ;
        RECT -61.895 89.710 -61.635 89.970 ;
        RECT -51.975 89.710 -51.715 89.970 ;
        RECT -42.055 89.710 -41.795 89.970 ;
        RECT -32.135 89.710 -31.875 89.970 ;
        RECT -22.215 89.710 -21.955 89.970 ;
        RECT -12.295 89.710 -12.035 89.970 ;
        RECT -2.375 89.710 -2.115 89.970 ;
        RECT 7.545 89.710 7.805 89.970 ;
        RECT 17.465 89.710 17.725 89.970 ;
        RECT -287.445 6.360 -287.185 6.620 ;
        RECT -277.525 6.360 -277.265 6.620 ;
        RECT -267.605 6.360 -267.345 6.620 ;
        RECT -257.685 6.360 -257.425 6.620 ;
        RECT -247.765 6.360 -247.505 6.620 ;
        RECT -237.845 6.360 -237.585 6.620 ;
        RECT -227.925 6.360 -227.665 6.620 ;
        RECT -218.005 6.360 -217.745 6.620 ;
        RECT -208.085 6.360 -207.825 6.620 ;
        RECT -198.165 6.360 -197.905 6.620 ;
        RECT -188.245 6.360 -187.985 6.620 ;
        RECT -178.325 6.360 -178.065 6.620 ;
        RECT -168.405 6.360 -168.145 6.620 ;
        RECT -158.485 6.360 -158.225 6.620 ;
        RECT -148.565 6.360 -148.305 6.620 ;
        RECT -138.645 6.360 -138.385 6.620 ;
        RECT -128.725 6.360 -128.465 6.620 ;
        RECT -118.805 6.360 -118.545 6.620 ;
        RECT -108.885 6.360 -108.625 6.620 ;
        RECT -98.965 6.360 -98.705 6.620 ;
        RECT -89.045 6.360 -88.785 6.620 ;
        RECT -79.125 6.360 -78.865 6.620 ;
        RECT -69.205 6.360 -68.945 6.620 ;
        RECT -59.285 6.360 -59.025 6.620 ;
        RECT -49.365 6.360 -49.105 6.620 ;
        RECT -39.445 6.360 -39.185 6.620 ;
        RECT -29.525 6.360 -29.265 6.620 ;
        RECT -19.605 6.360 -19.345 6.620 ;
        RECT -9.685 6.360 -9.425 6.620 ;
        RECT 0.235 6.360 0.495 6.620 ;
        RECT 10.155 6.360 10.415 6.620 ;
        RECT 20.075 6.360 20.335 6.620 ;
        RECT -280.275 5.490 -280.015 5.750 ;
        RECT -279.805 5.490 -279.545 5.750 ;
        RECT -270.355 5.490 -270.095 5.750 ;
        RECT -269.885 5.490 -269.625 5.750 ;
        RECT -260.435 5.490 -260.175 5.750 ;
        RECT -259.965 5.490 -259.705 5.750 ;
        RECT -250.515 5.490 -250.255 5.750 ;
        RECT -250.045 5.490 -249.785 5.750 ;
        RECT -240.595 5.490 -240.335 5.750 ;
        RECT -240.125 5.490 -239.865 5.750 ;
        RECT -230.675 5.490 -230.415 5.750 ;
        RECT -230.205 5.490 -229.945 5.750 ;
        RECT -220.755 5.490 -220.495 5.750 ;
        RECT -220.285 5.490 -220.025 5.750 ;
        RECT -210.835 5.490 -210.575 5.750 ;
        RECT -210.365 5.490 -210.105 5.750 ;
        RECT -200.915 5.490 -200.655 5.750 ;
        RECT -200.445 5.490 -200.185 5.750 ;
        RECT -190.995 5.490 -190.735 5.750 ;
        RECT -190.525 5.490 -190.265 5.750 ;
        RECT -181.075 5.490 -180.815 5.750 ;
        RECT -180.605 5.490 -180.345 5.750 ;
        RECT -171.155 5.490 -170.895 5.750 ;
        RECT -170.685 5.490 -170.425 5.750 ;
        RECT -161.235 5.490 -160.975 5.750 ;
        RECT -160.765 5.490 -160.505 5.750 ;
        RECT -151.315 5.490 -151.055 5.750 ;
        RECT -150.845 5.490 -150.585 5.750 ;
        RECT -141.395 5.490 -141.135 5.750 ;
        RECT -140.925 5.490 -140.665 5.750 ;
        RECT -131.475 5.490 -131.215 5.750 ;
        RECT -131.005 5.490 -130.745 5.750 ;
        RECT -121.555 5.490 -121.295 5.750 ;
        RECT -121.085 5.490 -120.825 5.750 ;
        RECT -111.635 5.490 -111.375 5.750 ;
        RECT -111.165 5.490 -110.905 5.750 ;
        RECT -101.715 5.490 -101.455 5.750 ;
        RECT -101.245 5.490 -100.985 5.750 ;
        RECT -91.795 5.490 -91.535 5.750 ;
        RECT -91.325 5.490 -91.065 5.750 ;
        RECT -81.875 5.490 -81.615 5.750 ;
        RECT -81.405 5.490 -81.145 5.750 ;
        RECT -71.955 5.490 -71.695 5.750 ;
        RECT -71.485 5.490 -71.225 5.750 ;
        RECT -62.035 5.490 -61.775 5.750 ;
        RECT -61.565 5.490 -61.305 5.750 ;
        RECT -52.115 5.490 -51.855 5.750 ;
        RECT -51.645 5.490 -51.385 5.750 ;
        RECT -42.195 5.490 -41.935 5.750 ;
        RECT -41.725 5.490 -41.465 5.750 ;
        RECT -32.275 5.490 -32.015 5.750 ;
        RECT -31.805 5.490 -31.545 5.750 ;
        RECT -22.355 5.490 -22.095 5.750 ;
        RECT -21.885 5.490 -21.625 5.750 ;
        RECT -12.435 5.490 -12.175 5.750 ;
        RECT -11.965 5.490 -11.705 5.750 ;
        RECT -2.515 5.490 -2.255 5.750 ;
        RECT -2.045 5.490 -1.785 5.750 ;
        RECT 7.405 5.490 7.665 5.750 ;
        RECT 7.875 5.490 8.135 5.750 ;
        RECT 17.325 5.490 17.585 5.750 ;
        RECT 17.795 5.490 18.055 5.750 ;
        RECT -287.535 2.760 -287.275 3.020 ;
        RECT -287.075 2.770 -286.815 3.030 ;
        RECT -277.615 2.760 -277.355 3.020 ;
        RECT -277.155 2.770 -276.895 3.030 ;
        RECT -267.695 2.760 -267.435 3.020 ;
        RECT -267.235 2.770 -266.975 3.030 ;
        RECT -257.775 2.760 -257.515 3.020 ;
        RECT -257.315 2.770 -257.055 3.030 ;
        RECT -247.855 2.760 -247.595 3.020 ;
        RECT -247.395 2.770 -247.135 3.030 ;
        RECT -237.935 2.760 -237.675 3.020 ;
        RECT -237.475 2.770 -237.215 3.030 ;
        RECT -228.015 2.760 -227.755 3.020 ;
        RECT -227.555 2.770 -227.295 3.030 ;
        RECT -218.095 2.760 -217.835 3.020 ;
        RECT -217.635 2.770 -217.375 3.030 ;
        RECT -208.175 2.760 -207.915 3.020 ;
        RECT -207.715 2.770 -207.455 3.030 ;
        RECT -198.255 2.760 -197.995 3.020 ;
        RECT -197.795 2.770 -197.535 3.030 ;
        RECT -188.335 2.760 -188.075 3.020 ;
        RECT -187.875 2.770 -187.615 3.030 ;
        RECT -178.415 2.760 -178.155 3.020 ;
        RECT -177.955 2.770 -177.695 3.030 ;
        RECT -168.495 2.760 -168.235 3.020 ;
        RECT -168.035 2.770 -167.775 3.030 ;
        RECT -158.575 2.760 -158.315 3.020 ;
        RECT -158.115 2.770 -157.855 3.030 ;
        RECT -148.655 2.760 -148.395 3.020 ;
        RECT -148.195 2.770 -147.935 3.030 ;
        RECT -138.735 2.760 -138.475 3.020 ;
        RECT -138.275 2.770 -138.015 3.030 ;
        RECT -128.815 2.760 -128.555 3.020 ;
        RECT -128.355 2.770 -128.095 3.030 ;
        RECT -118.895 2.760 -118.635 3.020 ;
        RECT -118.435 2.770 -118.175 3.030 ;
        RECT -108.975 2.760 -108.715 3.020 ;
        RECT -108.515 2.770 -108.255 3.030 ;
        RECT -99.055 2.760 -98.795 3.020 ;
        RECT -98.595 2.770 -98.335 3.030 ;
        RECT -89.135 2.760 -88.875 3.020 ;
        RECT -88.675 2.770 -88.415 3.030 ;
        RECT -79.215 2.760 -78.955 3.020 ;
        RECT -78.755 2.770 -78.495 3.030 ;
        RECT -69.295 2.760 -69.035 3.020 ;
        RECT -68.835 2.770 -68.575 3.030 ;
        RECT -59.375 2.760 -59.115 3.020 ;
        RECT -58.915 2.770 -58.655 3.030 ;
        RECT -49.455 2.760 -49.195 3.020 ;
        RECT -48.995 2.770 -48.735 3.030 ;
        RECT -39.535 2.760 -39.275 3.020 ;
        RECT -39.075 2.770 -38.815 3.030 ;
        RECT -29.615 2.760 -29.355 3.020 ;
        RECT -29.155 2.770 -28.895 3.030 ;
        RECT -19.695 2.760 -19.435 3.020 ;
        RECT -19.235 2.770 -18.975 3.030 ;
        RECT -9.775 2.760 -9.515 3.020 ;
        RECT -9.315 2.770 -9.055 3.030 ;
        RECT 0.145 2.760 0.405 3.020 ;
        RECT 0.605 2.770 0.865 3.030 ;
        RECT 10.065 2.760 10.325 3.020 ;
        RECT 10.525 2.770 10.785 3.030 ;
        RECT 19.985 2.760 20.245 3.020 ;
        RECT 20.445 2.770 20.705 3.030 ;
        RECT -279.885 2.000 -279.625 2.260 ;
        RECT -269.965 2.000 -269.705 2.260 ;
        RECT -260.045 2.000 -259.785 2.260 ;
        RECT -250.125 2.000 -249.865 2.260 ;
        RECT -240.205 2.000 -239.945 2.260 ;
        RECT -230.285 2.000 -230.025 2.260 ;
        RECT -220.365 2.000 -220.105 2.260 ;
        RECT -210.445 2.000 -210.185 2.260 ;
        RECT -200.525 2.000 -200.265 2.260 ;
        RECT -190.605 2.000 -190.345 2.260 ;
        RECT -180.685 2.000 -180.425 2.260 ;
        RECT -170.765 2.000 -170.505 2.260 ;
        RECT -160.845 2.000 -160.585 2.260 ;
        RECT -150.925 2.000 -150.665 2.260 ;
        RECT -141.005 2.000 -140.745 2.260 ;
        RECT -131.085 2.000 -130.825 2.260 ;
        RECT -121.165 2.000 -120.905 2.260 ;
        RECT -111.245 2.000 -110.985 2.260 ;
        RECT -101.325 2.000 -101.065 2.260 ;
        RECT -91.405 2.000 -91.145 2.260 ;
        RECT -81.485 2.000 -81.225 2.260 ;
        RECT -71.565 2.000 -71.305 2.260 ;
        RECT -61.645 2.000 -61.385 2.260 ;
        RECT -51.725 2.000 -51.465 2.260 ;
        RECT -41.805 2.000 -41.545 2.260 ;
        RECT -31.885 2.000 -31.625 2.260 ;
        RECT -21.965 2.000 -21.705 2.260 ;
        RECT -12.045 2.000 -11.785 2.260 ;
        RECT -2.125 2.000 -1.865 2.260 ;
        RECT 7.795 2.000 8.055 2.260 ;
        RECT 17.715 2.000 17.975 2.260 ;
        RECT -285.685 -86.990 -285.425 -86.730 ;
        RECT -275.765 -86.990 -275.505 -86.730 ;
        RECT -265.845 -86.990 -265.585 -86.730 ;
        RECT -255.925 -86.990 -255.665 -86.730 ;
        RECT -246.005 -86.990 -245.745 -86.730 ;
        RECT -236.085 -86.990 -235.825 -86.730 ;
        RECT -226.165 -86.990 -225.905 -86.730 ;
        RECT -216.245 -86.990 -215.985 -86.730 ;
        RECT -206.325 -86.990 -206.065 -86.730 ;
        RECT -196.405 -86.990 -196.145 -86.730 ;
        RECT -186.485 -86.990 -186.225 -86.730 ;
        RECT -176.565 -86.990 -176.305 -86.730 ;
        RECT -166.645 -86.990 -166.385 -86.730 ;
        RECT -156.725 -86.990 -156.465 -86.730 ;
        RECT -146.805 -86.990 -146.545 -86.730 ;
        RECT -136.885 -86.990 -136.625 -86.730 ;
        RECT -126.965 -86.990 -126.705 -86.730 ;
        RECT -117.045 -86.990 -116.785 -86.730 ;
        RECT -107.125 -86.990 -106.865 -86.730 ;
        RECT -97.205 -86.990 -96.945 -86.730 ;
        RECT -87.285 -86.990 -87.025 -86.730 ;
        RECT -77.365 -86.990 -77.105 -86.730 ;
        RECT -67.445 -86.990 -67.185 -86.730 ;
        RECT -57.525 -86.990 -57.265 -86.730 ;
        RECT -47.605 -86.990 -47.345 -86.730 ;
        RECT -37.685 -86.990 -37.425 -86.730 ;
        RECT -27.765 -86.990 -27.505 -86.730 ;
        RECT -17.845 -86.990 -17.585 -86.730 ;
        RECT -7.925 -86.990 -7.665 -86.730 ;
        RECT 1.995 -86.990 2.255 -86.730 ;
        RECT 11.915 -86.990 12.175 -86.730 ;
        RECT 21.835 -86.990 22.095 -86.730 ;
        RECT -278.515 -87.860 -278.255 -87.600 ;
        RECT -278.045 -87.860 -277.785 -87.600 ;
        RECT -268.595 -87.860 -268.335 -87.600 ;
        RECT -268.125 -87.860 -267.865 -87.600 ;
        RECT -258.675 -87.860 -258.415 -87.600 ;
        RECT -258.205 -87.860 -257.945 -87.600 ;
        RECT -248.755 -87.860 -248.495 -87.600 ;
        RECT -248.285 -87.860 -248.025 -87.600 ;
        RECT -238.835 -87.860 -238.575 -87.600 ;
        RECT -238.365 -87.860 -238.105 -87.600 ;
        RECT -228.915 -87.860 -228.655 -87.600 ;
        RECT -228.445 -87.860 -228.185 -87.600 ;
        RECT -218.995 -87.860 -218.735 -87.600 ;
        RECT -218.525 -87.860 -218.265 -87.600 ;
        RECT -209.075 -87.860 -208.815 -87.600 ;
        RECT -208.605 -87.860 -208.345 -87.600 ;
        RECT -199.155 -87.860 -198.895 -87.600 ;
        RECT -198.685 -87.860 -198.425 -87.600 ;
        RECT -189.235 -87.860 -188.975 -87.600 ;
        RECT -188.765 -87.860 -188.505 -87.600 ;
        RECT -179.315 -87.860 -179.055 -87.600 ;
        RECT -178.845 -87.860 -178.585 -87.600 ;
        RECT -169.395 -87.860 -169.135 -87.600 ;
        RECT -168.925 -87.860 -168.665 -87.600 ;
        RECT -159.475 -87.860 -159.215 -87.600 ;
        RECT -159.005 -87.860 -158.745 -87.600 ;
        RECT -149.555 -87.860 -149.295 -87.600 ;
        RECT -149.085 -87.860 -148.825 -87.600 ;
        RECT -139.635 -87.860 -139.375 -87.600 ;
        RECT -139.165 -87.860 -138.905 -87.600 ;
        RECT -129.715 -87.860 -129.455 -87.600 ;
        RECT -129.245 -87.860 -128.985 -87.600 ;
        RECT -119.795 -87.860 -119.535 -87.600 ;
        RECT -119.325 -87.860 -119.065 -87.600 ;
        RECT -109.875 -87.860 -109.615 -87.600 ;
        RECT -109.405 -87.860 -109.145 -87.600 ;
        RECT -99.955 -87.860 -99.695 -87.600 ;
        RECT -99.485 -87.860 -99.225 -87.600 ;
        RECT -90.035 -87.860 -89.775 -87.600 ;
        RECT -89.565 -87.860 -89.305 -87.600 ;
        RECT -80.115 -87.860 -79.855 -87.600 ;
        RECT -79.645 -87.860 -79.385 -87.600 ;
        RECT -70.195 -87.860 -69.935 -87.600 ;
        RECT -69.725 -87.860 -69.465 -87.600 ;
        RECT -60.275 -87.860 -60.015 -87.600 ;
        RECT -59.805 -87.860 -59.545 -87.600 ;
        RECT -50.355 -87.860 -50.095 -87.600 ;
        RECT -49.885 -87.860 -49.625 -87.600 ;
        RECT -40.435 -87.860 -40.175 -87.600 ;
        RECT -39.965 -87.860 -39.705 -87.600 ;
        RECT -30.515 -87.860 -30.255 -87.600 ;
        RECT -30.045 -87.860 -29.785 -87.600 ;
        RECT -20.595 -87.860 -20.335 -87.600 ;
        RECT -20.125 -87.860 -19.865 -87.600 ;
        RECT -10.675 -87.860 -10.415 -87.600 ;
        RECT -10.205 -87.860 -9.945 -87.600 ;
        RECT -0.755 -87.860 -0.495 -87.600 ;
        RECT -0.285 -87.860 -0.025 -87.600 ;
        RECT 9.165 -87.860 9.425 -87.600 ;
        RECT 9.635 -87.860 9.895 -87.600 ;
        RECT 19.085 -87.860 19.345 -87.600 ;
        RECT 19.555 -87.860 19.815 -87.600 ;
        RECT -285.775 -90.590 -285.515 -90.330 ;
        RECT -285.315 -90.580 -285.055 -90.320 ;
        RECT -275.855 -90.590 -275.595 -90.330 ;
        RECT -275.395 -90.580 -275.135 -90.320 ;
        RECT -265.935 -90.590 -265.675 -90.330 ;
        RECT -265.475 -90.580 -265.215 -90.320 ;
        RECT -256.015 -90.590 -255.755 -90.330 ;
        RECT -255.555 -90.580 -255.295 -90.320 ;
        RECT -246.095 -90.590 -245.835 -90.330 ;
        RECT -245.635 -90.580 -245.375 -90.320 ;
        RECT -236.175 -90.590 -235.915 -90.330 ;
        RECT -235.715 -90.580 -235.455 -90.320 ;
        RECT -226.255 -90.590 -225.995 -90.330 ;
        RECT -225.795 -90.580 -225.535 -90.320 ;
        RECT -216.335 -90.590 -216.075 -90.330 ;
        RECT -215.875 -90.580 -215.615 -90.320 ;
        RECT -206.415 -90.590 -206.155 -90.330 ;
        RECT -205.955 -90.580 -205.695 -90.320 ;
        RECT -196.495 -90.590 -196.235 -90.330 ;
        RECT -196.035 -90.580 -195.775 -90.320 ;
        RECT -186.575 -90.590 -186.315 -90.330 ;
        RECT -186.115 -90.580 -185.855 -90.320 ;
        RECT -176.655 -90.590 -176.395 -90.330 ;
        RECT -176.195 -90.580 -175.935 -90.320 ;
        RECT -166.735 -90.590 -166.475 -90.330 ;
        RECT -166.275 -90.580 -166.015 -90.320 ;
        RECT -156.815 -90.590 -156.555 -90.330 ;
        RECT -156.355 -90.580 -156.095 -90.320 ;
        RECT -146.895 -90.590 -146.635 -90.330 ;
        RECT -146.435 -90.580 -146.175 -90.320 ;
        RECT -136.975 -90.590 -136.715 -90.330 ;
        RECT -136.515 -90.580 -136.255 -90.320 ;
        RECT -127.055 -90.590 -126.795 -90.330 ;
        RECT -126.595 -90.580 -126.335 -90.320 ;
        RECT -117.135 -90.590 -116.875 -90.330 ;
        RECT -116.675 -90.580 -116.415 -90.320 ;
        RECT -107.215 -90.590 -106.955 -90.330 ;
        RECT -106.755 -90.580 -106.495 -90.320 ;
        RECT -97.295 -90.590 -97.035 -90.330 ;
        RECT -96.835 -90.580 -96.575 -90.320 ;
        RECT -87.375 -90.590 -87.115 -90.330 ;
        RECT -86.915 -90.580 -86.655 -90.320 ;
        RECT -77.455 -90.590 -77.195 -90.330 ;
        RECT -76.995 -90.580 -76.735 -90.320 ;
        RECT -67.535 -90.590 -67.275 -90.330 ;
        RECT -67.075 -90.580 -66.815 -90.320 ;
        RECT -57.615 -90.590 -57.355 -90.330 ;
        RECT -57.155 -90.580 -56.895 -90.320 ;
        RECT -47.695 -90.590 -47.435 -90.330 ;
        RECT -47.235 -90.580 -46.975 -90.320 ;
        RECT -37.775 -90.590 -37.515 -90.330 ;
        RECT -37.315 -90.580 -37.055 -90.320 ;
        RECT -27.855 -90.590 -27.595 -90.330 ;
        RECT -27.395 -90.580 -27.135 -90.320 ;
        RECT -17.935 -90.590 -17.675 -90.330 ;
        RECT -17.475 -90.580 -17.215 -90.320 ;
        RECT -8.015 -90.590 -7.755 -90.330 ;
        RECT -7.555 -90.580 -7.295 -90.320 ;
        RECT 1.905 -90.590 2.165 -90.330 ;
        RECT 2.365 -90.580 2.625 -90.320 ;
        RECT 11.825 -90.590 12.085 -90.330 ;
        RECT 12.285 -90.580 12.545 -90.320 ;
        RECT 21.745 -90.590 22.005 -90.330 ;
        RECT 22.205 -90.580 22.465 -90.320 ;
        RECT -278.125 -91.350 -277.865 -91.090 ;
        RECT -268.205 -91.350 -267.945 -91.090 ;
        RECT -258.285 -91.350 -258.025 -91.090 ;
        RECT -248.365 -91.350 -248.105 -91.090 ;
        RECT -238.445 -91.350 -238.185 -91.090 ;
        RECT -228.525 -91.350 -228.265 -91.090 ;
        RECT -218.605 -91.350 -218.345 -91.090 ;
        RECT -208.685 -91.350 -208.425 -91.090 ;
        RECT -198.765 -91.350 -198.505 -91.090 ;
        RECT -188.845 -91.350 -188.585 -91.090 ;
        RECT -178.925 -91.350 -178.665 -91.090 ;
        RECT -169.005 -91.350 -168.745 -91.090 ;
        RECT -159.085 -91.350 -158.825 -91.090 ;
        RECT -149.165 -91.350 -148.905 -91.090 ;
        RECT -139.245 -91.350 -138.985 -91.090 ;
        RECT -129.325 -91.350 -129.065 -91.090 ;
        RECT -119.405 -91.350 -119.145 -91.090 ;
        RECT -109.485 -91.350 -109.225 -91.090 ;
        RECT -99.565 -91.350 -99.305 -91.090 ;
        RECT -89.645 -91.350 -89.385 -91.090 ;
        RECT -79.725 -91.350 -79.465 -91.090 ;
        RECT -69.805 -91.350 -69.545 -91.090 ;
        RECT -59.885 -91.350 -59.625 -91.090 ;
        RECT -49.965 -91.350 -49.705 -91.090 ;
        RECT -40.045 -91.350 -39.785 -91.090 ;
        RECT -30.125 -91.350 -29.865 -91.090 ;
        RECT -20.205 -91.350 -19.945 -91.090 ;
        RECT -10.285 -91.350 -10.025 -91.090 ;
        RECT -0.365 -91.350 -0.105 -91.090 ;
        RECT 9.555 -91.350 9.815 -91.090 ;
        RECT 19.475 -91.350 19.735 -91.090 ;
        RECT -285.435 -174.700 -285.175 -174.440 ;
        RECT -275.515 -174.700 -275.255 -174.440 ;
        RECT -265.595 -174.700 -265.335 -174.440 ;
        RECT -255.675 -174.700 -255.415 -174.440 ;
        RECT -245.755 -174.700 -245.495 -174.440 ;
        RECT -235.835 -174.700 -235.575 -174.440 ;
        RECT -225.915 -174.700 -225.655 -174.440 ;
        RECT -215.995 -174.700 -215.735 -174.440 ;
        RECT -206.075 -174.700 -205.815 -174.440 ;
        RECT -196.155 -174.700 -195.895 -174.440 ;
        RECT -186.235 -174.700 -185.975 -174.440 ;
        RECT -176.315 -174.700 -176.055 -174.440 ;
        RECT -166.395 -174.700 -166.135 -174.440 ;
        RECT -156.475 -174.700 -156.215 -174.440 ;
        RECT -146.555 -174.700 -146.295 -174.440 ;
        RECT -136.635 -174.700 -136.375 -174.440 ;
        RECT -126.715 -174.700 -126.455 -174.440 ;
        RECT -116.795 -174.700 -116.535 -174.440 ;
        RECT -106.875 -174.700 -106.615 -174.440 ;
        RECT -96.955 -174.700 -96.695 -174.440 ;
        RECT -87.035 -174.700 -86.775 -174.440 ;
        RECT -77.115 -174.700 -76.855 -174.440 ;
        RECT -67.195 -174.700 -66.935 -174.440 ;
        RECT -57.275 -174.700 -57.015 -174.440 ;
        RECT -47.355 -174.700 -47.095 -174.440 ;
        RECT -37.435 -174.700 -37.175 -174.440 ;
        RECT -27.515 -174.700 -27.255 -174.440 ;
        RECT -17.595 -174.700 -17.335 -174.440 ;
        RECT -7.675 -174.700 -7.415 -174.440 ;
        RECT 2.245 -174.700 2.505 -174.440 ;
        RECT 12.165 -174.700 12.425 -174.440 ;
        RECT 22.085 -174.700 22.345 -174.440 ;
        RECT -278.265 -175.570 -278.005 -175.310 ;
        RECT -277.795 -175.570 -277.535 -175.310 ;
        RECT -268.345 -175.570 -268.085 -175.310 ;
        RECT -267.875 -175.570 -267.615 -175.310 ;
        RECT -258.425 -175.570 -258.165 -175.310 ;
        RECT -257.955 -175.570 -257.695 -175.310 ;
        RECT -248.505 -175.570 -248.245 -175.310 ;
        RECT -248.035 -175.570 -247.775 -175.310 ;
        RECT -238.585 -175.570 -238.325 -175.310 ;
        RECT -238.115 -175.570 -237.855 -175.310 ;
        RECT -228.665 -175.570 -228.405 -175.310 ;
        RECT -228.195 -175.570 -227.935 -175.310 ;
        RECT -218.745 -175.570 -218.485 -175.310 ;
        RECT -218.275 -175.570 -218.015 -175.310 ;
        RECT -208.825 -175.570 -208.565 -175.310 ;
        RECT -208.355 -175.570 -208.095 -175.310 ;
        RECT -198.905 -175.570 -198.645 -175.310 ;
        RECT -198.435 -175.570 -198.175 -175.310 ;
        RECT -188.985 -175.570 -188.725 -175.310 ;
        RECT -188.515 -175.570 -188.255 -175.310 ;
        RECT -179.065 -175.570 -178.805 -175.310 ;
        RECT -178.595 -175.570 -178.335 -175.310 ;
        RECT -169.145 -175.570 -168.885 -175.310 ;
        RECT -168.675 -175.570 -168.415 -175.310 ;
        RECT -159.225 -175.570 -158.965 -175.310 ;
        RECT -158.755 -175.570 -158.495 -175.310 ;
        RECT -149.305 -175.570 -149.045 -175.310 ;
        RECT -148.835 -175.570 -148.575 -175.310 ;
        RECT -139.385 -175.570 -139.125 -175.310 ;
        RECT -138.915 -175.570 -138.655 -175.310 ;
        RECT -129.465 -175.570 -129.205 -175.310 ;
        RECT -128.995 -175.570 -128.735 -175.310 ;
        RECT -119.545 -175.570 -119.285 -175.310 ;
        RECT -119.075 -175.570 -118.815 -175.310 ;
        RECT -109.625 -175.570 -109.365 -175.310 ;
        RECT -109.155 -175.570 -108.895 -175.310 ;
        RECT -99.705 -175.570 -99.445 -175.310 ;
        RECT -99.235 -175.570 -98.975 -175.310 ;
        RECT -89.785 -175.570 -89.525 -175.310 ;
        RECT -89.315 -175.570 -89.055 -175.310 ;
        RECT -79.865 -175.570 -79.605 -175.310 ;
        RECT -79.395 -175.570 -79.135 -175.310 ;
        RECT -69.945 -175.570 -69.685 -175.310 ;
        RECT -69.475 -175.570 -69.215 -175.310 ;
        RECT -60.025 -175.570 -59.765 -175.310 ;
        RECT -59.555 -175.570 -59.295 -175.310 ;
        RECT -50.105 -175.570 -49.845 -175.310 ;
        RECT -49.635 -175.570 -49.375 -175.310 ;
        RECT -40.185 -175.570 -39.925 -175.310 ;
        RECT -39.715 -175.570 -39.455 -175.310 ;
        RECT -30.265 -175.570 -30.005 -175.310 ;
        RECT -29.795 -175.570 -29.535 -175.310 ;
        RECT -20.345 -175.570 -20.085 -175.310 ;
        RECT -19.875 -175.570 -19.615 -175.310 ;
        RECT -10.425 -175.570 -10.165 -175.310 ;
        RECT -9.955 -175.570 -9.695 -175.310 ;
        RECT -0.505 -175.570 -0.245 -175.310 ;
        RECT -0.035 -175.570 0.225 -175.310 ;
        RECT 9.415 -175.570 9.675 -175.310 ;
        RECT 9.885 -175.570 10.145 -175.310 ;
        RECT 19.335 -175.570 19.595 -175.310 ;
        RECT 19.805 -175.570 20.065 -175.310 ;
        RECT -285.525 -178.300 -285.265 -178.040 ;
        RECT -285.065 -178.290 -284.805 -178.030 ;
        RECT -275.605 -178.300 -275.345 -178.040 ;
        RECT -275.145 -178.290 -274.885 -178.030 ;
        RECT -265.685 -178.300 -265.425 -178.040 ;
        RECT -265.225 -178.290 -264.965 -178.030 ;
        RECT -255.765 -178.300 -255.505 -178.040 ;
        RECT -255.305 -178.290 -255.045 -178.030 ;
        RECT -245.845 -178.300 -245.585 -178.040 ;
        RECT -245.385 -178.290 -245.125 -178.030 ;
        RECT -235.925 -178.300 -235.665 -178.040 ;
        RECT -235.465 -178.290 -235.205 -178.030 ;
        RECT -226.005 -178.300 -225.745 -178.040 ;
        RECT -225.545 -178.290 -225.285 -178.030 ;
        RECT -216.085 -178.300 -215.825 -178.040 ;
        RECT -215.625 -178.290 -215.365 -178.030 ;
        RECT -206.165 -178.300 -205.905 -178.040 ;
        RECT -205.705 -178.290 -205.445 -178.030 ;
        RECT -196.245 -178.300 -195.985 -178.040 ;
        RECT -195.785 -178.290 -195.525 -178.030 ;
        RECT -186.325 -178.300 -186.065 -178.040 ;
        RECT -185.865 -178.290 -185.605 -178.030 ;
        RECT -176.405 -178.300 -176.145 -178.040 ;
        RECT -175.945 -178.290 -175.685 -178.030 ;
        RECT -166.485 -178.300 -166.225 -178.040 ;
        RECT -166.025 -178.290 -165.765 -178.030 ;
        RECT -156.565 -178.300 -156.305 -178.040 ;
        RECT -156.105 -178.290 -155.845 -178.030 ;
        RECT -146.645 -178.300 -146.385 -178.040 ;
        RECT -146.185 -178.290 -145.925 -178.030 ;
        RECT -136.725 -178.300 -136.465 -178.040 ;
        RECT -136.265 -178.290 -136.005 -178.030 ;
        RECT -126.805 -178.300 -126.545 -178.040 ;
        RECT -126.345 -178.290 -126.085 -178.030 ;
        RECT -116.885 -178.300 -116.625 -178.040 ;
        RECT -116.425 -178.290 -116.165 -178.030 ;
        RECT -106.965 -178.300 -106.705 -178.040 ;
        RECT -106.505 -178.290 -106.245 -178.030 ;
        RECT -97.045 -178.300 -96.785 -178.040 ;
        RECT -96.585 -178.290 -96.325 -178.030 ;
        RECT -87.125 -178.300 -86.865 -178.040 ;
        RECT -86.665 -178.290 -86.405 -178.030 ;
        RECT -77.205 -178.300 -76.945 -178.040 ;
        RECT -76.745 -178.290 -76.485 -178.030 ;
        RECT -67.285 -178.300 -67.025 -178.040 ;
        RECT -66.825 -178.290 -66.565 -178.030 ;
        RECT -57.365 -178.300 -57.105 -178.040 ;
        RECT -56.905 -178.290 -56.645 -178.030 ;
        RECT -47.445 -178.300 -47.185 -178.040 ;
        RECT -46.985 -178.290 -46.725 -178.030 ;
        RECT -37.525 -178.300 -37.265 -178.040 ;
        RECT -37.065 -178.290 -36.805 -178.030 ;
        RECT -27.605 -178.300 -27.345 -178.040 ;
        RECT -27.145 -178.290 -26.885 -178.030 ;
        RECT -17.685 -178.300 -17.425 -178.040 ;
        RECT -17.225 -178.290 -16.965 -178.030 ;
        RECT -7.765 -178.300 -7.505 -178.040 ;
        RECT -7.305 -178.290 -7.045 -178.030 ;
        RECT 2.155 -178.300 2.415 -178.040 ;
        RECT 2.615 -178.290 2.875 -178.030 ;
        RECT 12.075 -178.300 12.335 -178.040 ;
        RECT 12.535 -178.290 12.795 -178.030 ;
        RECT 21.995 -178.300 22.255 -178.040 ;
        RECT 22.455 -178.290 22.715 -178.030 ;
        RECT -277.875 -179.060 -277.615 -178.800 ;
        RECT -267.955 -179.060 -267.695 -178.800 ;
        RECT -258.035 -179.060 -257.775 -178.800 ;
        RECT -248.115 -179.060 -247.855 -178.800 ;
        RECT -238.195 -179.060 -237.935 -178.800 ;
        RECT -228.275 -179.060 -228.015 -178.800 ;
        RECT -218.355 -179.060 -218.095 -178.800 ;
        RECT -208.435 -179.060 -208.175 -178.800 ;
        RECT -198.515 -179.060 -198.255 -178.800 ;
        RECT -188.595 -179.060 -188.335 -178.800 ;
        RECT -178.675 -179.060 -178.415 -178.800 ;
        RECT -168.755 -179.060 -168.495 -178.800 ;
        RECT -158.835 -179.060 -158.575 -178.800 ;
        RECT -148.915 -179.060 -148.655 -178.800 ;
        RECT -138.995 -179.060 -138.735 -178.800 ;
        RECT -129.075 -179.060 -128.815 -178.800 ;
        RECT -119.155 -179.060 -118.895 -178.800 ;
        RECT -109.235 -179.060 -108.975 -178.800 ;
        RECT -99.315 -179.060 -99.055 -178.800 ;
        RECT -89.395 -179.060 -89.135 -178.800 ;
        RECT -79.475 -179.060 -79.215 -178.800 ;
        RECT -69.555 -179.060 -69.295 -178.800 ;
        RECT -59.635 -179.060 -59.375 -178.800 ;
        RECT -49.715 -179.060 -49.455 -178.800 ;
        RECT -39.795 -179.060 -39.535 -178.800 ;
        RECT -29.875 -179.060 -29.615 -178.800 ;
        RECT -19.955 -179.060 -19.695 -178.800 ;
        RECT -10.035 -179.060 -9.775 -178.800 ;
        RECT -0.115 -179.060 0.145 -178.800 ;
        RECT 9.805 -179.060 10.065 -178.800 ;
        RECT 19.725 -179.060 19.985 -178.800 ;
      LAYER met2 ;
        RECT -288.280 93.760 -287.110 94.560 ;
        RECT -278.360 93.760 -277.190 94.560 ;
        RECT -268.440 93.760 -267.270 94.560 ;
        RECT -258.520 93.760 -257.350 94.560 ;
        RECT -248.600 93.760 -247.430 94.560 ;
        RECT -238.680 93.760 -237.510 94.560 ;
        RECT -228.760 93.760 -227.590 94.560 ;
        RECT -218.840 93.760 -217.670 94.560 ;
        RECT -208.920 93.760 -207.750 94.560 ;
        RECT -199.000 93.760 -197.830 94.560 ;
        RECT -189.080 93.760 -187.910 94.560 ;
        RECT -179.160 93.760 -177.990 94.560 ;
        RECT -169.240 93.760 -168.070 94.560 ;
        RECT -159.320 93.760 -158.150 94.560 ;
        RECT -149.400 93.760 -148.230 94.560 ;
        RECT -139.480 93.760 -138.310 94.560 ;
        RECT -129.560 93.760 -128.390 94.560 ;
        RECT -119.640 93.760 -118.470 94.560 ;
        RECT -109.720 93.760 -108.550 94.560 ;
        RECT -99.800 93.760 -98.630 94.560 ;
        RECT -89.880 93.760 -88.710 94.560 ;
        RECT -79.960 93.760 -78.790 94.560 ;
        RECT -70.040 93.760 -68.870 94.560 ;
        RECT -60.120 93.760 -58.950 94.560 ;
        RECT -50.200 93.760 -49.030 94.560 ;
        RECT -40.280 93.760 -39.110 94.560 ;
        RECT -30.360 93.760 -29.190 94.560 ;
        RECT -20.440 93.760 -19.270 94.560 ;
        RECT -10.520 93.760 -9.350 94.560 ;
        RECT -0.600 93.760 0.570 94.560 ;
        RECT 9.320 93.760 10.490 94.560 ;
        RECT 19.240 93.760 20.410 94.560 ;
        RECT -280.620 93.090 -279.700 93.570 ;
        RECT -270.700 93.090 -269.780 93.570 ;
        RECT -260.780 93.090 -259.860 93.570 ;
        RECT -250.860 93.090 -249.940 93.570 ;
        RECT -240.940 93.090 -240.020 93.570 ;
        RECT -231.020 93.090 -230.100 93.570 ;
        RECT -221.100 93.090 -220.180 93.570 ;
        RECT -211.180 93.090 -210.260 93.570 ;
        RECT -201.260 93.090 -200.340 93.570 ;
        RECT -191.340 93.090 -190.420 93.570 ;
        RECT -181.420 93.090 -180.500 93.570 ;
        RECT -171.500 93.090 -170.580 93.570 ;
        RECT -161.580 93.090 -160.660 93.570 ;
        RECT -151.660 93.090 -150.740 93.570 ;
        RECT -141.740 93.090 -140.820 93.570 ;
        RECT -131.820 93.090 -130.900 93.570 ;
        RECT -121.900 93.090 -120.980 93.570 ;
        RECT -111.980 93.090 -111.060 93.570 ;
        RECT -102.060 93.090 -101.140 93.570 ;
        RECT -92.140 93.090 -91.220 93.570 ;
        RECT -82.220 93.090 -81.300 93.570 ;
        RECT -72.300 93.090 -71.380 93.570 ;
        RECT -62.380 93.090 -61.460 93.570 ;
        RECT -52.460 93.090 -51.540 93.570 ;
        RECT -42.540 93.090 -41.620 93.570 ;
        RECT -32.620 93.090 -31.700 93.570 ;
        RECT -22.700 93.090 -21.780 93.570 ;
        RECT -12.780 93.090 -11.860 93.570 ;
        RECT -2.860 93.090 -1.940 93.570 ;
        RECT 7.060 93.090 7.980 93.570 ;
        RECT 16.980 93.090 17.900 93.570 ;
        RECT -287.880 90.370 -286.960 90.850 ;
        RECT -277.960 90.370 -277.040 90.850 ;
        RECT -268.040 90.370 -267.120 90.850 ;
        RECT -258.120 90.370 -257.200 90.850 ;
        RECT -248.200 90.370 -247.280 90.850 ;
        RECT -238.280 90.370 -237.360 90.850 ;
        RECT -228.360 90.370 -227.440 90.850 ;
        RECT -218.440 90.370 -217.520 90.850 ;
        RECT -208.520 90.370 -207.600 90.850 ;
        RECT -198.600 90.370 -197.680 90.850 ;
        RECT -188.680 90.370 -187.760 90.850 ;
        RECT -178.760 90.370 -177.840 90.850 ;
        RECT -168.840 90.370 -167.920 90.850 ;
        RECT -158.920 90.370 -158.000 90.850 ;
        RECT -149.000 90.370 -148.080 90.850 ;
        RECT -139.080 90.370 -138.160 90.850 ;
        RECT -129.160 90.370 -128.240 90.850 ;
        RECT -119.240 90.370 -118.320 90.850 ;
        RECT -109.320 90.370 -108.400 90.850 ;
        RECT -99.400 90.370 -98.480 90.850 ;
        RECT -89.480 90.370 -88.560 90.850 ;
        RECT -79.560 90.370 -78.640 90.850 ;
        RECT -69.640 90.370 -68.720 90.850 ;
        RECT -59.720 90.370 -58.800 90.850 ;
        RECT -49.800 90.370 -48.880 90.850 ;
        RECT -39.880 90.370 -38.960 90.850 ;
        RECT -29.960 90.370 -29.040 90.850 ;
        RECT -20.040 90.370 -19.120 90.850 ;
        RECT -10.120 90.370 -9.200 90.850 ;
        RECT -0.200 90.370 0.720 90.850 ;
        RECT 9.720 90.370 10.640 90.850 ;
        RECT 19.640 90.370 20.560 90.850 ;
        RECT -280.460 89.390 -279.290 90.190 ;
        RECT -270.540 89.390 -269.370 90.190 ;
        RECT -260.620 89.390 -259.450 90.190 ;
        RECT -250.700 89.390 -249.530 90.190 ;
        RECT -240.780 89.390 -239.610 90.190 ;
        RECT -230.860 89.390 -229.690 90.190 ;
        RECT -220.940 89.390 -219.770 90.190 ;
        RECT -211.020 89.390 -209.850 90.190 ;
        RECT -201.100 89.390 -199.930 90.190 ;
        RECT -191.180 89.390 -190.010 90.190 ;
        RECT -181.260 89.390 -180.090 90.190 ;
        RECT -171.340 89.390 -170.170 90.190 ;
        RECT -161.420 89.390 -160.250 90.190 ;
        RECT -151.500 89.390 -150.330 90.190 ;
        RECT -141.580 89.390 -140.410 90.190 ;
        RECT -131.660 89.390 -130.490 90.190 ;
        RECT -121.740 89.390 -120.570 90.190 ;
        RECT -111.820 89.390 -110.650 90.190 ;
        RECT -101.900 89.390 -100.730 90.190 ;
        RECT -91.980 89.390 -90.810 90.190 ;
        RECT -82.060 89.390 -80.890 90.190 ;
        RECT -72.140 89.390 -70.970 90.190 ;
        RECT -62.220 89.390 -61.050 90.190 ;
        RECT -52.300 89.390 -51.130 90.190 ;
        RECT -42.380 89.390 -41.210 90.190 ;
        RECT -32.460 89.390 -31.290 90.190 ;
        RECT -22.540 89.390 -21.370 90.190 ;
        RECT -12.620 89.390 -11.450 90.190 ;
        RECT -2.700 89.390 -1.530 90.190 ;
        RECT 7.220 89.390 8.390 90.190 ;
        RECT 17.140 89.390 18.310 90.190 ;
        RECT -288.030 6.050 -286.860 6.850 ;
        RECT -278.110 6.050 -276.940 6.850 ;
        RECT -268.190 6.050 -267.020 6.850 ;
        RECT -258.270 6.050 -257.100 6.850 ;
        RECT -248.350 6.050 -247.180 6.850 ;
        RECT -238.430 6.050 -237.260 6.850 ;
        RECT -228.510 6.050 -227.340 6.850 ;
        RECT -218.590 6.050 -217.420 6.850 ;
        RECT -208.670 6.050 -207.500 6.850 ;
        RECT -198.750 6.050 -197.580 6.850 ;
        RECT -188.830 6.050 -187.660 6.850 ;
        RECT -178.910 6.050 -177.740 6.850 ;
        RECT -168.990 6.050 -167.820 6.850 ;
        RECT -159.070 6.050 -157.900 6.850 ;
        RECT -149.150 6.050 -147.980 6.850 ;
        RECT -139.230 6.050 -138.060 6.850 ;
        RECT -129.310 6.050 -128.140 6.850 ;
        RECT -119.390 6.050 -118.220 6.850 ;
        RECT -109.470 6.050 -108.300 6.850 ;
        RECT -99.550 6.050 -98.380 6.850 ;
        RECT -89.630 6.050 -88.460 6.850 ;
        RECT -79.710 6.050 -78.540 6.850 ;
        RECT -69.790 6.050 -68.620 6.850 ;
        RECT -59.870 6.050 -58.700 6.850 ;
        RECT -49.950 6.050 -48.780 6.850 ;
        RECT -40.030 6.050 -38.860 6.850 ;
        RECT -30.110 6.050 -28.940 6.850 ;
        RECT -20.190 6.050 -19.020 6.850 ;
        RECT -10.270 6.050 -9.100 6.850 ;
        RECT -0.350 6.050 0.820 6.850 ;
        RECT 9.570 6.050 10.740 6.850 ;
        RECT 19.490 6.050 20.660 6.850 ;
        RECT -280.370 5.380 -279.450 5.860 ;
        RECT -270.450 5.380 -269.530 5.860 ;
        RECT -260.530 5.380 -259.610 5.860 ;
        RECT -250.610 5.380 -249.690 5.860 ;
        RECT -240.690 5.380 -239.770 5.860 ;
        RECT -230.770 5.380 -229.850 5.860 ;
        RECT -220.850 5.380 -219.930 5.860 ;
        RECT -210.930 5.380 -210.010 5.860 ;
        RECT -201.010 5.380 -200.090 5.860 ;
        RECT -191.090 5.380 -190.170 5.860 ;
        RECT -181.170 5.380 -180.250 5.860 ;
        RECT -171.250 5.380 -170.330 5.860 ;
        RECT -161.330 5.380 -160.410 5.860 ;
        RECT -151.410 5.380 -150.490 5.860 ;
        RECT -141.490 5.380 -140.570 5.860 ;
        RECT -131.570 5.380 -130.650 5.860 ;
        RECT -121.650 5.380 -120.730 5.860 ;
        RECT -111.730 5.380 -110.810 5.860 ;
        RECT -101.810 5.380 -100.890 5.860 ;
        RECT -91.890 5.380 -90.970 5.860 ;
        RECT -81.970 5.380 -81.050 5.860 ;
        RECT -72.050 5.380 -71.130 5.860 ;
        RECT -62.130 5.380 -61.210 5.860 ;
        RECT -52.210 5.380 -51.290 5.860 ;
        RECT -42.290 5.380 -41.370 5.860 ;
        RECT -32.370 5.380 -31.450 5.860 ;
        RECT -22.450 5.380 -21.530 5.860 ;
        RECT -12.530 5.380 -11.610 5.860 ;
        RECT -2.610 5.380 -1.690 5.860 ;
        RECT 7.310 5.380 8.230 5.860 ;
        RECT 17.230 5.380 18.150 5.860 ;
        RECT -287.630 2.660 -286.710 3.140 ;
        RECT -277.710 2.660 -276.790 3.140 ;
        RECT -267.790 2.660 -266.870 3.140 ;
        RECT -257.870 2.660 -256.950 3.140 ;
        RECT -247.950 2.660 -247.030 3.140 ;
        RECT -238.030 2.660 -237.110 3.140 ;
        RECT -228.110 2.660 -227.190 3.140 ;
        RECT -218.190 2.660 -217.270 3.140 ;
        RECT -208.270 2.660 -207.350 3.140 ;
        RECT -198.350 2.660 -197.430 3.140 ;
        RECT -188.430 2.660 -187.510 3.140 ;
        RECT -178.510 2.660 -177.590 3.140 ;
        RECT -168.590 2.660 -167.670 3.140 ;
        RECT -158.670 2.660 -157.750 3.140 ;
        RECT -148.750 2.660 -147.830 3.140 ;
        RECT -138.830 2.660 -137.910 3.140 ;
        RECT -128.910 2.660 -127.990 3.140 ;
        RECT -118.990 2.660 -118.070 3.140 ;
        RECT -109.070 2.660 -108.150 3.140 ;
        RECT -99.150 2.660 -98.230 3.140 ;
        RECT -89.230 2.660 -88.310 3.140 ;
        RECT -79.310 2.660 -78.390 3.140 ;
        RECT -69.390 2.660 -68.470 3.140 ;
        RECT -59.470 2.660 -58.550 3.140 ;
        RECT -49.550 2.660 -48.630 3.140 ;
        RECT -39.630 2.660 -38.710 3.140 ;
        RECT -29.710 2.660 -28.790 3.140 ;
        RECT -19.790 2.660 -18.870 3.140 ;
        RECT -9.870 2.660 -8.950 3.140 ;
        RECT 0.050 2.660 0.970 3.140 ;
        RECT 9.970 2.660 10.890 3.140 ;
        RECT 19.890 2.660 20.810 3.140 ;
        RECT -280.210 1.680 -279.040 2.480 ;
        RECT -270.290 1.680 -269.120 2.480 ;
        RECT -260.370 1.680 -259.200 2.480 ;
        RECT -250.450 1.680 -249.280 2.480 ;
        RECT -240.530 1.680 -239.360 2.480 ;
        RECT -230.610 1.680 -229.440 2.480 ;
        RECT -220.690 1.680 -219.520 2.480 ;
        RECT -210.770 1.680 -209.600 2.480 ;
        RECT -200.850 1.680 -199.680 2.480 ;
        RECT -190.930 1.680 -189.760 2.480 ;
        RECT -181.010 1.680 -179.840 2.480 ;
        RECT -171.090 1.680 -169.920 2.480 ;
        RECT -161.170 1.680 -160.000 2.480 ;
        RECT -151.250 1.680 -150.080 2.480 ;
        RECT -141.330 1.680 -140.160 2.480 ;
        RECT -131.410 1.680 -130.240 2.480 ;
        RECT -121.490 1.680 -120.320 2.480 ;
        RECT -111.570 1.680 -110.400 2.480 ;
        RECT -101.650 1.680 -100.480 2.480 ;
        RECT -91.730 1.680 -90.560 2.480 ;
        RECT -81.810 1.680 -80.640 2.480 ;
        RECT -71.890 1.680 -70.720 2.480 ;
        RECT -61.970 1.680 -60.800 2.480 ;
        RECT -52.050 1.680 -50.880 2.480 ;
        RECT -42.130 1.680 -40.960 2.480 ;
        RECT -32.210 1.680 -31.040 2.480 ;
        RECT -22.290 1.680 -21.120 2.480 ;
        RECT -12.370 1.680 -11.200 2.480 ;
        RECT -2.450 1.680 -1.280 2.480 ;
        RECT 7.470 1.680 8.640 2.480 ;
        RECT 17.390 1.680 18.560 2.480 ;
        RECT -286.270 -87.300 -285.100 -86.500 ;
        RECT -276.350 -87.300 -275.180 -86.500 ;
        RECT -266.430 -87.300 -265.260 -86.500 ;
        RECT -256.510 -87.300 -255.340 -86.500 ;
        RECT -246.590 -87.300 -245.420 -86.500 ;
        RECT -236.670 -87.300 -235.500 -86.500 ;
        RECT -226.750 -87.300 -225.580 -86.500 ;
        RECT -216.830 -87.300 -215.660 -86.500 ;
        RECT -206.910 -87.300 -205.740 -86.500 ;
        RECT -196.990 -87.300 -195.820 -86.500 ;
        RECT -187.070 -87.300 -185.900 -86.500 ;
        RECT -177.150 -87.300 -175.980 -86.500 ;
        RECT -167.230 -87.300 -166.060 -86.500 ;
        RECT -157.310 -87.300 -156.140 -86.500 ;
        RECT -147.390 -87.300 -146.220 -86.500 ;
        RECT -137.470 -87.300 -136.300 -86.500 ;
        RECT -127.550 -87.300 -126.380 -86.500 ;
        RECT -117.630 -87.300 -116.460 -86.500 ;
        RECT -107.710 -87.300 -106.540 -86.500 ;
        RECT -97.790 -87.300 -96.620 -86.500 ;
        RECT -87.870 -87.300 -86.700 -86.500 ;
        RECT -77.950 -87.300 -76.780 -86.500 ;
        RECT -68.030 -87.300 -66.860 -86.500 ;
        RECT -58.110 -87.300 -56.940 -86.500 ;
        RECT -48.190 -87.300 -47.020 -86.500 ;
        RECT -38.270 -87.300 -37.100 -86.500 ;
        RECT -28.350 -87.300 -27.180 -86.500 ;
        RECT -18.430 -87.300 -17.260 -86.500 ;
        RECT -8.510 -87.300 -7.340 -86.500 ;
        RECT 1.410 -87.300 2.580 -86.500 ;
        RECT 11.330 -87.300 12.500 -86.500 ;
        RECT 21.250 -87.300 22.420 -86.500 ;
        RECT -278.610 -87.970 -277.690 -87.490 ;
        RECT -268.690 -87.970 -267.770 -87.490 ;
        RECT -258.770 -87.970 -257.850 -87.490 ;
        RECT -248.850 -87.970 -247.930 -87.490 ;
        RECT -238.930 -87.970 -238.010 -87.490 ;
        RECT -229.010 -87.970 -228.090 -87.490 ;
        RECT -219.090 -87.970 -218.170 -87.490 ;
        RECT -209.170 -87.970 -208.250 -87.490 ;
        RECT -199.250 -87.970 -198.330 -87.490 ;
        RECT -189.330 -87.970 -188.410 -87.490 ;
        RECT -179.410 -87.970 -178.490 -87.490 ;
        RECT -169.490 -87.970 -168.570 -87.490 ;
        RECT -159.570 -87.970 -158.650 -87.490 ;
        RECT -149.650 -87.970 -148.730 -87.490 ;
        RECT -139.730 -87.970 -138.810 -87.490 ;
        RECT -129.810 -87.970 -128.890 -87.490 ;
        RECT -119.890 -87.970 -118.970 -87.490 ;
        RECT -109.970 -87.970 -109.050 -87.490 ;
        RECT -100.050 -87.970 -99.130 -87.490 ;
        RECT -90.130 -87.970 -89.210 -87.490 ;
        RECT -80.210 -87.970 -79.290 -87.490 ;
        RECT -70.290 -87.970 -69.370 -87.490 ;
        RECT -60.370 -87.970 -59.450 -87.490 ;
        RECT -50.450 -87.970 -49.530 -87.490 ;
        RECT -40.530 -87.970 -39.610 -87.490 ;
        RECT -30.610 -87.970 -29.690 -87.490 ;
        RECT -20.690 -87.970 -19.770 -87.490 ;
        RECT -10.770 -87.970 -9.850 -87.490 ;
        RECT -0.850 -87.970 0.070 -87.490 ;
        RECT 9.070 -87.970 9.990 -87.490 ;
        RECT 18.990 -87.970 19.910 -87.490 ;
        RECT -285.870 -90.690 -284.950 -90.210 ;
        RECT -275.950 -90.690 -275.030 -90.210 ;
        RECT -266.030 -90.690 -265.110 -90.210 ;
        RECT -256.110 -90.690 -255.190 -90.210 ;
        RECT -246.190 -90.690 -245.270 -90.210 ;
        RECT -236.270 -90.690 -235.350 -90.210 ;
        RECT -226.350 -90.690 -225.430 -90.210 ;
        RECT -216.430 -90.690 -215.510 -90.210 ;
        RECT -206.510 -90.690 -205.590 -90.210 ;
        RECT -196.590 -90.690 -195.670 -90.210 ;
        RECT -186.670 -90.690 -185.750 -90.210 ;
        RECT -176.750 -90.690 -175.830 -90.210 ;
        RECT -166.830 -90.690 -165.910 -90.210 ;
        RECT -156.910 -90.690 -155.990 -90.210 ;
        RECT -146.990 -90.690 -146.070 -90.210 ;
        RECT -137.070 -90.690 -136.150 -90.210 ;
        RECT -127.150 -90.690 -126.230 -90.210 ;
        RECT -117.230 -90.690 -116.310 -90.210 ;
        RECT -107.310 -90.690 -106.390 -90.210 ;
        RECT -97.390 -90.690 -96.470 -90.210 ;
        RECT -87.470 -90.690 -86.550 -90.210 ;
        RECT -77.550 -90.690 -76.630 -90.210 ;
        RECT -67.630 -90.690 -66.710 -90.210 ;
        RECT -57.710 -90.690 -56.790 -90.210 ;
        RECT -47.790 -90.690 -46.870 -90.210 ;
        RECT -37.870 -90.690 -36.950 -90.210 ;
        RECT -27.950 -90.690 -27.030 -90.210 ;
        RECT -18.030 -90.690 -17.110 -90.210 ;
        RECT -8.110 -90.690 -7.190 -90.210 ;
        RECT 1.810 -90.690 2.730 -90.210 ;
        RECT 11.730 -90.690 12.650 -90.210 ;
        RECT 21.650 -90.690 22.570 -90.210 ;
        RECT -278.450 -91.670 -277.280 -90.870 ;
        RECT -268.530 -91.670 -267.360 -90.870 ;
        RECT -258.610 -91.670 -257.440 -90.870 ;
        RECT -248.690 -91.670 -247.520 -90.870 ;
        RECT -238.770 -91.670 -237.600 -90.870 ;
        RECT -228.850 -91.670 -227.680 -90.870 ;
        RECT -218.930 -91.670 -217.760 -90.870 ;
        RECT -209.010 -91.670 -207.840 -90.870 ;
        RECT -199.090 -91.670 -197.920 -90.870 ;
        RECT -189.170 -91.670 -188.000 -90.870 ;
        RECT -179.250 -91.670 -178.080 -90.870 ;
        RECT -169.330 -91.670 -168.160 -90.870 ;
        RECT -159.410 -91.670 -158.240 -90.870 ;
        RECT -149.490 -91.670 -148.320 -90.870 ;
        RECT -139.570 -91.670 -138.400 -90.870 ;
        RECT -129.650 -91.670 -128.480 -90.870 ;
        RECT -119.730 -91.670 -118.560 -90.870 ;
        RECT -109.810 -91.670 -108.640 -90.870 ;
        RECT -99.890 -91.670 -98.720 -90.870 ;
        RECT -89.970 -91.670 -88.800 -90.870 ;
        RECT -80.050 -91.670 -78.880 -90.870 ;
        RECT -70.130 -91.670 -68.960 -90.870 ;
        RECT -60.210 -91.670 -59.040 -90.870 ;
        RECT -50.290 -91.670 -49.120 -90.870 ;
        RECT -40.370 -91.670 -39.200 -90.870 ;
        RECT -30.450 -91.670 -29.280 -90.870 ;
        RECT -20.530 -91.670 -19.360 -90.870 ;
        RECT -10.610 -91.670 -9.440 -90.870 ;
        RECT -0.690 -91.670 0.480 -90.870 ;
        RECT 9.230 -91.670 10.400 -90.870 ;
        RECT 19.150 -91.670 20.320 -90.870 ;
        RECT -286.020 -175.010 -284.850 -174.210 ;
        RECT -276.100 -175.010 -274.930 -174.210 ;
        RECT -266.180 -175.010 -265.010 -174.210 ;
        RECT -256.260 -175.010 -255.090 -174.210 ;
        RECT -246.340 -175.010 -245.170 -174.210 ;
        RECT -236.420 -175.010 -235.250 -174.210 ;
        RECT -226.500 -175.010 -225.330 -174.210 ;
        RECT -216.580 -175.010 -215.410 -174.210 ;
        RECT -206.660 -175.010 -205.490 -174.210 ;
        RECT -196.740 -175.010 -195.570 -174.210 ;
        RECT -186.820 -175.010 -185.650 -174.210 ;
        RECT -176.900 -175.010 -175.730 -174.210 ;
        RECT -166.980 -175.010 -165.810 -174.210 ;
        RECT -157.060 -175.010 -155.890 -174.210 ;
        RECT -147.140 -175.010 -145.970 -174.210 ;
        RECT -137.220 -175.010 -136.050 -174.210 ;
        RECT -127.300 -175.010 -126.130 -174.210 ;
        RECT -117.380 -175.010 -116.210 -174.210 ;
        RECT -107.460 -175.010 -106.290 -174.210 ;
        RECT -97.540 -175.010 -96.370 -174.210 ;
        RECT -87.620 -175.010 -86.450 -174.210 ;
        RECT -77.700 -175.010 -76.530 -174.210 ;
        RECT -67.780 -175.010 -66.610 -174.210 ;
        RECT -57.860 -175.010 -56.690 -174.210 ;
        RECT -47.940 -175.010 -46.770 -174.210 ;
        RECT -38.020 -175.010 -36.850 -174.210 ;
        RECT -28.100 -175.010 -26.930 -174.210 ;
        RECT -18.180 -175.010 -17.010 -174.210 ;
        RECT -8.260 -175.010 -7.090 -174.210 ;
        RECT 1.660 -175.010 2.830 -174.210 ;
        RECT 11.580 -175.010 12.750 -174.210 ;
        RECT 21.500 -175.010 22.670 -174.210 ;
        RECT -278.360 -175.680 -277.440 -175.200 ;
        RECT -268.440 -175.680 -267.520 -175.200 ;
        RECT -258.520 -175.680 -257.600 -175.200 ;
        RECT -248.600 -175.680 -247.680 -175.200 ;
        RECT -238.680 -175.680 -237.760 -175.200 ;
        RECT -228.760 -175.680 -227.840 -175.200 ;
        RECT -218.840 -175.680 -217.920 -175.200 ;
        RECT -208.920 -175.680 -208.000 -175.200 ;
        RECT -199.000 -175.680 -198.080 -175.200 ;
        RECT -189.080 -175.680 -188.160 -175.200 ;
        RECT -179.160 -175.680 -178.240 -175.200 ;
        RECT -169.240 -175.680 -168.320 -175.200 ;
        RECT -159.320 -175.680 -158.400 -175.200 ;
        RECT -149.400 -175.680 -148.480 -175.200 ;
        RECT -139.480 -175.680 -138.560 -175.200 ;
        RECT -129.560 -175.680 -128.640 -175.200 ;
        RECT -119.640 -175.680 -118.720 -175.200 ;
        RECT -109.720 -175.680 -108.800 -175.200 ;
        RECT -99.800 -175.680 -98.880 -175.200 ;
        RECT -89.880 -175.680 -88.960 -175.200 ;
        RECT -79.960 -175.680 -79.040 -175.200 ;
        RECT -70.040 -175.680 -69.120 -175.200 ;
        RECT -60.120 -175.680 -59.200 -175.200 ;
        RECT -50.200 -175.680 -49.280 -175.200 ;
        RECT -40.280 -175.680 -39.360 -175.200 ;
        RECT -30.360 -175.680 -29.440 -175.200 ;
        RECT -20.440 -175.680 -19.520 -175.200 ;
        RECT -10.520 -175.680 -9.600 -175.200 ;
        RECT -0.600 -175.680 0.320 -175.200 ;
        RECT 9.320 -175.680 10.240 -175.200 ;
        RECT 19.240 -175.680 20.160 -175.200 ;
        RECT -285.620 -178.400 -284.700 -177.920 ;
        RECT -275.700 -178.400 -274.780 -177.920 ;
        RECT -265.780 -178.400 -264.860 -177.920 ;
        RECT -255.860 -178.400 -254.940 -177.920 ;
        RECT -245.940 -178.400 -245.020 -177.920 ;
        RECT -236.020 -178.400 -235.100 -177.920 ;
        RECT -226.100 -178.400 -225.180 -177.920 ;
        RECT -216.180 -178.400 -215.260 -177.920 ;
        RECT -206.260 -178.400 -205.340 -177.920 ;
        RECT -196.340 -178.400 -195.420 -177.920 ;
        RECT -186.420 -178.400 -185.500 -177.920 ;
        RECT -176.500 -178.400 -175.580 -177.920 ;
        RECT -166.580 -178.400 -165.660 -177.920 ;
        RECT -156.660 -178.400 -155.740 -177.920 ;
        RECT -146.740 -178.400 -145.820 -177.920 ;
        RECT -136.820 -178.400 -135.900 -177.920 ;
        RECT -126.900 -178.400 -125.980 -177.920 ;
        RECT -116.980 -178.400 -116.060 -177.920 ;
        RECT -107.060 -178.400 -106.140 -177.920 ;
        RECT -97.140 -178.400 -96.220 -177.920 ;
        RECT -87.220 -178.400 -86.300 -177.920 ;
        RECT -77.300 -178.400 -76.380 -177.920 ;
        RECT -67.380 -178.400 -66.460 -177.920 ;
        RECT -57.460 -178.400 -56.540 -177.920 ;
        RECT -47.540 -178.400 -46.620 -177.920 ;
        RECT -37.620 -178.400 -36.700 -177.920 ;
        RECT -27.700 -178.400 -26.780 -177.920 ;
        RECT -17.780 -178.400 -16.860 -177.920 ;
        RECT -7.860 -178.400 -6.940 -177.920 ;
        RECT 2.060 -178.400 2.980 -177.920 ;
        RECT 11.980 -178.400 12.900 -177.920 ;
        RECT 21.900 -178.400 22.820 -177.920 ;
        RECT -278.200 -179.380 -277.030 -178.580 ;
        RECT -268.280 -179.380 -267.110 -178.580 ;
        RECT -258.360 -179.380 -257.190 -178.580 ;
        RECT -248.440 -179.380 -247.270 -178.580 ;
        RECT -238.520 -179.380 -237.350 -178.580 ;
        RECT -228.600 -179.380 -227.430 -178.580 ;
        RECT -218.680 -179.380 -217.510 -178.580 ;
        RECT -208.760 -179.380 -207.590 -178.580 ;
        RECT -198.840 -179.380 -197.670 -178.580 ;
        RECT -188.920 -179.380 -187.750 -178.580 ;
        RECT -179.000 -179.380 -177.830 -178.580 ;
        RECT -169.080 -179.380 -167.910 -178.580 ;
        RECT -159.160 -179.380 -157.990 -178.580 ;
        RECT -149.240 -179.380 -148.070 -178.580 ;
        RECT -139.320 -179.380 -138.150 -178.580 ;
        RECT -129.400 -179.380 -128.230 -178.580 ;
        RECT -119.480 -179.380 -118.310 -178.580 ;
        RECT -109.560 -179.380 -108.390 -178.580 ;
        RECT -99.640 -179.380 -98.470 -178.580 ;
        RECT -89.720 -179.380 -88.550 -178.580 ;
        RECT -79.800 -179.380 -78.630 -178.580 ;
        RECT -69.880 -179.380 -68.710 -178.580 ;
        RECT -59.960 -179.380 -58.790 -178.580 ;
        RECT -50.040 -179.380 -48.870 -178.580 ;
        RECT -40.120 -179.380 -38.950 -178.580 ;
        RECT -30.200 -179.380 -29.030 -178.580 ;
        RECT -20.280 -179.380 -19.110 -178.580 ;
        RECT -10.360 -179.380 -9.190 -178.580 ;
        RECT -0.440 -179.380 0.730 -178.580 ;
        RECT 9.480 -179.380 10.650 -178.580 ;
        RECT 19.400 -179.380 20.570 -178.580 ;
      LAYER via2 ;
        RECT -287.705 94.060 -287.425 94.340 ;
        RECT -277.785 94.060 -277.505 94.340 ;
        RECT -267.865 94.060 -267.585 94.340 ;
        RECT -257.945 94.060 -257.665 94.340 ;
        RECT -248.025 94.060 -247.745 94.340 ;
        RECT -238.105 94.060 -237.825 94.340 ;
        RECT -228.185 94.060 -227.905 94.340 ;
        RECT -218.265 94.060 -217.985 94.340 ;
        RECT -208.345 94.060 -208.065 94.340 ;
        RECT -198.425 94.060 -198.145 94.340 ;
        RECT -188.505 94.060 -188.225 94.340 ;
        RECT -178.585 94.060 -178.305 94.340 ;
        RECT -168.665 94.060 -168.385 94.340 ;
        RECT -158.745 94.060 -158.465 94.340 ;
        RECT -148.825 94.060 -148.545 94.340 ;
        RECT -138.905 94.060 -138.625 94.340 ;
        RECT -128.985 94.060 -128.705 94.340 ;
        RECT -119.065 94.060 -118.785 94.340 ;
        RECT -109.145 94.060 -108.865 94.340 ;
        RECT -99.225 94.060 -98.945 94.340 ;
        RECT -89.305 94.060 -89.025 94.340 ;
        RECT -79.385 94.060 -79.105 94.340 ;
        RECT -69.465 94.060 -69.185 94.340 ;
        RECT -59.545 94.060 -59.265 94.340 ;
        RECT -49.625 94.060 -49.345 94.340 ;
        RECT -39.705 94.060 -39.425 94.340 ;
        RECT -29.785 94.060 -29.505 94.340 ;
        RECT -19.865 94.060 -19.585 94.340 ;
        RECT -9.945 94.060 -9.665 94.340 ;
        RECT -0.025 94.060 0.255 94.340 ;
        RECT 9.895 94.060 10.175 94.340 ;
        RECT 19.815 94.060 20.095 94.340 ;
        RECT -280.535 93.190 -280.255 93.470 ;
        RECT -280.065 93.190 -279.785 93.470 ;
        RECT -270.615 93.190 -270.335 93.470 ;
        RECT -270.145 93.190 -269.865 93.470 ;
        RECT -260.695 93.190 -260.415 93.470 ;
        RECT -260.225 93.190 -259.945 93.470 ;
        RECT -250.775 93.190 -250.495 93.470 ;
        RECT -250.305 93.190 -250.025 93.470 ;
        RECT -240.855 93.190 -240.575 93.470 ;
        RECT -240.385 93.190 -240.105 93.470 ;
        RECT -230.935 93.190 -230.655 93.470 ;
        RECT -230.465 93.190 -230.185 93.470 ;
        RECT -221.015 93.190 -220.735 93.470 ;
        RECT -220.545 93.190 -220.265 93.470 ;
        RECT -211.095 93.190 -210.815 93.470 ;
        RECT -210.625 93.190 -210.345 93.470 ;
        RECT -201.175 93.190 -200.895 93.470 ;
        RECT -200.705 93.190 -200.425 93.470 ;
        RECT -191.255 93.190 -190.975 93.470 ;
        RECT -190.785 93.190 -190.505 93.470 ;
        RECT -181.335 93.190 -181.055 93.470 ;
        RECT -180.865 93.190 -180.585 93.470 ;
        RECT -171.415 93.190 -171.135 93.470 ;
        RECT -170.945 93.190 -170.665 93.470 ;
        RECT -161.495 93.190 -161.215 93.470 ;
        RECT -161.025 93.190 -160.745 93.470 ;
        RECT -151.575 93.190 -151.295 93.470 ;
        RECT -151.105 93.190 -150.825 93.470 ;
        RECT -141.655 93.190 -141.375 93.470 ;
        RECT -141.185 93.190 -140.905 93.470 ;
        RECT -131.735 93.190 -131.455 93.470 ;
        RECT -131.265 93.190 -130.985 93.470 ;
        RECT -121.815 93.190 -121.535 93.470 ;
        RECT -121.345 93.190 -121.065 93.470 ;
        RECT -111.895 93.190 -111.615 93.470 ;
        RECT -111.425 93.190 -111.145 93.470 ;
        RECT -101.975 93.190 -101.695 93.470 ;
        RECT -101.505 93.190 -101.225 93.470 ;
        RECT -92.055 93.190 -91.775 93.470 ;
        RECT -91.585 93.190 -91.305 93.470 ;
        RECT -82.135 93.190 -81.855 93.470 ;
        RECT -81.665 93.190 -81.385 93.470 ;
        RECT -72.215 93.190 -71.935 93.470 ;
        RECT -71.745 93.190 -71.465 93.470 ;
        RECT -62.295 93.190 -62.015 93.470 ;
        RECT -61.825 93.190 -61.545 93.470 ;
        RECT -52.375 93.190 -52.095 93.470 ;
        RECT -51.905 93.190 -51.625 93.470 ;
        RECT -42.455 93.190 -42.175 93.470 ;
        RECT -41.985 93.190 -41.705 93.470 ;
        RECT -32.535 93.190 -32.255 93.470 ;
        RECT -32.065 93.190 -31.785 93.470 ;
        RECT -22.615 93.190 -22.335 93.470 ;
        RECT -22.145 93.190 -21.865 93.470 ;
        RECT -12.695 93.190 -12.415 93.470 ;
        RECT -12.225 93.190 -11.945 93.470 ;
        RECT -2.775 93.190 -2.495 93.470 ;
        RECT -2.305 93.190 -2.025 93.470 ;
        RECT 7.145 93.190 7.425 93.470 ;
        RECT 7.615 93.190 7.895 93.470 ;
        RECT 17.065 93.190 17.345 93.470 ;
        RECT 17.535 93.190 17.815 93.470 ;
        RECT -287.795 90.460 -287.515 90.740 ;
        RECT -287.335 90.470 -287.055 90.750 ;
        RECT -277.875 90.460 -277.595 90.740 ;
        RECT -277.415 90.470 -277.135 90.750 ;
        RECT -267.955 90.460 -267.675 90.740 ;
        RECT -267.495 90.470 -267.215 90.750 ;
        RECT -258.035 90.460 -257.755 90.740 ;
        RECT -257.575 90.470 -257.295 90.750 ;
        RECT -248.115 90.460 -247.835 90.740 ;
        RECT -247.655 90.470 -247.375 90.750 ;
        RECT -238.195 90.460 -237.915 90.740 ;
        RECT -237.735 90.470 -237.455 90.750 ;
        RECT -228.275 90.460 -227.995 90.740 ;
        RECT -227.815 90.470 -227.535 90.750 ;
        RECT -218.355 90.460 -218.075 90.740 ;
        RECT -217.895 90.470 -217.615 90.750 ;
        RECT -208.435 90.460 -208.155 90.740 ;
        RECT -207.975 90.470 -207.695 90.750 ;
        RECT -198.515 90.460 -198.235 90.740 ;
        RECT -198.055 90.470 -197.775 90.750 ;
        RECT -188.595 90.460 -188.315 90.740 ;
        RECT -188.135 90.470 -187.855 90.750 ;
        RECT -178.675 90.460 -178.395 90.740 ;
        RECT -178.215 90.470 -177.935 90.750 ;
        RECT -168.755 90.460 -168.475 90.740 ;
        RECT -168.295 90.470 -168.015 90.750 ;
        RECT -158.835 90.460 -158.555 90.740 ;
        RECT -158.375 90.470 -158.095 90.750 ;
        RECT -148.915 90.460 -148.635 90.740 ;
        RECT -148.455 90.470 -148.175 90.750 ;
        RECT -138.995 90.460 -138.715 90.740 ;
        RECT -138.535 90.470 -138.255 90.750 ;
        RECT -129.075 90.460 -128.795 90.740 ;
        RECT -128.615 90.470 -128.335 90.750 ;
        RECT -119.155 90.460 -118.875 90.740 ;
        RECT -118.695 90.470 -118.415 90.750 ;
        RECT -109.235 90.460 -108.955 90.740 ;
        RECT -108.775 90.470 -108.495 90.750 ;
        RECT -99.315 90.460 -99.035 90.740 ;
        RECT -98.855 90.470 -98.575 90.750 ;
        RECT -89.395 90.460 -89.115 90.740 ;
        RECT -88.935 90.470 -88.655 90.750 ;
        RECT -79.475 90.460 -79.195 90.740 ;
        RECT -79.015 90.470 -78.735 90.750 ;
        RECT -69.555 90.460 -69.275 90.740 ;
        RECT -69.095 90.470 -68.815 90.750 ;
        RECT -59.635 90.460 -59.355 90.740 ;
        RECT -59.175 90.470 -58.895 90.750 ;
        RECT -49.715 90.460 -49.435 90.740 ;
        RECT -49.255 90.470 -48.975 90.750 ;
        RECT -39.795 90.460 -39.515 90.740 ;
        RECT -39.335 90.470 -39.055 90.750 ;
        RECT -29.875 90.460 -29.595 90.740 ;
        RECT -29.415 90.470 -29.135 90.750 ;
        RECT -19.955 90.460 -19.675 90.740 ;
        RECT -19.495 90.470 -19.215 90.750 ;
        RECT -10.035 90.460 -9.755 90.740 ;
        RECT -9.575 90.470 -9.295 90.750 ;
        RECT -0.115 90.460 0.165 90.740 ;
        RECT 0.345 90.470 0.625 90.750 ;
        RECT 9.805 90.460 10.085 90.740 ;
        RECT 10.265 90.470 10.545 90.750 ;
        RECT 19.725 90.460 20.005 90.740 ;
        RECT 20.185 90.470 20.465 90.750 ;
        RECT -280.145 89.700 -279.865 89.980 ;
        RECT -270.225 89.700 -269.945 89.980 ;
        RECT -260.305 89.700 -260.025 89.980 ;
        RECT -250.385 89.700 -250.105 89.980 ;
        RECT -240.465 89.700 -240.185 89.980 ;
        RECT -230.545 89.700 -230.265 89.980 ;
        RECT -220.625 89.700 -220.345 89.980 ;
        RECT -210.705 89.700 -210.425 89.980 ;
        RECT -200.785 89.700 -200.505 89.980 ;
        RECT -190.865 89.700 -190.585 89.980 ;
        RECT -180.945 89.700 -180.665 89.980 ;
        RECT -171.025 89.700 -170.745 89.980 ;
        RECT -161.105 89.700 -160.825 89.980 ;
        RECT -151.185 89.700 -150.905 89.980 ;
        RECT -141.265 89.700 -140.985 89.980 ;
        RECT -131.345 89.700 -131.065 89.980 ;
        RECT -121.425 89.700 -121.145 89.980 ;
        RECT -111.505 89.700 -111.225 89.980 ;
        RECT -101.585 89.700 -101.305 89.980 ;
        RECT -91.665 89.700 -91.385 89.980 ;
        RECT -81.745 89.700 -81.465 89.980 ;
        RECT -71.825 89.700 -71.545 89.980 ;
        RECT -61.905 89.700 -61.625 89.980 ;
        RECT -51.985 89.700 -51.705 89.980 ;
        RECT -42.065 89.700 -41.785 89.980 ;
        RECT -32.145 89.700 -31.865 89.980 ;
        RECT -22.225 89.700 -21.945 89.980 ;
        RECT -12.305 89.700 -12.025 89.980 ;
        RECT -2.385 89.700 -2.105 89.980 ;
        RECT 7.535 89.700 7.815 89.980 ;
        RECT 17.455 89.700 17.735 89.980 ;
        RECT -287.455 6.350 -287.175 6.630 ;
        RECT -277.535 6.350 -277.255 6.630 ;
        RECT -267.615 6.350 -267.335 6.630 ;
        RECT -257.695 6.350 -257.415 6.630 ;
        RECT -247.775 6.350 -247.495 6.630 ;
        RECT -237.855 6.350 -237.575 6.630 ;
        RECT -227.935 6.350 -227.655 6.630 ;
        RECT -218.015 6.350 -217.735 6.630 ;
        RECT -208.095 6.350 -207.815 6.630 ;
        RECT -198.175 6.350 -197.895 6.630 ;
        RECT -188.255 6.350 -187.975 6.630 ;
        RECT -178.335 6.350 -178.055 6.630 ;
        RECT -168.415 6.350 -168.135 6.630 ;
        RECT -158.495 6.350 -158.215 6.630 ;
        RECT -148.575 6.350 -148.295 6.630 ;
        RECT -138.655 6.350 -138.375 6.630 ;
        RECT -128.735 6.350 -128.455 6.630 ;
        RECT -118.815 6.350 -118.535 6.630 ;
        RECT -108.895 6.350 -108.615 6.630 ;
        RECT -98.975 6.350 -98.695 6.630 ;
        RECT -89.055 6.350 -88.775 6.630 ;
        RECT -79.135 6.350 -78.855 6.630 ;
        RECT -69.215 6.350 -68.935 6.630 ;
        RECT -59.295 6.350 -59.015 6.630 ;
        RECT -49.375 6.350 -49.095 6.630 ;
        RECT -39.455 6.350 -39.175 6.630 ;
        RECT -29.535 6.350 -29.255 6.630 ;
        RECT -19.615 6.350 -19.335 6.630 ;
        RECT -9.695 6.350 -9.415 6.630 ;
        RECT 0.225 6.350 0.505 6.630 ;
        RECT 10.145 6.350 10.425 6.630 ;
        RECT 20.065 6.350 20.345 6.630 ;
        RECT -280.285 5.480 -280.005 5.760 ;
        RECT -279.815 5.480 -279.535 5.760 ;
        RECT -270.365 5.480 -270.085 5.760 ;
        RECT -269.895 5.480 -269.615 5.760 ;
        RECT -260.445 5.480 -260.165 5.760 ;
        RECT -259.975 5.480 -259.695 5.760 ;
        RECT -250.525 5.480 -250.245 5.760 ;
        RECT -250.055 5.480 -249.775 5.760 ;
        RECT -240.605 5.480 -240.325 5.760 ;
        RECT -240.135 5.480 -239.855 5.760 ;
        RECT -230.685 5.480 -230.405 5.760 ;
        RECT -230.215 5.480 -229.935 5.760 ;
        RECT -220.765 5.480 -220.485 5.760 ;
        RECT -220.295 5.480 -220.015 5.760 ;
        RECT -210.845 5.480 -210.565 5.760 ;
        RECT -210.375 5.480 -210.095 5.760 ;
        RECT -200.925 5.480 -200.645 5.760 ;
        RECT -200.455 5.480 -200.175 5.760 ;
        RECT -191.005 5.480 -190.725 5.760 ;
        RECT -190.535 5.480 -190.255 5.760 ;
        RECT -181.085 5.480 -180.805 5.760 ;
        RECT -180.615 5.480 -180.335 5.760 ;
        RECT -171.165 5.480 -170.885 5.760 ;
        RECT -170.695 5.480 -170.415 5.760 ;
        RECT -161.245 5.480 -160.965 5.760 ;
        RECT -160.775 5.480 -160.495 5.760 ;
        RECT -151.325 5.480 -151.045 5.760 ;
        RECT -150.855 5.480 -150.575 5.760 ;
        RECT -141.405 5.480 -141.125 5.760 ;
        RECT -140.935 5.480 -140.655 5.760 ;
        RECT -131.485 5.480 -131.205 5.760 ;
        RECT -131.015 5.480 -130.735 5.760 ;
        RECT -121.565 5.480 -121.285 5.760 ;
        RECT -121.095 5.480 -120.815 5.760 ;
        RECT -111.645 5.480 -111.365 5.760 ;
        RECT -111.175 5.480 -110.895 5.760 ;
        RECT -101.725 5.480 -101.445 5.760 ;
        RECT -101.255 5.480 -100.975 5.760 ;
        RECT -91.805 5.480 -91.525 5.760 ;
        RECT -91.335 5.480 -91.055 5.760 ;
        RECT -81.885 5.480 -81.605 5.760 ;
        RECT -81.415 5.480 -81.135 5.760 ;
        RECT -71.965 5.480 -71.685 5.760 ;
        RECT -71.495 5.480 -71.215 5.760 ;
        RECT -62.045 5.480 -61.765 5.760 ;
        RECT -61.575 5.480 -61.295 5.760 ;
        RECT -52.125 5.480 -51.845 5.760 ;
        RECT -51.655 5.480 -51.375 5.760 ;
        RECT -42.205 5.480 -41.925 5.760 ;
        RECT -41.735 5.480 -41.455 5.760 ;
        RECT -32.285 5.480 -32.005 5.760 ;
        RECT -31.815 5.480 -31.535 5.760 ;
        RECT -22.365 5.480 -22.085 5.760 ;
        RECT -21.895 5.480 -21.615 5.760 ;
        RECT -12.445 5.480 -12.165 5.760 ;
        RECT -11.975 5.480 -11.695 5.760 ;
        RECT -2.525 5.480 -2.245 5.760 ;
        RECT -2.055 5.480 -1.775 5.760 ;
        RECT 7.395 5.480 7.675 5.760 ;
        RECT 7.865 5.480 8.145 5.760 ;
        RECT 17.315 5.480 17.595 5.760 ;
        RECT 17.785 5.480 18.065 5.760 ;
        RECT -287.545 2.750 -287.265 3.030 ;
        RECT -287.085 2.760 -286.805 3.040 ;
        RECT -277.625 2.750 -277.345 3.030 ;
        RECT -277.165 2.760 -276.885 3.040 ;
        RECT -267.705 2.750 -267.425 3.030 ;
        RECT -267.245 2.760 -266.965 3.040 ;
        RECT -257.785 2.750 -257.505 3.030 ;
        RECT -257.325 2.760 -257.045 3.040 ;
        RECT -247.865 2.750 -247.585 3.030 ;
        RECT -247.405 2.760 -247.125 3.040 ;
        RECT -237.945 2.750 -237.665 3.030 ;
        RECT -237.485 2.760 -237.205 3.040 ;
        RECT -228.025 2.750 -227.745 3.030 ;
        RECT -227.565 2.760 -227.285 3.040 ;
        RECT -218.105 2.750 -217.825 3.030 ;
        RECT -217.645 2.760 -217.365 3.040 ;
        RECT -208.185 2.750 -207.905 3.030 ;
        RECT -207.725 2.760 -207.445 3.040 ;
        RECT -198.265 2.750 -197.985 3.030 ;
        RECT -197.805 2.760 -197.525 3.040 ;
        RECT -188.345 2.750 -188.065 3.030 ;
        RECT -187.885 2.760 -187.605 3.040 ;
        RECT -178.425 2.750 -178.145 3.030 ;
        RECT -177.965 2.760 -177.685 3.040 ;
        RECT -168.505 2.750 -168.225 3.030 ;
        RECT -168.045 2.760 -167.765 3.040 ;
        RECT -158.585 2.750 -158.305 3.030 ;
        RECT -158.125 2.760 -157.845 3.040 ;
        RECT -148.665 2.750 -148.385 3.030 ;
        RECT -148.205 2.760 -147.925 3.040 ;
        RECT -138.745 2.750 -138.465 3.030 ;
        RECT -138.285 2.760 -138.005 3.040 ;
        RECT -128.825 2.750 -128.545 3.030 ;
        RECT -128.365 2.760 -128.085 3.040 ;
        RECT -118.905 2.750 -118.625 3.030 ;
        RECT -118.445 2.760 -118.165 3.040 ;
        RECT -108.985 2.750 -108.705 3.030 ;
        RECT -108.525 2.760 -108.245 3.040 ;
        RECT -99.065 2.750 -98.785 3.030 ;
        RECT -98.605 2.760 -98.325 3.040 ;
        RECT -89.145 2.750 -88.865 3.030 ;
        RECT -88.685 2.760 -88.405 3.040 ;
        RECT -79.225 2.750 -78.945 3.030 ;
        RECT -78.765 2.760 -78.485 3.040 ;
        RECT -69.305 2.750 -69.025 3.030 ;
        RECT -68.845 2.760 -68.565 3.040 ;
        RECT -59.385 2.750 -59.105 3.030 ;
        RECT -58.925 2.760 -58.645 3.040 ;
        RECT -49.465 2.750 -49.185 3.030 ;
        RECT -49.005 2.760 -48.725 3.040 ;
        RECT -39.545 2.750 -39.265 3.030 ;
        RECT -39.085 2.760 -38.805 3.040 ;
        RECT -29.625 2.750 -29.345 3.030 ;
        RECT -29.165 2.760 -28.885 3.040 ;
        RECT -19.705 2.750 -19.425 3.030 ;
        RECT -19.245 2.760 -18.965 3.040 ;
        RECT -9.785 2.750 -9.505 3.030 ;
        RECT -9.325 2.760 -9.045 3.040 ;
        RECT 0.135 2.750 0.415 3.030 ;
        RECT 0.595 2.760 0.875 3.040 ;
        RECT 10.055 2.750 10.335 3.030 ;
        RECT 10.515 2.760 10.795 3.040 ;
        RECT 19.975 2.750 20.255 3.030 ;
        RECT 20.435 2.760 20.715 3.040 ;
        RECT -279.895 1.990 -279.615 2.270 ;
        RECT -269.975 1.990 -269.695 2.270 ;
        RECT -260.055 1.990 -259.775 2.270 ;
        RECT -250.135 1.990 -249.855 2.270 ;
        RECT -240.215 1.990 -239.935 2.270 ;
        RECT -230.295 1.990 -230.015 2.270 ;
        RECT -220.375 1.990 -220.095 2.270 ;
        RECT -210.455 1.990 -210.175 2.270 ;
        RECT -200.535 1.990 -200.255 2.270 ;
        RECT -190.615 1.990 -190.335 2.270 ;
        RECT -180.695 1.990 -180.415 2.270 ;
        RECT -170.775 1.990 -170.495 2.270 ;
        RECT -160.855 1.990 -160.575 2.270 ;
        RECT -150.935 1.990 -150.655 2.270 ;
        RECT -141.015 1.990 -140.735 2.270 ;
        RECT -131.095 1.990 -130.815 2.270 ;
        RECT -121.175 1.990 -120.895 2.270 ;
        RECT -111.255 1.990 -110.975 2.270 ;
        RECT -101.335 1.990 -101.055 2.270 ;
        RECT -91.415 1.990 -91.135 2.270 ;
        RECT -81.495 1.990 -81.215 2.270 ;
        RECT -71.575 1.990 -71.295 2.270 ;
        RECT -61.655 1.990 -61.375 2.270 ;
        RECT -51.735 1.990 -51.455 2.270 ;
        RECT -41.815 1.990 -41.535 2.270 ;
        RECT -31.895 1.990 -31.615 2.270 ;
        RECT -21.975 1.990 -21.695 2.270 ;
        RECT -12.055 1.990 -11.775 2.270 ;
        RECT -2.135 1.990 -1.855 2.270 ;
        RECT 7.785 1.990 8.065 2.270 ;
        RECT 17.705 1.990 17.985 2.270 ;
        RECT -285.695 -87.000 -285.415 -86.720 ;
        RECT -275.775 -87.000 -275.495 -86.720 ;
        RECT -265.855 -87.000 -265.575 -86.720 ;
        RECT -255.935 -87.000 -255.655 -86.720 ;
        RECT -246.015 -87.000 -245.735 -86.720 ;
        RECT -236.095 -87.000 -235.815 -86.720 ;
        RECT -226.175 -87.000 -225.895 -86.720 ;
        RECT -216.255 -87.000 -215.975 -86.720 ;
        RECT -206.335 -87.000 -206.055 -86.720 ;
        RECT -196.415 -87.000 -196.135 -86.720 ;
        RECT -186.495 -87.000 -186.215 -86.720 ;
        RECT -176.575 -87.000 -176.295 -86.720 ;
        RECT -166.655 -87.000 -166.375 -86.720 ;
        RECT -156.735 -87.000 -156.455 -86.720 ;
        RECT -146.815 -87.000 -146.535 -86.720 ;
        RECT -136.895 -87.000 -136.615 -86.720 ;
        RECT -126.975 -87.000 -126.695 -86.720 ;
        RECT -117.055 -87.000 -116.775 -86.720 ;
        RECT -107.135 -87.000 -106.855 -86.720 ;
        RECT -97.215 -87.000 -96.935 -86.720 ;
        RECT -87.295 -87.000 -87.015 -86.720 ;
        RECT -77.375 -87.000 -77.095 -86.720 ;
        RECT -67.455 -87.000 -67.175 -86.720 ;
        RECT -57.535 -87.000 -57.255 -86.720 ;
        RECT -47.615 -87.000 -47.335 -86.720 ;
        RECT -37.695 -87.000 -37.415 -86.720 ;
        RECT -27.775 -87.000 -27.495 -86.720 ;
        RECT -17.855 -87.000 -17.575 -86.720 ;
        RECT -7.935 -87.000 -7.655 -86.720 ;
        RECT 1.985 -87.000 2.265 -86.720 ;
        RECT 11.905 -87.000 12.185 -86.720 ;
        RECT 21.825 -87.000 22.105 -86.720 ;
        RECT -278.525 -87.870 -278.245 -87.590 ;
        RECT -278.055 -87.870 -277.775 -87.590 ;
        RECT -268.605 -87.870 -268.325 -87.590 ;
        RECT -268.135 -87.870 -267.855 -87.590 ;
        RECT -258.685 -87.870 -258.405 -87.590 ;
        RECT -258.215 -87.870 -257.935 -87.590 ;
        RECT -248.765 -87.870 -248.485 -87.590 ;
        RECT -248.295 -87.870 -248.015 -87.590 ;
        RECT -238.845 -87.870 -238.565 -87.590 ;
        RECT -238.375 -87.870 -238.095 -87.590 ;
        RECT -228.925 -87.870 -228.645 -87.590 ;
        RECT -228.455 -87.870 -228.175 -87.590 ;
        RECT -219.005 -87.870 -218.725 -87.590 ;
        RECT -218.535 -87.870 -218.255 -87.590 ;
        RECT -209.085 -87.870 -208.805 -87.590 ;
        RECT -208.615 -87.870 -208.335 -87.590 ;
        RECT -199.165 -87.870 -198.885 -87.590 ;
        RECT -198.695 -87.870 -198.415 -87.590 ;
        RECT -189.245 -87.870 -188.965 -87.590 ;
        RECT -188.775 -87.870 -188.495 -87.590 ;
        RECT -179.325 -87.870 -179.045 -87.590 ;
        RECT -178.855 -87.870 -178.575 -87.590 ;
        RECT -169.405 -87.870 -169.125 -87.590 ;
        RECT -168.935 -87.870 -168.655 -87.590 ;
        RECT -159.485 -87.870 -159.205 -87.590 ;
        RECT -159.015 -87.870 -158.735 -87.590 ;
        RECT -149.565 -87.870 -149.285 -87.590 ;
        RECT -149.095 -87.870 -148.815 -87.590 ;
        RECT -139.645 -87.870 -139.365 -87.590 ;
        RECT -139.175 -87.870 -138.895 -87.590 ;
        RECT -129.725 -87.870 -129.445 -87.590 ;
        RECT -129.255 -87.870 -128.975 -87.590 ;
        RECT -119.805 -87.870 -119.525 -87.590 ;
        RECT -119.335 -87.870 -119.055 -87.590 ;
        RECT -109.885 -87.870 -109.605 -87.590 ;
        RECT -109.415 -87.870 -109.135 -87.590 ;
        RECT -99.965 -87.870 -99.685 -87.590 ;
        RECT -99.495 -87.870 -99.215 -87.590 ;
        RECT -90.045 -87.870 -89.765 -87.590 ;
        RECT -89.575 -87.870 -89.295 -87.590 ;
        RECT -80.125 -87.870 -79.845 -87.590 ;
        RECT -79.655 -87.870 -79.375 -87.590 ;
        RECT -70.205 -87.870 -69.925 -87.590 ;
        RECT -69.735 -87.870 -69.455 -87.590 ;
        RECT -60.285 -87.870 -60.005 -87.590 ;
        RECT -59.815 -87.870 -59.535 -87.590 ;
        RECT -50.365 -87.870 -50.085 -87.590 ;
        RECT -49.895 -87.870 -49.615 -87.590 ;
        RECT -40.445 -87.870 -40.165 -87.590 ;
        RECT -39.975 -87.870 -39.695 -87.590 ;
        RECT -30.525 -87.870 -30.245 -87.590 ;
        RECT -30.055 -87.870 -29.775 -87.590 ;
        RECT -20.605 -87.870 -20.325 -87.590 ;
        RECT -20.135 -87.870 -19.855 -87.590 ;
        RECT -10.685 -87.870 -10.405 -87.590 ;
        RECT -10.215 -87.870 -9.935 -87.590 ;
        RECT -0.765 -87.870 -0.485 -87.590 ;
        RECT -0.295 -87.870 -0.015 -87.590 ;
        RECT 9.155 -87.870 9.435 -87.590 ;
        RECT 9.625 -87.870 9.905 -87.590 ;
        RECT 19.075 -87.870 19.355 -87.590 ;
        RECT 19.545 -87.870 19.825 -87.590 ;
        RECT -285.785 -90.600 -285.505 -90.320 ;
        RECT -285.325 -90.590 -285.045 -90.310 ;
        RECT -275.865 -90.600 -275.585 -90.320 ;
        RECT -275.405 -90.590 -275.125 -90.310 ;
        RECT -265.945 -90.600 -265.665 -90.320 ;
        RECT -265.485 -90.590 -265.205 -90.310 ;
        RECT -256.025 -90.600 -255.745 -90.320 ;
        RECT -255.565 -90.590 -255.285 -90.310 ;
        RECT -246.105 -90.600 -245.825 -90.320 ;
        RECT -245.645 -90.590 -245.365 -90.310 ;
        RECT -236.185 -90.600 -235.905 -90.320 ;
        RECT -235.725 -90.590 -235.445 -90.310 ;
        RECT -226.265 -90.600 -225.985 -90.320 ;
        RECT -225.805 -90.590 -225.525 -90.310 ;
        RECT -216.345 -90.600 -216.065 -90.320 ;
        RECT -215.885 -90.590 -215.605 -90.310 ;
        RECT -206.425 -90.600 -206.145 -90.320 ;
        RECT -205.965 -90.590 -205.685 -90.310 ;
        RECT -196.505 -90.600 -196.225 -90.320 ;
        RECT -196.045 -90.590 -195.765 -90.310 ;
        RECT -186.585 -90.600 -186.305 -90.320 ;
        RECT -186.125 -90.590 -185.845 -90.310 ;
        RECT -176.665 -90.600 -176.385 -90.320 ;
        RECT -176.205 -90.590 -175.925 -90.310 ;
        RECT -166.745 -90.600 -166.465 -90.320 ;
        RECT -166.285 -90.590 -166.005 -90.310 ;
        RECT -156.825 -90.600 -156.545 -90.320 ;
        RECT -156.365 -90.590 -156.085 -90.310 ;
        RECT -146.905 -90.600 -146.625 -90.320 ;
        RECT -146.445 -90.590 -146.165 -90.310 ;
        RECT -136.985 -90.600 -136.705 -90.320 ;
        RECT -136.525 -90.590 -136.245 -90.310 ;
        RECT -127.065 -90.600 -126.785 -90.320 ;
        RECT -126.605 -90.590 -126.325 -90.310 ;
        RECT -117.145 -90.600 -116.865 -90.320 ;
        RECT -116.685 -90.590 -116.405 -90.310 ;
        RECT -107.225 -90.600 -106.945 -90.320 ;
        RECT -106.765 -90.590 -106.485 -90.310 ;
        RECT -97.305 -90.600 -97.025 -90.320 ;
        RECT -96.845 -90.590 -96.565 -90.310 ;
        RECT -87.385 -90.600 -87.105 -90.320 ;
        RECT -86.925 -90.590 -86.645 -90.310 ;
        RECT -77.465 -90.600 -77.185 -90.320 ;
        RECT -77.005 -90.590 -76.725 -90.310 ;
        RECT -67.545 -90.600 -67.265 -90.320 ;
        RECT -67.085 -90.590 -66.805 -90.310 ;
        RECT -57.625 -90.600 -57.345 -90.320 ;
        RECT -57.165 -90.590 -56.885 -90.310 ;
        RECT -47.705 -90.600 -47.425 -90.320 ;
        RECT -47.245 -90.590 -46.965 -90.310 ;
        RECT -37.785 -90.600 -37.505 -90.320 ;
        RECT -37.325 -90.590 -37.045 -90.310 ;
        RECT -27.865 -90.600 -27.585 -90.320 ;
        RECT -27.405 -90.590 -27.125 -90.310 ;
        RECT -17.945 -90.600 -17.665 -90.320 ;
        RECT -17.485 -90.590 -17.205 -90.310 ;
        RECT -8.025 -90.600 -7.745 -90.320 ;
        RECT -7.565 -90.590 -7.285 -90.310 ;
        RECT 1.895 -90.600 2.175 -90.320 ;
        RECT 2.355 -90.590 2.635 -90.310 ;
        RECT 11.815 -90.600 12.095 -90.320 ;
        RECT 12.275 -90.590 12.555 -90.310 ;
        RECT 21.735 -90.600 22.015 -90.320 ;
        RECT 22.195 -90.590 22.475 -90.310 ;
        RECT -278.135 -91.360 -277.855 -91.080 ;
        RECT -268.215 -91.360 -267.935 -91.080 ;
        RECT -258.295 -91.360 -258.015 -91.080 ;
        RECT -248.375 -91.360 -248.095 -91.080 ;
        RECT -238.455 -91.360 -238.175 -91.080 ;
        RECT -228.535 -91.360 -228.255 -91.080 ;
        RECT -218.615 -91.360 -218.335 -91.080 ;
        RECT -208.695 -91.360 -208.415 -91.080 ;
        RECT -198.775 -91.360 -198.495 -91.080 ;
        RECT -188.855 -91.360 -188.575 -91.080 ;
        RECT -178.935 -91.360 -178.655 -91.080 ;
        RECT -169.015 -91.360 -168.735 -91.080 ;
        RECT -159.095 -91.360 -158.815 -91.080 ;
        RECT -149.175 -91.360 -148.895 -91.080 ;
        RECT -139.255 -91.360 -138.975 -91.080 ;
        RECT -129.335 -91.360 -129.055 -91.080 ;
        RECT -119.415 -91.360 -119.135 -91.080 ;
        RECT -109.495 -91.360 -109.215 -91.080 ;
        RECT -99.575 -91.360 -99.295 -91.080 ;
        RECT -89.655 -91.360 -89.375 -91.080 ;
        RECT -79.735 -91.360 -79.455 -91.080 ;
        RECT -69.815 -91.360 -69.535 -91.080 ;
        RECT -59.895 -91.360 -59.615 -91.080 ;
        RECT -49.975 -91.360 -49.695 -91.080 ;
        RECT -40.055 -91.360 -39.775 -91.080 ;
        RECT -30.135 -91.360 -29.855 -91.080 ;
        RECT -20.215 -91.360 -19.935 -91.080 ;
        RECT -10.295 -91.360 -10.015 -91.080 ;
        RECT -0.375 -91.360 -0.095 -91.080 ;
        RECT 9.545 -91.360 9.825 -91.080 ;
        RECT 19.465 -91.360 19.745 -91.080 ;
        RECT -285.445 -174.710 -285.165 -174.430 ;
        RECT -275.525 -174.710 -275.245 -174.430 ;
        RECT -265.605 -174.710 -265.325 -174.430 ;
        RECT -255.685 -174.710 -255.405 -174.430 ;
        RECT -245.765 -174.710 -245.485 -174.430 ;
        RECT -235.845 -174.710 -235.565 -174.430 ;
        RECT -225.925 -174.710 -225.645 -174.430 ;
        RECT -216.005 -174.710 -215.725 -174.430 ;
        RECT -206.085 -174.710 -205.805 -174.430 ;
        RECT -196.165 -174.710 -195.885 -174.430 ;
        RECT -186.245 -174.710 -185.965 -174.430 ;
        RECT -176.325 -174.710 -176.045 -174.430 ;
        RECT -166.405 -174.710 -166.125 -174.430 ;
        RECT -156.485 -174.710 -156.205 -174.430 ;
        RECT -146.565 -174.710 -146.285 -174.430 ;
        RECT -136.645 -174.710 -136.365 -174.430 ;
        RECT -126.725 -174.710 -126.445 -174.430 ;
        RECT -116.805 -174.710 -116.525 -174.430 ;
        RECT -106.885 -174.710 -106.605 -174.430 ;
        RECT -96.965 -174.710 -96.685 -174.430 ;
        RECT -87.045 -174.710 -86.765 -174.430 ;
        RECT -77.125 -174.710 -76.845 -174.430 ;
        RECT -67.205 -174.710 -66.925 -174.430 ;
        RECT -57.285 -174.710 -57.005 -174.430 ;
        RECT -47.365 -174.710 -47.085 -174.430 ;
        RECT -37.445 -174.710 -37.165 -174.430 ;
        RECT -27.525 -174.710 -27.245 -174.430 ;
        RECT -17.605 -174.710 -17.325 -174.430 ;
        RECT -7.685 -174.710 -7.405 -174.430 ;
        RECT 2.235 -174.710 2.515 -174.430 ;
        RECT 12.155 -174.710 12.435 -174.430 ;
        RECT 22.075 -174.710 22.355 -174.430 ;
        RECT -278.275 -175.580 -277.995 -175.300 ;
        RECT -277.805 -175.580 -277.525 -175.300 ;
        RECT -268.355 -175.580 -268.075 -175.300 ;
        RECT -267.885 -175.580 -267.605 -175.300 ;
        RECT -258.435 -175.580 -258.155 -175.300 ;
        RECT -257.965 -175.580 -257.685 -175.300 ;
        RECT -248.515 -175.580 -248.235 -175.300 ;
        RECT -248.045 -175.580 -247.765 -175.300 ;
        RECT -238.595 -175.580 -238.315 -175.300 ;
        RECT -238.125 -175.580 -237.845 -175.300 ;
        RECT -228.675 -175.580 -228.395 -175.300 ;
        RECT -228.205 -175.580 -227.925 -175.300 ;
        RECT -218.755 -175.580 -218.475 -175.300 ;
        RECT -218.285 -175.580 -218.005 -175.300 ;
        RECT -208.835 -175.580 -208.555 -175.300 ;
        RECT -208.365 -175.580 -208.085 -175.300 ;
        RECT -198.915 -175.580 -198.635 -175.300 ;
        RECT -198.445 -175.580 -198.165 -175.300 ;
        RECT -188.995 -175.580 -188.715 -175.300 ;
        RECT -188.525 -175.580 -188.245 -175.300 ;
        RECT -179.075 -175.580 -178.795 -175.300 ;
        RECT -178.605 -175.580 -178.325 -175.300 ;
        RECT -169.155 -175.580 -168.875 -175.300 ;
        RECT -168.685 -175.580 -168.405 -175.300 ;
        RECT -159.235 -175.580 -158.955 -175.300 ;
        RECT -158.765 -175.580 -158.485 -175.300 ;
        RECT -149.315 -175.580 -149.035 -175.300 ;
        RECT -148.845 -175.580 -148.565 -175.300 ;
        RECT -139.395 -175.580 -139.115 -175.300 ;
        RECT -138.925 -175.580 -138.645 -175.300 ;
        RECT -129.475 -175.580 -129.195 -175.300 ;
        RECT -129.005 -175.580 -128.725 -175.300 ;
        RECT -119.555 -175.580 -119.275 -175.300 ;
        RECT -119.085 -175.580 -118.805 -175.300 ;
        RECT -109.635 -175.580 -109.355 -175.300 ;
        RECT -109.165 -175.580 -108.885 -175.300 ;
        RECT -99.715 -175.580 -99.435 -175.300 ;
        RECT -99.245 -175.580 -98.965 -175.300 ;
        RECT -89.795 -175.580 -89.515 -175.300 ;
        RECT -89.325 -175.580 -89.045 -175.300 ;
        RECT -79.875 -175.580 -79.595 -175.300 ;
        RECT -79.405 -175.580 -79.125 -175.300 ;
        RECT -69.955 -175.580 -69.675 -175.300 ;
        RECT -69.485 -175.580 -69.205 -175.300 ;
        RECT -60.035 -175.580 -59.755 -175.300 ;
        RECT -59.565 -175.580 -59.285 -175.300 ;
        RECT -50.115 -175.580 -49.835 -175.300 ;
        RECT -49.645 -175.580 -49.365 -175.300 ;
        RECT -40.195 -175.580 -39.915 -175.300 ;
        RECT -39.725 -175.580 -39.445 -175.300 ;
        RECT -30.275 -175.580 -29.995 -175.300 ;
        RECT -29.805 -175.580 -29.525 -175.300 ;
        RECT -20.355 -175.580 -20.075 -175.300 ;
        RECT -19.885 -175.580 -19.605 -175.300 ;
        RECT -10.435 -175.580 -10.155 -175.300 ;
        RECT -9.965 -175.580 -9.685 -175.300 ;
        RECT -0.515 -175.580 -0.235 -175.300 ;
        RECT -0.045 -175.580 0.235 -175.300 ;
        RECT 9.405 -175.580 9.685 -175.300 ;
        RECT 9.875 -175.580 10.155 -175.300 ;
        RECT 19.325 -175.580 19.605 -175.300 ;
        RECT 19.795 -175.580 20.075 -175.300 ;
        RECT -285.535 -178.310 -285.255 -178.030 ;
        RECT -285.075 -178.300 -284.795 -178.020 ;
        RECT -275.615 -178.310 -275.335 -178.030 ;
        RECT -275.155 -178.300 -274.875 -178.020 ;
        RECT -265.695 -178.310 -265.415 -178.030 ;
        RECT -265.235 -178.300 -264.955 -178.020 ;
        RECT -255.775 -178.310 -255.495 -178.030 ;
        RECT -255.315 -178.300 -255.035 -178.020 ;
        RECT -245.855 -178.310 -245.575 -178.030 ;
        RECT -245.395 -178.300 -245.115 -178.020 ;
        RECT -235.935 -178.310 -235.655 -178.030 ;
        RECT -235.475 -178.300 -235.195 -178.020 ;
        RECT -226.015 -178.310 -225.735 -178.030 ;
        RECT -225.555 -178.300 -225.275 -178.020 ;
        RECT -216.095 -178.310 -215.815 -178.030 ;
        RECT -215.635 -178.300 -215.355 -178.020 ;
        RECT -206.175 -178.310 -205.895 -178.030 ;
        RECT -205.715 -178.300 -205.435 -178.020 ;
        RECT -196.255 -178.310 -195.975 -178.030 ;
        RECT -195.795 -178.300 -195.515 -178.020 ;
        RECT -186.335 -178.310 -186.055 -178.030 ;
        RECT -185.875 -178.300 -185.595 -178.020 ;
        RECT -176.415 -178.310 -176.135 -178.030 ;
        RECT -175.955 -178.300 -175.675 -178.020 ;
        RECT -166.495 -178.310 -166.215 -178.030 ;
        RECT -166.035 -178.300 -165.755 -178.020 ;
        RECT -156.575 -178.310 -156.295 -178.030 ;
        RECT -156.115 -178.300 -155.835 -178.020 ;
        RECT -146.655 -178.310 -146.375 -178.030 ;
        RECT -146.195 -178.300 -145.915 -178.020 ;
        RECT -136.735 -178.310 -136.455 -178.030 ;
        RECT -136.275 -178.300 -135.995 -178.020 ;
        RECT -126.815 -178.310 -126.535 -178.030 ;
        RECT -126.355 -178.300 -126.075 -178.020 ;
        RECT -116.895 -178.310 -116.615 -178.030 ;
        RECT -116.435 -178.300 -116.155 -178.020 ;
        RECT -106.975 -178.310 -106.695 -178.030 ;
        RECT -106.515 -178.300 -106.235 -178.020 ;
        RECT -97.055 -178.310 -96.775 -178.030 ;
        RECT -96.595 -178.300 -96.315 -178.020 ;
        RECT -87.135 -178.310 -86.855 -178.030 ;
        RECT -86.675 -178.300 -86.395 -178.020 ;
        RECT -77.215 -178.310 -76.935 -178.030 ;
        RECT -76.755 -178.300 -76.475 -178.020 ;
        RECT -67.295 -178.310 -67.015 -178.030 ;
        RECT -66.835 -178.300 -66.555 -178.020 ;
        RECT -57.375 -178.310 -57.095 -178.030 ;
        RECT -56.915 -178.300 -56.635 -178.020 ;
        RECT -47.455 -178.310 -47.175 -178.030 ;
        RECT -46.995 -178.300 -46.715 -178.020 ;
        RECT -37.535 -178.310 -37.255 -178.030 ;
        RECT -37.075 -178.300 -36.795 -178.020 ;
        RECT -27.615 -178.310 -27.335 -178.030 ;
        RECT -27.155 -178.300 -26.875 -178.020 ;
        RECT -17.695 -178.310 -17.415 -178.030 ;
        RECT -17.235 -178.300 -16.955 -178.020 ;
        RECT -7.775 -178.310 -7.495 -178.030 ;
        RECT -7.315 -178.300 -7.035 -178.020 ;
        RECT 2.145 -178.310 2.425 -178.030 ;
        RECT 2.605 -178.300 2.885 -178.020 ;
        RECT 12.065 -178.310 12.345 -178.030 ;
        RECT 12.525 -178.300 12.805 -178.020 ;
        RECT 21.985 -178.310 22.265 -178.030 ;
        RECT 22.445 -178.300 22.725 -178.020 ;
        RECT -277.885 -179.070 -277.605 -178.790 ;
        RECT -267.965 -179.070 -267.685 -178.790 ;
        RECT -258.045 -179.070 -257.765 -178.790 ;
        RECT -248.125 -179.070 -247.845 -178.790 ;
        RECT -238.205 -179.070 -237.925 -178.790 ;
        RECT -228.285 -179.070 -228.005 -178.790 ;
        RECT -218.365 -179.070 -218.085 -178.790 ;
        RECT -208.445 -179.070 -208.165 -178.790 ;
        RECT -198.525 -179.070 -198.245 -178.790 ;
        RECT -188.605 -179.070 -188.325 -178.790 ;
        RECT -178.685 -179.070 -178.405 -178.790 ;
        RECT -168.765 -179.070 -168.485 -178.790 ;
        RECT -158.845 -179.070 -158.565 -178.790 ;
        RECT -148.925 -179.070 -148.645 -178.790 ;
        RECT -139.005 -179.070 -138.725 -178.790 ;
        RECT -129.085 -179.070 -128.805 -178.790 ;
        RECT -119.165 -179.070 -118.885 -178.790 ;
        RECT -109.245 -179.070 -108.965 -178.790 ;
        RECT -99.325 -179.070 -99.045 -178.790 ;
        RECT -89.405 -179.070 -89.125 -178.790 ;
        RECT -79.485 -179.070 -79.205 -178.790 ;
        RECT -69.565 -179.070 -69.285 -178.790 ;
        RECT -59.645 -179.070 -59.365 -178.790 ;
        RECT -49.725 -179.070 -49.445 -178.790 ;
        RECT -39.805 -179.070 -39.525 -178.790 ;
        RECT -29.885 -179.070 -29.605 -178.790 ;
        RECT -19.965 -179.070 -19.685 -178.790 ;
        RECT -10.045 -179.070 -9.765 -178.790 ;
        RECT -0.125 -179.070 0.155 -178.790 ;
        RECT 9.795 -179.070 10.075 -178.790 ;
        RECT 19.715 -179.070 19.995 -178.790 ;
      LAYER met3 ;
        RECT -288.280 93.760 -287.110 94.560 ;
        RECT -278.360 93.760 -277.190 94.560 ;
        RECT -268.440 93.760 -267.270 94.560 ;
        RECT -258.520 93.760 -257.350 94.560 ;
        RECT -248.600 93.760 -247.430 94.560 ;
        RECT -238.680 93.760 -237.510 94.560 ;
        RECT -228.760 93.760 -227.590 94.560 ;
        RECT -218.840 93.760 -217.670 94.560 ;
        RECT -208.920 93.760 -207.750 94.560 ;
        RECT -199.000 93.760 -197.830 94.560 ;
        RECT -189.080 93.760 -187.910 94.560 ;
        RECT -179.160 93.760 -177.990 94.560 ;
        RECT -169.240 93.760 -168.070 94.560 ;
        RECT -159.320 93.760 -158.150 94.560 ;
        RECT -149.400 93.760 -148.230 94.560 ;
        RECT -139.480 93.760 -138.310 94.560 ;
        RECT -129.560 93.760 -128.390 94.560 ;
        RECT -119.640 93.760 -118.470 94.560 ;
        RECT -109.720 93.760 -108.550 94.560 ;
        RECT -99.800 93.760 -98.630 94.560 ;
        RECT -89.880 93.760 -88.710 94.560 ;
        RECT -79.960 93.760 -78.790 94.560 ;
        RECT -70.040 93.760 -68.870 94.560 ;
        RECT -60.120 93.760 -58.950 94.560 ;
        RECT -50.200 93.760 -49.030 94.560 ;
        RECT -40.280 93.760 -39.110 94.560 ;
        RECT -30.360 93.760 -29.190 94.560 ;
        RECT -20.440 93.760 -19.270 94.560 ;
        RECT -10.520 93.760 -9.350 94.560 ;
        RECT -0.600 93.760 0.570 94.560 ;
        RECT 9.320 93.760 10.490 94.560 ;
        RECT 19.240 93.760 20.410 94.560 ;
        RECT -280.620 93.090 -279.700 93.570 ;
        RECT -270.700 93.090 -269.780 93.570 ;
        RECT -260.740 93.090 -259.860 93.570 ;
        RECT -250.860 93.090 -249.940 93.570 ;
        RECT -240.940 93.090 -240.020 93.570 ;
        RECT -231.020 93.090 -230.100 93.570 ;
        RECT -221.100 93.090 -220.180 93.570 ;
        RECT -211.160 93.090 -210.260 93.570 ;
        RECT -201.260 93.090 -200.340 93.570 ;
        RECT -191.340 93.090 -190.420 93.570 ;
        RECT -181.420 93.090 -180.500 93.570 ;
        RECT -171.480 93.090 -170.580 93.570 ;
        RECT -161.550 93.090 -160.660 93.570 ;
        RECT -151.660 93.090 -150.740 93.570 ;
        RECT -141.740 93.090 -140.820 93.570 ;
        RECT -131.820 93.090 -130.900 93.570 ;
        RECT -121.880 93.090 -120.980 93.570 ;
        RECT -111.980 93.090 -111.060 93.570 ;
        RECT -102.060 93.090 -101.140 93.570 ;
        RECT -92.140 93.090 -91.220 93.570 ;
        RECT -82.200 93.090 -81.300 93.570 ;
        RECT -72.300 93.090 -71.380 93.570 ;
        RECT -62.360 93.090 -61.460 93.570 ;
        RECT -52.450 93.090 -51.540 93.570 ;
        RECT -42.540 93.090 -41.620 93.570 ;
        RECT -32.620 93.090 -31.700 93.570 ;
        RECT -22.700 93.090 -21.780 93.570 ;
        RECT -12.780 93.090 -11.860 93.570 ;
        RECT -2.860 93.090 -1.940 93.570 ;
        RECT 7.060 93.090 7.980 93.570 ;
        RECT 16.980 93.090 17.900 93.570 ;
        RECT -287.880 90.370 -286.960 90.850 ;
        RECT -277.960 90.370 -277.060 90.850 ;
        RECT -268.040 90.370 -267.120 90.850 ;
        RECT -258.120 90.370 -257.220 90.850 ;
        RECT -248.200 90.370 -247.290 90.850 ;
        RECT -238.280 90.370 -237.380 90.850 ;
        RECT -228.360 90.370 -227.450 90.850 ;
        RECT -218.440 90.370 -217.520 90.850 ;
        RECT -208.520 90.370 -207.600 90.850 ;
        RECT -198.600 90.370 -197.720 90.850 ;
        RECT -188.680 90.370 -187.760 90.850 ;
        RECT -178.760 90.370 -177.850 90.850 ;
        RECT -168.840 90.370 -167.920 90.850 ;
        RECT -158.920 90.370 -158.010 90.850 ;
        RECT -149.000 90.370 -148.090 90.850 ;
        RECT -139.080 90.370 -138.160 90.850 ;
        RECT -129.160 90.370 -128.240 90.850 ;
        RECT -119.240 90.370 -118.340 90.850 ;
        RECT -109.320 90.370 -108.420 90.850 ;
        RECT -99.400 90.370 -98.480 90.850 ;
        RECT -89.480 90.370 -88.560 90.850 ;
        RECT -79.560 90.370 -78.650 90.850 ;
        RECT -69.640 90.370 -68.720 90.850 ;
        RECT -59.720 90.370 -58.820 90.850 ;
        RECT -49.800 90.370 -48.880 90.850 ;
        RECT -39.880 90.370 -38.980 90.850 ;
        RECT -29.960 90.370 -29.050 90.850 ;
        RECT -20.040 90.370 -19.120 90.850 ;
        RECT -10.120 90.370 -9.220 90.850 ;
        RECT -0.200 90.370 0.700 90.850 ;
        RECT 9.720 90.370 10.640 90.850 ;
        RECT 19.640 90.370 20.560 90.850 ;
        RECT -280.460 89.390 -279.290 90.190 ;
        RECT -270.540 89.390 -269.370 90.190 ;
        RECT -260.620 89.390 -259.450 90.190 ;
        RECT -250.700 89.390 -249.530 90.190 ;
        RECT -240.780 89.390 -239.610 90.190 ;
        RECT -230.860 89.390 -229.690 90.190 ;
        RECT -220.940 89.390 -219.770 90.190 ;
        RECT -211.020 89.390 -209.850 90.190 ;
        RECT -201.100 89.390 -199.930 90.190 ;
        RECT -191.180 89.390 -190.010 90.190 ;
        RECT -181.260 89.390 -180.090 90.190 ;
        RECT -171.340 89.390 -170.170 90.190 ;
        RECT -161.420 89.390 -160.250 90.190 ;
        RECT -151.500 89.390 -150.330 90.190 ;
        RECT -141.580 89.390 -140.410 90.190 ;
        RECT -131.660 89.390 -130.490 90.190 ;
        RECT -121.740 89.390 -120.570 90.190 ;
        RECT -111.820 89.390 -110.650 90.190 ;
        RECT -101.900 89.390 -100.730 90.190 ;
        RECT -91.980 89.390 -90.810 90.190 ;
        RECT -82.060 89.390 -80.890 90.190 ;
        RECT -72.140 89.390 -70.970 90.190 ;
        RECT -62.220 89.390 -61.050 90.190 ;
        RECT -52.300 89.390 -51.130 90.190 ;
        RECT -42.380 89.390 -41.210 90.190 ;
        RECT -32.460 89.390 -31.290 90.190 ;
        RECT -22.540 89.390 -21.370 90.190 ;
        RECT -12.620 89.390 -11.450 90.190 ;
        RECT -2.700 89.390 -1.530 90.190 ;
        RECT 7.220 89.390 8.390 90.190 ;
        RECT 17.140 89.390 18.310 90.190 ;
        RECT -288.030 6.050 -286.860 6.850 ;
        RECT -278.110 6.050 -276.940 6.850 ;
        RECT -268.190 6.050 -267.020 6.850 ;
        RECT -258.270 6.050 -257.100 6.850 ;
        RECT -248.350 6.050 -247.180 6.850 ;
        RECT -238.430 6.050 -237.260 6.850 ;
        RECT -228.510 6.050 -227.340 6.850 ;
        RECT -218.590 6.050 -217.420 6.850 ;
        RECT -208.670 6.050 -207.500 6.850 ;
        RECT -198.750 6.050 -197.580 6.850 ;
        RECT -188.830 6.050 -187.660 6.850 ;
        RECT -178.910 6.050 -177.740 6.850 ;
        RECT -168.990 6.050 -167.820 6.850 ;
        RECT -159.070 6.050 -157.900 6.850 ;
        RECT -149.150 6.050 -147.980 6.850 ;
        RECT -139.230 6.050 -138.060 6.850 ;
        RECT -129.310 6.050 -128.140 6.850 ;
        RECT -119.390 6.050 -118.220 6.850 ;
        RECT -109.470 6.050 -108.300 6.850 ;
        RECT -99.550 6.050 -98.380 6.850 ;
        RECT -89.630 6.050 -88.460 6.850 ;
        RECT -79.710 6.050 -78.540 6.850 ;
        RECT -69.790 6.050 -68.620 6.850 ;
        RECT -59.870 6.050 -58.700 6.850 ;
        RECT -49.950 6.050 -48.780 6.850 ;
        RECT -40.030 6.050 -38.860 6.850 ;
        RECT -30.110 6.050 -28.940 6.850 ;
        RECT -20.190 6.050 -19.020 6.850 ;
        RECT -10.270 6.050 -9.100 6.850 ;
        RECT -0.350 6.050 0.820 6.850 ;
        RECT 9.570 6.050 10.740 6.850 ;
        RECT 19.490 6.050 20.660 6.850 ;
        RECT -280.370 5.380 -279.450 5.860 ;
        RECT -270.450 5.380 -269.530 5.860 ;
        RECT -260.490 5.380 -259.610 5.860 ;
        RECT -250.610 5.380 -249.690 5.860 ;
        RECT -240.690 5.380 -239.770 5.860 ;
        RECT -230.770 5.380 -229.850 5.860 ;
        RECT -220.850 5.380 -219.930 5.860 ;
        RECT -210.910 5.380 -210.010 5.860 ;
        RECT -201.010 5.380 -200.090 5.860 ;
        RECT -191.090 5.380 -190.170 5.860 ;
        RECT -181.170 5.380 -180.250 5.860 ;
        RECT -171.230 5.380 -170.330 5.860 ;
        RECT -161.300 5.380 -160.410 5.860 ;
        RECT -151.410 5.380 -150.490 5.860 ;
        RECT -141.490 5.380 -140.570 5.860 ;
        RECT -131.570 5.380 -130.650 5.860 ;
        RECT -121.630 5.380 -120.730 5.860 ;
        RECT -111.730 5.380 -110.810 5.860 ;
        RECT -101.810 5.380 -100.890 5.860 ;
        RECT -91.890 5.380 -90.970 5.860 ;
        RECT -81.950 5.380 -81.050 5.860 ;
        RECT -72.050 5.380 -71.130 5.860 ;
        RECT -62.110 5.380 -61.210 5.860 ;
        RECT -52.200 5.380 -51.290 5.860 ;
        RECT -42.290 5.380 -41.370 5.860 ;
        RECT -32.370 5.380 -31.450 5.860 ;
        RECT -22.450 5.380 -21.530 5.860 ;
        RECT -12.530 5.380 -11.610 5.860 ;
        RECT -2.610 5.380 -1.690 5.860 ;
        RECT 7.310 5.380 8.230 5.860 ;
        RECT 17.230 5.380 18.150 5.860 ;
        RECT -287.630 2.660 -286.710 3.140 ;
        RECT -277.710 2.660 -276.810 3.140 ;
        RECT -267.790 2.660 -266.870 3.140 ;
        RECT -257.870 2.660 -256.970 3.140 ;
        RECT -247.950 2.660 -247.040 3.140 ;
        RECT -238.030 2.660 -237.130 3.140 ;
        RECT -228.110 2.660 -227.200 3.140 ;
        RECT -218.190 2.660 -217.270 3.140 ;
        RECT -208.270 2.660 -207.350 3.140 ;
        RECT -198.350 2.660 -197.470 3.140 ;
        RECT -188.430 2.660 -187.510 3.140 ;
        RECT -178.510 2.660 -177.600 3.140 ;
        RECT -168.590 2.660 -167.670 3.140 ;
        RECT -158.670 2.660 -157.760 3.140 ;
        RECT -148.750 2.660 -147.840 3.140 ;
        RECT -138.830 2.660 -137.910 3.140 ;
        RECT -128.910 2.660 -127.990 3.140 ;
        RECT -118.990 2.660 -118.090 3.140 ;
        RECT -109.070 2.660 -108.170 3.140 ;
        RECT -99.150 2.660 -98.230 3.140 ;
        RECT -89.230 2.660 -88.310 3.140 ;
        RECT -79.310 2.660 -78.400 3.140 ;
        RECT -69.390 2.660 -68.470 3.140 ;
        RECT -59.470 2.660 -58.570 3.140 ;
        RECT -49.550 2.660 -48.630 3.140 ;
        RECT -39.630 2.660 -38.730 3.140 ;
        RECT -29.710 2.660 -28.800 3.140 ;
        RECT -19.790 2.660 -18.870 3.140 ;
        RECT -9.870 2.660 -8.970 3.140 ;
        RECT 0.050 2.660 0.950 3.140 ;
        RECT 9.970 2.660 10.890 3.140 ;
        RECT 19.890 2.660 20.810 3.140 ;
        RECT -280.210 1.680 -279.040 2.480 ;
        RECT -270.290 1.680 -269.120 2.480 ;
        RECT -260.370 1.680 -259.200 2.480 ;
        RECT -250.450 1.680 -249.280 2.480 ;
        RECT -240.530 1.680 -239.360 2.480 ;
        RECT -230.610 1.680 -229.440 2.480 ;
        RECT -220.690 1.680 -219.520 2.480 ;
        RECT -210.770 1.680 -209.600 2.480 ;
        RECT -200.850 1.680 -199.680 2.480 ;
        RECT -190.930 1.680 -189.760 2.480 ;
        RECT -181.010 1.680 -179.840 2.480 ;
        RECT -171.090 1.680 -169.920 2.480 ;
        RECT -161.170 1.680 -160.000 2.480 ;
        RECT -151.250 1.680 -150.080 2.480 ;
        RECT -141.330 1.680 -140.160 2.480 ;
        RECT -131.410 1.680 -130.240 2.480 ;
        RECT -121.490 1.680 -120.320 2.480 ;
        RECT -111.570 1.680 -110.400 2.480 ;
        RECT -101.650 1.680 -100.480 2.480 ;
        RECT -91.730 1.680 -90.560 2.480 ;
        RECT -81.810 1.680 -80.640 2.480 ;
        RECT -71.890 1.680 -70.720 2.480 ;
        RECT -61.970 1.680 -60.800 2.480 ;
        RECT -52.050 1.680 -50.880 2.480 ;
        RECT -42.130 1.680 -40.960 2.480 ;
        RECT -32.210 1.680 -31.040 2.480 ;
        RECT -22.290 1.680 -21.120 2.480 ;
        RECT -12.370 1.680 -11.200 2.480 ;
        RECT -2.450 1.680 -1.280 2.480 ;
        RECT 7.470 1.680 8.640 2.480 ;
        RECT 17.390 1.680 18.560 2.480 ;
        RECT -286.270 -87.300 -285.100 -86.500 ;
        RECT -276.350 -87.300 -275.180 -86.500 ;
        RECT -266.430 -87.300 -265.260 -86.500 ;
        RECT -256.510 -87.300 -255.340 -86.500 ;
        RECT -246.590 -87.300 -245.420 -86.500 ;
        RECT -236.670 -87.300 -235.500 -86.500 ;
        RECT -226.750 -87.300 -225.580 -86.500 ;
        RECT -216.830 -87.300 -215.660 -86.500 ;
        RECT -206.910 -87.300 -205.740 -86.500 ;
        RECT -196.990 -87.300 -195.820 -86.500 ;
        RECT -187.070 -87.300 -185.900 -86.500 ;
        RECT -177.150 -87.300 -175.980 -86.500 ;
        RECT -167.230 -87.300 -166.060 -86.500 ;
        RECT -157.310 -87.300 -156.140 -86.500 ;
        RECT -147.390 -87.300 -146.220 -86.500 ;
        RECT -137.470 -87.300 -136.300 -86.500 ;
        RECT -127.550 -87.300 -126.380 -86.500 ;
        RECT -117.630 -87.300 -116.460 -86.500 ;
        RECT -107.710 -87.300 -106.540 -86.500 ;
        RECT -97.790 -87.300 -96.620 -86.500 ;
        RECT -87.870 -87.300 -86.700 -86.500 ;
        RECT -77.950 -87.300 -76.780 -86.500 ;
        RECT -68.030 -87.300 -66.860 -86.500 ;
        RECT -58.110 -87.300 -56.940 -86.500 ;
        RECT -48.190 -87.300 -47.020 -86.500 ;
        RECT -38.270 -87.300 -37.100 -86.500 ;
        RECT -28.350 -87.300 -27.180 -86.500 ;
        RECT -18.430 -87.300 -17.260 -86.500 ;
        RECT -8.510 -87.300 -7.340 -86.500 ;
        RECT 1.410 -87.300 2.580 -86.500 ;
        RECT 11.330 -87.300 12.500 -86.500 ;
        RECT 21.250 -87.300 22.420 -86.500 ;
        RECT -278.610 -87.970 -277.690 -87.490 ;
        RECT -268.690 -87.970 -267.770 -87.490 ;
        RECT -258.730 -87.970 -257.850 -87.490 ;
        RECT -248.850 -87.970 -247.930 -87.490 ;
        RECT -238.930 -87.970 -238.010 -87.490 ;
        RECT -229.010 -87.970 -228.090 -87.490 ;
        RECT -219.090 -87.970 -218.170 -87.490 ;
        RECT -209.150 -87.970 -208.250 -87.490 ;
        RECT -199.250 -87.970 -198.330 -87.490 ;
        RECT -189.330 -87.970 -188.410 -87.490 ;
        RECT -179.410 -87.970 -178.490 -87.490 ;
        RECT -169.470 -87.970 -168.570 -87.490 ;
        RECT -159.540 -87.970 -158.650 -87.490 ;
        RECT -149.650 -87.970 -148.730 -87.490 ;
        RECT -139.730 -87.970 -138.810 -87.490 ;
        RECT -129.810 -87.970 -128.890 -87.490 ;
        RECT -119.870 -87.970 -118.970 -87.490 ;
        RECT -109.970 -87.970 -109.050 -87.490 ;
        RECT -100.050 -87.970 -99.130 -87.490 ;
        RECT -90.130 -87.970 -89.210 -87.490 ;
        RECT -80.190 -87.970 -79.290 -87.490 ;
        RECT -70.290 -87.970 -69.370 -87.490 ;
        RECT -60.350 -87.970 -59.450 -87.490 ;
        RECT -50.440 -87.970 -49.530 -87.490 ;
        RECT -40.530 -87.970 -39.610 -87.490 ;
        RECT -30.610 -87.970 -29.690 -87.490 ;
        RECT -20.690 -87.970 -19.770 -87.490 ;
        RECT -10.770 -87.970 -9.850 -87.490 ;
        RECT -0.850 -87.970 0.070 -87.490 ;
        RECT 9.070 -87.970 9.990 -87.490 ;
        RECT 18.990 -87.970 19.910 -87.490 ;
        RECT -285.870 -90.690 -284.950 -90.210 ;
        RECT -275.950 -90.690 -275.050 -90.210 ;
        RECT -266.030 -90.690 -265.110 -90.210 ;
        RECT -256.110 -90.690 -255.210 -90.210 ;
        RECT -246.190 -90.690 -245.280 -90.210 ;
        RECT -236.270 -90.690 -235.370 -90.210 ;
        RECT -226.350 -90.690 -225.440 -90.210 ;
        RECT -216.430 -90.690 -215.510 -90.210 ;
        RECT -206.510 -90.690 -205.590 -90.210 ;
        RECT -196.590 -90.690 -195.710 -90.210 ;
        RECT -186.670 -90.690 -185.750 -90.210 ;
        RECT -176.750 -90.690 -175.840 -90.210 ;
        RECT -166.830 -90.690 -165.910 -90.210 ;
        RECT -156.910 -90.690 -156.000 -90.210 ;
        RECT -146.990 -90.690 -146.080 -90.210 ;
        RECT -137.070 -90.690 -136.150 -90.210 ;
        RECT -127.150 -90.690 -126.230 -90.210 ;
        RECT -117.230 -90.690 -116.330 -90.210 ;
        RECT -107.310 -90.690 -106.410 -90.210 ;
        RECT -97.390 -90.690 -96.470 -90.210 ;
        RECT -87.470 -90.690 -86.550 -90.210 ;
        RECT -77.550 -90.690 -76.640 -90.210 ;
        RECT -67.630 -90.690 -66.710 -90.210 ;
        RECT -57.710 -90.690 -56.810 -90.210 ;
        RECT -47.790 -90.690 -46.870 -90.210 ;
        RECT -37.870 -90.690 -36.970 -90.210 ;
        RECT -27.950 -90.690 -27.040 -90.210 ;
        RECT -18.030 -90.690 -17.110 -90.210 ;
        RECT -8.110 -90.690 -7.210 -90.210 ;
        RECT 1.810 -90.690 2.710 -90.210 ;
        RECT 11.730 -90.690 12.650 -90.210 ;
        RECT 21.650 -90.690 22.570 -90.210 ;
        RECT -278.450 -91.670 -277.280 -90.870 ;
        RECT -268.530 -91.670 -267.360 -90.870 ;
        RECT -258.610 -91.670 -257.440 -90.870 ;
        RECT -248.690 -91.670 -247.520 -90.870 ;
        RECT -238.770 -91.670 -237.600 -90.870 ;
        RECT -228.850 -91.670 -227.680 -90.870 ;
        RECT -218.930 -91.670 -217.760 -90.870 ;
        RECT -209.010 -91.670 -207.840 -90.870 ;
        RECT -199.090 -91.670 -197.920 -90.870 ;
        RECT -189.170 -91.670 -188.000 -90.870 ;
        RECT -179.250 -91.670 -178.080 -90.870 ;
        RECT -169.330 -91.670 -168.160 -90.870 ;
        RECT -159.410 -91.670 -158.240 -90.870 ;
        RECT -149.490 -91.670 -148.320 -90.870 ;
        RECT -139.570 -91.670 -138.400 -90.870 ;
        RECT -129.650 -91.670 -128.480 -90.870 ;
        RECT -119.730 -91.670 -118.560 -90.870 ;
        RECT -109.810 -91.670 -108.640 -90.870 ;
        RECT -99.890 -91.670 -98.720 -90.870 ;
        RECT -89.970 -91.670 -88.800 -90.870 ;
        RECT -80.050 -91.670 -78.880 -90.870 ;
        RECT -70.130 -91.670 -68.960 -90.870 ;
        RECT -60.210 -91.670 -59.040 -90.870 ;
        RECT -50.290 -91.670 -49.120 -90.870 ;
        RECT -40.370 -91.670 -39.200 -90.870 ;
        RECT -30.450 -91.670 -29.280 -90.870 ;
        RECT -20.530 -91.670 -19.360 -90.870 ;
        RECT -10.610 -91.670 -9.440 -90.870 ;
        RECT -0.690 -91.670 0.480 -90.870 ;
        RECT 9.230 -91.670 10.400 -90.870 ;
        RECT 19.150 -91.670 20.320 -90.870 ;
        RECT -286.020 -175.010 -284.850 -174.210 ;
        RECT -276.100 -175.010 -274.930 -174.210 ;
        RECT -266.180 -175.010 -265.010 -174.210 ;
        RECT -256.260 -175.010 -255.090 -174.210 ;
        RECT -246.340 -175.010 -245.170 -174.210 ;
        RECT -236.420 -175.010 -235.250 -174.210 ;
        RECT -226.500 -175.010 -225.330 -174.210 ;
        RECT -216.580 -175.010 -215.410 -174.210 ;
        RECT -206.660 -175.010 -205.490 -174.210 ;
        RECT -196.740 -175.010 -195.570 -174.210 ;
        RECT -186.820 -175.010 -185.650 -174.210 ;
        RECT -176.900 -175.010 -175.730 -174.210 ;
        RECT -166.980 -175.010 -165.810 -174.210 ;
        RECT -157.060 -175.010 -155.890 -174.210 ;
        RECT -147.140 -175.010 -145.970 -174.210 ;
        RECT -137.220 -175.010 -136.050 -174.210 ;
        RECT -127.300 -175.010 -126.130 -174.210 ;
        RECT -117.380 -175.010 -116.210 -174.210 ;
        RECT -107.460 -175.010 -106.290 -174.210 ;
        RECT -97.540 -175.010 -96.370 -174.210 ;
        RECT -87.620 -175.010 -86.450 -174.210 ;
        RECT -77.700 -175.010 -76.530 -174.210 ;
        RECT -67.780 -175.010 -66.610 -174.210 ;
        RECT -57.860 -175.010 -56.690 -174.210 ;
        RECT -47.940 -175.010 -46.770 -174.210 ;
        RECT -38.020 -175.010 -36.850 -174.210 ;
        RECT -28.100 -175.010 -26.930 -174.210 ;
        RECT -18.180 -175.010 -17.010 -174.210 ;
        RECT -8.260 -175.010 -7.090 -174.210 ;
        RECT 1.660 -175.010 2.830 -174.210 ;
        RECT 11.580 -175.010 12.750 -174.210 ;
        RECT 21.500 -175.010 22.670 -174.210 ;
        RECT -278.360 -175.680 -277.440 -175.200 ;
        RECT -268.440 -175.680 -267.520 -175.200 ;
        RECT -258.480 -175.680 -257.600 -175.200 ;
        RECT -248.600 -175.680 -247.680 -175.200 ;
        RECT -238.680 -175.680 -237.760 -175.200 ;
        RECT -228.760 -175.680 -227.840 -175.200 ;
        RECT -218.840 -175.680 -217.920 -175.200 ;
        RECT -208.900 -175.680 -208.000 -175.200 ;
        RECT -199.000 -175.680 -198.080 -175.200 ;
        RECT -189.080 -175.680 -188.160 -175.200 ;
        RECT -179.160 -175.680 -178.240 -175.200 ;
        RECT -169.220 -175.680 -168.320 -175.200 ;
        RECT -159.290 -175.680 -158.400 -175.200 ;
        RECT -149.400 -175.680 -148.480 -175.200 ;
        RECT -139.480 -175.680 -138.560 -175.200 ;
        RECT -129.560 -175.680 -128.640 -175.200 ;
        RECT -119.620 -175.680 -118.720 -175.200 ;
        RECT -109.720 -175.680 -108.800 -175.200 ;
        RECT -99.800 -175.680 -98.880 -175.200 ;
        RECT -89.880 -175.680 -88.960 -175.200 ;
        RECT -79.940 -175.680 -79.040 -175.200 ;
        RECT -70.040 -175.680 -69.120 -175.200 ;
        RECT -60.100 -175.680 -59.200 -175.200 ;
        RECT -50.190 -175.680 -49.280 -175.200 ;
        RECT -40.280 -175.680 -39.360 -175.200 ;
        RECT -30.360 -175.680 -29.440 -175.200 ;
        RECT -20.440 -175.680 -19.520 -175.200 ;
        RECT -10.520 -175.680 -9.600 -175.200 ;
        RECT -0.600 -175.680 0.320 -175.200 ;
        RECT 9.320 -175.680 10.240 -175.200 ;
        RECT 19.240 -175.680 20.160 -175.200 ;
        RECT -285.620 -178.400 -284.700 -177.920 ;
        RECT -275.700 -178.400 -274.800 -177.920 ;
        RECT -265.780 -178.400 -264.860 -177.920 ;
        RECT -255.860 -178.400 -254.960 -177.920 ;
        RECT -245.940 -178.400 -245.030 -177.920 ;
        RECT -236.020 -178.400 -235.120 -177.920 ;
        RECT -226.100 -178.400 -225.190 -177.920 ;
        RECT -216.180 -178.400 -215.260 -177.920 ;
        RECT -206.260 -178.400 -205.340 -177.920 ;
        RECT -196.340 -178.400 -195.460 -177.920 ;
        RECT -186.420 -178.400 -185.500 -177.920 ;
        RECT -176.500 -178.400 -175.590 -177.920 ;
        RECT -166.580 -178.400 -165.660 -177.920 ;
        RECT -156.660 -178.400 -155.750 -177.920 ;
        RECT -146.740 -178.400 -145.830 -177.920 ;
        RECT -136.820 -178.400 -135.900 -177.920 ;
        RECT -126.900 -178.400 -125.980 -177.920 ;
        RECT -116.980 -178.400 -116.080 -177.920 ;
        RECT -107.060 -178.400 -106.160 -177.920 ;
        RECT -97.140 -178.400 -96.220 -177.920 ;
        RECT -87.220 -178.400 -86.300 -177.920 ;
        RECT -77.300 -178.400 -76.390 -177.920 ;
        RECT -67.380 -178.400 -66.460 -177.920 ;
        RECT -57.460 -178.400 -56.560 -177.920 ;
        RECT -47.540 -178.400 -46.620 -177.920 ;
        RECT -37.620 -178.400 -36.720 -177.920 ;
        RECT -27.700 -178.400 -26.790 -177.920 ;
        RECT -17.780 -178.400 -16.860 -177.920 ;
        RECT -7.860 -178.400 -6.960 -177.920 ;
        RECT 2.060 -178.400 2.960 -177.920 ;
        RECT 11.980 -178.400 12.900 -177.920 ;
        RECT 21.900 -178.400 22.820 -177.920 ;
        RECT -278.200 -179.380 -277.030 -178.580 ;
        RECT -268.280 -179.380 -267.110 -178.580 ;
        RECT -258.360 -179.380 -257.190 -178.580 ;
        RECT -248.440 -179.380 -247.270 -178.580 ;
        RECT -238.520 -179.380 -237.350 -178.580 ;
        RECT -228.600 -179.380 -227.430 -178.580 ;
        RECT -218.680 -179.380 -217.510 -178.580 ;
        RECT -208.760 -179.380 -207.590 -178.580 ;
        RECT -198.840 -179.380 -197.670 -178.580 ;
        RECT -188.920 -179.380 -187.750 -178.580 ;
        RECT -179.000 -179.380 -177.830 -178.580 ;
        RECT -169.080 -179.380 -167.910 -178.580 ;
        RECT -159.160 -179.380 -157.990 -178.580 ;
        RECT -149.240 -179.380 -148.070 -178.580 ;
        RECT -139.320 -179.380 -138.150 -178.580 ;
        RECT -129.400 -179.380 -128.230 -178.580 ;
        RECT -119.480 -179.380 -118.310 -178.580 ;
        RECT -109.560 -179.380 -108.390 -178.580 ;
        RECT -99.640 -179.380 -98.470 -178.580 ;
        RECT -89.720 -179.380 -88.550 -178.580 ;
        RECT -79.800 -179.380 -78.630 -178.580 ;
        RECT -69.880 -179.380 -68.710 -178.580 ;
        RECT -59.960 -179.380 -58.790 -178.580 ;
        RECT -50.040 -179.380 -48.870 -178.580 ;
        RECT -40.120 -179.380 -38.950 -178.580 ;
        RECT -30.200 -179.380 -29.030 -178.580 ;
        RECT -20.280 -179.380 -19.110 -178.580 ;
        RECT -10.360 -179.380 -9.190 -178.580 ;
        RECT -0.440 -179.380 0.730 -178.580 ;
        RECT 9.480 -179.380 10.650 -178.580 ;
        RECT 19.400 -179.380 20.570 -178.580 ;
      LAYER via3 ;
        RECT -287.730 94.035 -287.410 94.355 ;
        RECT -277.810 94.035 -277.490 94.355 ;
        RECT -267.890 94.035 -267.570 94.355 ;
        RECT -257.970 94.035 -257.650 94.355 ;
        RECT -248.050 94.035 -247.730 94.355 ;
        RECT -238.130 94.035 -237.810 94.355 ;
        RECT -228.210 94.035 -227.890 94.355 ;
        RECT -218.290 94.035 -217.970 94.355 ;
        RECT -208.370 94.035 -208.050 94.355 ;
        RECT -198.450 94.035 -198.130 94.355 ;
        RECT -188.530 94.035 -188.210 94.355 ;
        RECT -178.610 94.035 -178.290 94.355 ;
        RECT -168.690 94.035 -168.370 94.355 ;
        RECT -158.770 94.035 -158.450 94.355 ;
        RECT -148.850 94.035 -148.530 94.355 ;
        RECT -138.930 94.035 -138.610 94.355 ;
        RECT -129.010 94.035 -128.690 94.355 ;
        RECT -119.090 94.035 -118.770 94.355 ;
        RECT -109.170 94.035 -108.850 94.355 ;
        RECT -99.250 94.035 -98.930 94.355 ;
        RECT -89.330 94.035 -89.010 94.355 ;
        RECT -79.410 94.035 -79.090 94.355 ;
        RECT -69.490 94.035 -69.170 94.355 ;
        RECT -59.570 94.035 -59.250 94.355 ;
        RECT -49.650 94.035 -49.330 94.355 ;
        RECT -39.730 94.035 -39.410 94.355 ;
        RECT -29.810 94.035 -29.490 94.355 ;
        RECT -19.890 94.035 -19.570 94.355 ;
        RECT -9.970 94.035 -9.650 94.355 ;
        RECT -0.050 94.035 0.270 94.355 ;
        RECT 9.870 94.035 10.190 94.355 ;
        RECT 19.790 94.035 20.110 94.355 ;
        RECT -280.550 93.165 -280.230 93.485 ;
        RECT -280.080 93.165 -279.760 93.485 ;
        RECT -270.630 93.165 -270.310 93.485 ;
        RECT -270.160 93.165 -269.840 93.485 ;
        RECT -260.710 93.165 -260.390 93.485 ;
        RECT -260.240 93.165 -259.920 93.485 ;
        RECT -250.790 93.165 -250.470 93.485 ;
        RECT -250.320 93.165 -250.000 93.485 ;
        RECT -240.870 93.165 -240.550 93.485 ;
        RECT -240.400 93.165 -240.080 93.485 ;
        RECT -230.950 93.165 -230.630 93.485 ;
        RECT -230.480 93.165 -230.160 93.485 ;
        RECT -221.030 93.165 -220.710 93.485 ;
        RECT -220.560 93.165 -220.240 93.485 ;
        RECT -211.110 93.165 -210.790 93.485 ;
        RECT -210.640 93.165 -210.320 93.485 ;
        RECT -201.190 93.165 -200.870 93.485 ;
        RECT -200.720 93.165 -200.400 93.485 ;
        RECT -191.270 93.165 -190.950 93.485 ;
        RECT -190.800 93.165 -190.480 93.485 ;
        RECT -181.350 93.165 -181.030 93.485 ;
        RECT -180.880 93.165 -180.560 93.485 ;
        RECT -171.430 93.165 -171.110 93.485 ;
        RECT -170.960 93.165 -170.640 93.485 ;
        RECT -161.510 93.165 -161.190 93.485 ;
        RECT -161.040 93.165 -160.720 93.485 ;
        RECT -151.590 93.165 -151.270 93.485 ;
        RECT -151.120 93.165 -150.800 93.485 ;
        RECT -141.670 93.165 -141.350 93.485 ;
        RECT -141.200 93.165 -140.880 93.485 ;
        RECT -131.750 93.165 -131.430 93.485 ;
        RECT -131.280 93.165 -130.960 93.485 ;
        RECT -121.830 93.165 -121.510 93.485 ;
        RECT -121.360 93.165 -121.040 93.485 ;
        RECT -111.910 93.165 -111.590 93.485 ;
        RECT -111.440 93.165 -111.120 93.485 ;
        RECT -101.990 93.165 -101.670 93.485 ;
        RECT -101.520 93.165 -101.200 93.485 ;
        RECT -92.070 93.165 -91.750 93.485 ;
        RECT -91.600 93.165 -91.280 93.485 ;
        RECT -82.150 93.165 -81.830 93.485 ;
        RECT -81.680 93.165 -81.360 93.485 ;
        RECT -72.230 93.165 -71.910 93.485 ;
        RECT -71.760 93.165 -71.440 93.485 ;
        RECT -62.310 93.165 -61.990 93.485 ;
        RECT -61.840 93.165 -61.520 93.485 ;
        RECT -52.390 93.165 -52.070 93.485 ;
        RECT -51.920 93.165 -51.600 93.485 ;
        RECT -42.470 93.165 -42.150 93.485 ;
        RECT -42.000 93.165 -41.680 93.485 ;
        RECT -32.550 93.165 -32.230 93.485 ;
        RECT -32.080 93.165 -31.760 93.485 ;
        RECT -22.630 93.165 -22.310 93.485 ;
        RECT -22.160 93.165 -21.840 93.485 ;
        RECT -12.710 93.165 -12.390 93.485 ;
        RECT -12.240 93.165 -11.920 93.485 ;
        RECT -2.790 93.165 -2.470 93.485 ;
        RECT -2.320 93.165 -2.000 93.485 ;
        RECT 7.130 93.165 7.450 93.485 ;
        RECT 7.600 93.165 7.920 93.485 ;
        RECT 17.050 93.165 17.370 93.485 ;
        RECT 17.520 93.165 17.840 93.485 ;
        RECT -287.810 90.445 -287.490 90.765 ;
        RECT -287.350 90.445 -287.030 90.765 ;
        RECT -277.890 90.445 -277.570 90.765 ;
        RECT -277.430 90.445 -277.110 90.765 ;
        RECT -267.970 90.445 -267.650 90.765 ;
        RECT -267.510 90.445 -267.190 90.765 ;
        RECT -258.050 90.445 -257.730 90.765 ;
        RECT -257.590 90.445 -257.270 90.765 ;
        RECT -248.130 90.445 -247.810 90.765 ;
        RECT -247.670 90.445 -247.350 90.765 ;
        RECT -238.210 90.445 -237.890 90.765 ;
        RECT -237.750 90.445 -237.430 90.765 ;
        RECT -228.290 90.445 -227.970 90.765 ;
        RECT -227.830 90.445 -227.510 90.765 ;
        RECT -218.370 90.445 -218.050 90.765 ;
        RECT -217.910 90.445 -217.590 90.765 ;
        RECT -208.450 90.445 -208.130 90.765 ;
        RECT -207.990 90.445 -207.670 90.765 ;
        RECT -198.530 90.445 -198.210 90.765 ;
        RECT -198.070 90.445 -197.750 90.765 ;
        RECT -188.610 90.445 -188.290 90.765 ;
        RECT -188.150 90.445 -187.830 90.765 ;
        RECT -178.690 90.445 -178.370 90.765 ;
        RECT -178.230 90.445 -177.910 90.765 ;
        RECT -168.770 90.445 -168.450 90.765 ;
        RECT -168.310 90.445 -167.990 90.765 ;
        RECT -158.850 90.445 -158.530 90.765 ;
        RECT -158.390 90.445 -158.070 90.765 ;
        RECT -148.930 90.445 -148.610 90.765 ;
        RECT -148.470 90.445 -148.150 90.765 ;
        RECT -139.010 90.445 -138.690 90.765 ;
        RECT -138.550 90.445 -138.230 90.765 ;
        RECT -129.090 90.445 -128.770 90.765 ;
        RECT -128.630 90.445 -128.310 90.765 ;
        RECT -119.170 90.445 -118.850 90.765 ;
        RECT -118.710 90.445 -118.390 90.765 ;
        RECT -109.250 90.445 -108.930 90.765 ;
        RECT -108.790 90.445 -108.470 90.765 ;
        RECT -99.330 90.445 -99.010 90.765 ;
        RECT -98.870 90.445 -98.550 90.765 ;
        RECT -89.410 90.445 -89.090 90.765 ;
        RECT -88.950 90.445 -88.630 90.765 ;
        RECT -79.490 90.445 -79.170 90.765 ;
        RECT -79.030 90.445 -78.710 90.765 ;
        RECT -69.570 90.445 -69.250 90.765 ;
        RECT -69.110 90.445 -68.790 90.765 ;
        RECT -59.650 90.445 -59.330 90.765 ;
        RECT -59.190 90.445 -58.870 90.765 ;
        RECT -49.730 90.445 -49.410 90.765 ;
        RECT -49.270 90.445 -48.950 90.765 ;
        RECT -39.810 90.445 -39.490 90.765 ;
        RECT -39.350 90.445 -39.030 90.765 ;
        RECT -29.890 90.445 -29.570 90.765 ;
        RECT -29.430 90.445 -29.110 90.765 ;
        RECT -19.970 90.445 -19.650 90.765 ;
        RECT -19.510 90.445 -19.190 90.765 ;
        RECT -10.050 90.445 -9.730 90.765 ;
        RECT -9.590 90.445 -9.270 90.765 ;
        RECT -0.130 90.445 0.190 90.765 ;
        RECT 0.330 90.445 0.650 90.765 ;
        RECT 9.790 90.445 10.110 90.765 ;
        RECT 10.250 90.445 10.570 90.765 ;
        RECT 19.710 90.445 20.030 90.765 ;
        RECT 20.170 90.445 20.490 90.765 ;
        RECT -280.160 89.685 -279.840 90.005 ;
        RECT -270.240 89.685 -269.920 90.005 ;
        RECT -260.320 89.685 -260.000 90.005 ;
        RECT -250.400 89.685 -250.080 90.005 ;
        RECT -240.480 89.685 -240.160 90.005 ;
        RECT -230.560 89.685 -230.240 90.005 ;
        RECT -220.640 89.685 -220.320 90.005 ;
        RECT -210.720 89.685 -210.400 90.005 ;
        RECT -200.800 89.685 -200.480 90.005 ;
        RECT -190.880 89.685 -190.560 90.005 ;
        RECT -180.960 89.685 -180.640 90.005 ;
        RECT -171.040 89.685 -170.720 90.005 ;
        RECT -161.120 89.685 -160.800 90.005 ;
        RECT -151.200 89.685 -150.880 90.005 ;
        RECT -141.280 89.685 -140.960 90.005 ;
        RECT -131.360 89.685 -131.040 90.005 ;
        RECT -121.440 89.685 -121.120 90.005 ;
        RECT -111.520 89.685 -111.200 90.005 ;
        RECT -101.600 89.685 -101.280 90.005 ;
        RECT -91.680 89.685 -91.360 90.005 ;
        RECT -81.760 89.685 -81.440 90.005 ;
        RECT -71.840 89.685 -71.520 90.005 ;
        RECT -61.920 89.685 -61.600 90.005 ;
        RECT -52.000 89.685 -51.680 90.005 ;
        RECT -42.080 89.685 -41.760 90.005 ;
        RECT -32.160 89.685 -31.840 90.005 ;
        RECT -22.240 89.685 -21.920 90.005 ;
        RECT -12.320 89.685 -12.000 90.005 ;
        RECT -2.400 89.685 -2.080 90.005 ;
        RECT 7.520 89.685 7.840 90.005 ;
        RECT 17.440 89.685 17.760 90.005 ;
        RECT -287.480 6.325 -287.160 6.645 ;
        RECT -277.560 6.325 -277.240 6.645 ;
        RECT -267.640 6.325 -267.320 6.645 ;
        RECT -257.720 6.325 -257.400 6.645 ;
        RECT -247.800 6.325 -247.480 6.645 ;
        RECT -237.880 6.325 -237.560 6.645 ;
        RECT -227.960 6.325 -227.640 6.645 ;
        RECT -218.040 6.325 -217.720 6.645 ;
        RECT -208.120 6.325 -207.800 6.645 ;
        RECT -198.200 6.325 -197.880 6.645 ;
        RECT -188.280 6.325 -187.960 6.645 ;
        RECT -178.360 6.325 -178.040 6.645 ;
        RECT -168.440 6.325 -168.120 6.645 ;
        RECT -158.520 6.325 -158.200 6.645 ;
        RECT -148.600 6.325 -148.280 6.645 ;
        RECT -138.680 6.325 -138.360 6.645 ;
        RECT -128.760 6.325 -128.440 6.645 ;
        RECT -118.840 6.325 -118.520 6.645 ;
        RECT -108.920 6.325 -108.600 6.645 ;
        RECT -99.000 6.325 -98.680 6.645 ;
        RECT -89.080 6.325 -88.760 6.645 ;
        RECT -79.160 6.325 -78.840 6.645 ;
        RECT -69.240 6.325 -68.920 6.645 ;
        RECT -59.320 6.325 -59.000 6.645 ;
        RECT -49.400 6.325 -49.080 6.645 ;
        RECT -39.480 6.325 -39.160 6.645 ;
        RECT -29.560 6.325 -29.240 6.645 ;
        RECT -19.640 6.325 -19.320 6.645 ;
        RECT -9.720 6.325 -9.400 6.645 ;
        RECT 0.200 6.325 0.520 6.645 ;
        RECT 10.120 6.325 10.440 6.645 ;
        RECT 20.040 6.325 20.360 6.645 ;
        RECT -280.300 5.455 -279.980 5.775 ;
        RECT -279.830 5.455 -279.510 5.775 ;
        RECT -270.380 5.455 -270.060 5.775 ;
        RECT -269.910 5.455 -269.590 5.775 ;
        RECT -260.460 5.455 -260.140 5.775 ;
        RECT -259.990 5.455 -259.670 5.775 ;
        RECT -250.540 5.455 -250.220 5.775 ;
        RECT -250.070 5.455 -249.750 5.775 ;
        RECT -240.620 5.455 -240.300 5.775 ;
        RECT -240.150 5.455 -239.830 5.775 ;
        RECT -230.700 5.455 -230.380 5.775 ;
        RECT -230.230 5.455 -229.910 5.775 ;
        RECT -220.780 5.455 -220.460 5.775 ;
        RECT -220.310 5.455 -219.990 5.775 ;
        RECT -210.860 5.455 -210.540 5.775 ;
        RECT -210.390 5.455 -210.070 5.775 ;
        RECT -200.940 5.455 -200.620 5.775 ;
        RECT -200.470 5.455 -200.150 5.775 ;
        RECT -191.020 5.455 -190.700 5.775 ;
        RECT -190.550 5.455 -190.230 5.775 ;
        RECT -181.100 5.455 -180.780 5.775 ;
        RECT -180.630 5.455 -180.310 5.775 ;
        RECT -171.180 5.455 -170.860 5.775 ;
        RECT -170.710 5.455 -170.390 5.775 ;
        RECT -161.260 5.455 -160.940 5.775 ;
        RECT -160.790 5.455 -160.470 5.775 ;
        RECT -151.340 5.455 -151.020 5.775 ;
        RECT -150.870 5.455 -150.550 5.775 ;
        RECT -141.420 5.455 -141.100 5.775 ;
        RECT -140.950 5.455 -140.630 5.775 ;
        RECT -131.500 5.455 -131.180 5.775 ;
        RECT -131.030 5.455 -130.710 5.775 ;
        RECT -121.580 5.455 -121.260 5.775 ;
        RECT -121.110 5.455 -120.790 5.775 ;
        RECT -111.660 5.455 -111.340 5.775 ;
        RECT -111.190 5.455 -110.870 5.775 ;
        RECT -101.740 5.455 -101.420 5.775 ;
        RECT -101.270 5.455 -100.950 5.775 ;
        RECT -91.820 5.455 -91.500 5.775 ;
        RECT -91.350 5.455 -91.030 5.775 ;
        RECT -81.900 5.455 -81.580 5.775 ;
        RECT -81.430 5.455 -81.110 5.775 ;
        RECT -71.980 5.455 -71.660 5.775 ;
        RECT -71.510 5.455 -71.190 5.775 ;
        RECT -62.060 5.455 -61.740 5.775 ;
        RECT -61.590 5.455 -61.270 5.775 ;
        RECT -52.140 5.455 -51.820 5.775 ;
        RECT -51.670 5.455 -51.350 5.775 ;
        RECT -42.220 5.455 -41.900 5.775 ;
        RECT -41.750 5.455 -41.430 5.775 ;
        RECT -32.300 5.455 -31.980 5.775 ;
        RECT -31.830 5.455 -31.510 5.775 ;
        RECT -22.380 5.455 -22.060 5.775 ;
        RECT -21.910 5.455 -21.590 5.775 ;
        RECT -12.460 5.455 -12.140 5.775 ;
        RECT -11.990 5.455 -11.670 5.775 ;
        RECT -2.540 5.455 -2.220 5.775 ;
        RECT -2.070 5.455 -1.750 5.775 ;
        RECT 7.380 5.455 7.700 5.775 ;
        RECT 7.850 5.455 8.170 5.775 ;
        RECT 17.300 5.455 17.620 5.775 ;
        RECT 17.770 5.455 18.090 5.775 ;
        RECT -287.560 2.735 -287.240 3.055 ;
        RECT -287.100 2.735 -286.780 3.055 ;
        RECT -277.640 2.735 -277.320 3.055 ;
        RECT -277.180 2.735 -276.860 3.055 ;
        RECT -267.720 2.735 -267.400 3.055 ;
        RECT -267.260 2.735 -266.940 3.055 ;
        RECT -257.800 2.735 -257.480 3.055 ;
        RECT -257.340 2.735 -257.020 3.055 ;
        RECT -247.880 2.735 -247.560 3.055 ;
        RECT -247.420 2.735 -247.100 3.055 ;
        RECT -237.960 2.735 -237.640 3.055 ;
        RECT -237.500 2.735 -237.180 3.055 ;
        RECT -228.040 2.735 -227.720 3.055 ;
        RECT -227.580 2.735 -227.260 3.055 ;
        RECT -218.120 2.735 -217.800 3.055 ;
        RECT -217.660 2.735 -217.340 3.055 ;
        RECT -208.200 2.735 -207.880 3.055 ;
        RECT -207.740 2.735 -207.420 3.055 ;
        RECT -198.280 2.735 -197.960 3.055 ;
        RECT -197.820 2.735 -197.500 3.055 ;
        RECT -188.360 2.735 -188.040 3.055 ;
        RECT -187.900 2.735 -187.580 3.055 ;
        RECT -178.440 2.735 -178.120 3.055 ;
        RECT -177.980 2.735 -177.660 3.055 ;
        RECT -168.520 2.735 -168.200 3.055 ;
        RECT -168.060 2.735 -167.740 3.055 ;
        RECT -158.600 2.735 -158.280 3.055 ;
        RECT -158.140 2.735 -157.820 3.055 ;
        RECT -148.680 2.735 -148.360 3.055 ;
        RECT -148.220 2.735 -147.900 3.055 ;
        RECT -138.760 2.735 -138.440 3.055 ;
        RECT -138.300 2.735 -137.980 3.055 ;
        RECT -128.840 2.735 -128.520 3.055 ;
        RECT -128.380 2.735 -128.060 3.055 ;
        RECT -118.920 2.735 -118.600 3.055 ;
        RECT -118.460 2.735 -118.140 3.055 ;
        RECT -109.000 2.735 -108.680 3.055 ;
        RECT -108.540 2.735 -108.220 3.055 ;
        RECT -99.080 2.735 -98.760 3.055 ;
        RECT -98.620 2.735 -98.300 3.055 ;
        RECT -89.160 2.735 -88.840 3.055 ;
        RECT -88.700 2.735 -88.380 3.055 ;
        RECT -79.240 2.735 -78.920 3.055 ;
        RECT -78.780 2.735 -78.460 3.055 ;
        RECT -69.320 2.735 -69.000 3.055 ;
        RECT -68.860 2.735 -68.540 3.055 ;
        RECT -59.400 2.735 -59.080 3.055 ;
        RECT -58.940 2.735 -58.620 3.055 ;
        RECT -49.480 2.735 -49.160 3.055 ;
        RECT -49.020 2.735 -48.700 3.055 ;
        RECT -39.560 2.735 -39.240 3.055 ;
        RECT -39.100 2.735 -38.780 3.055 ;
        RECT -29.640 2.735 -29.320 3.055 ;
        RECT -29.180 2.735 -28.860 3.055 ;
        RECT -19.720 2.735 -19.400 3.055 ;
        RECT -19.260 2.735 -18.940 3.055 ;
        RECT -9.800 2.735 -9.480 3.055 ;
        RECT -9.340 2.735 -9.020 3.055 ;
        RECT 0.120 2.735 0.440 3.055 ;
        RECT 0.580 2.735 0.900 3.055 ;
        RECT 10.040 2.735 10.360 3.055 ;
        RECT 10.500 2.735 10.820 3.055 ;
        RECT 19.960 2.735 20.280 3.055 ;
        RECT 20.420 2.735 20.740 3.055 ;
        RECT -279.910 1.975 -279.590 2.295 ;
        RECT -269.990 1.975 -269.670 2.295 ;
        RECT -260.070 1.975 -259.750 2.295 ;
        RECT -250.150 1.975 -249.830 2.295 ;
        RECT -240.230 1.975 -239.910 2.295 ;
        RECT -230.310 1.975 -229.990 2.295 ;
        RECT -220.390 1.975 -220.070 2.295 ;
        RECT -210.470 1.975 -210.150 2.295 ;
        RECT -200.550 1.975 -200.230 2.295 ;
        RECT -190.630 1.975 -190.310 2.295 ;
        RECT -180.710 1.975 -180.390 2.295 ;
        RECT -170.790 1.975 -170.470 2.295 ;
        RECT -160.870 1.975 -160.550 2.295 ;
        RECT -150.950 1.975 -150.630 2.295 ;
        RECT -141.030 1.975 -140.710 2.295 ;
        RECT -131.110 1.975 -130.790 2.295 ;
        RECT -121.190 1.975 -120.870 2.295 ;
        RECT -111.270 1.975 -110.950 2.295 ;
        RECT -101.350 1.975 -101.030 2.295 ;
        RECT -91.430 1.975 -91.110 2.295 ;
        RECT -81.510 1.975 -81.190 2.295 ;
        RECT -71.590 1.975 -71.270 2.295 ;
        RECT -61.670 1.975 -61.350 2.295 ;
        RECT -51.750 1.975 -51.430 2.295 ;
        RECT -41.830 1.975 -41.510 2.295 ;
        RECT -31.910 1.975 -31.590 2.295 ;
        RECT -21.990 1.975 -21.670 2.295 ;
        RECT -12.070 1.975 -11.750 2.295 ;
        RECT -2.150 1.975 -1.830 2.295 ;
        RECT 7.770 1.975 8.090 2.295 ;
        RECT 17.690 1.975 18.010 2.295 ;
        RECT -285.720 -87.025 -285.400 -86.705 ;
        RECT -275.800 -87.025 -275.480 -86.705 ;
        RECT -265.880 -87.025 -265.560 -86.705 ;
        RECT -255.960 -87.025 -255.640 -86.705 ;
        RECT -246.040 -87.025 -245.720 -86.705 ;
        RECT -236.120 -87.025 -235.800 -86.705 ;
        RECT -226.200 -87.025 -225.880 -86.705 ;
        RECT -216.280 -87.025 -215.960 -86.705 ;
        RECT -206.360 -87.025 -206.040 -86.705 ;
        RECT -196.440 -87.025 -196.120 -86.705 ;
        RECT -186.520 -87.025 -186.200 -86.705 ;
        RECT -176.600 -87.025 -176.280 -86.705 ;
        RECT -166.680 -87.025 -166.360 -86.705 ;
        RECT -156.760 -87.025 -156.440 -86.705 ;
        RECT -146.840 -87.025 -146.520 -86.705 ;
        RECT -136.920 -87.025 -136.600 -86.705 ;
        RECT -127.000 -87.025 -126.680 -86.705 ;
        RECT -117.080 -87.025 -116.760 -86.705 ;
        RECT -107.160 -87.025 -106.840 -86.705 ;
        RECT -97.240 -87.025 -96.920 -86.705 ;
        RECT -87.320 -87.025 -87.000 -86.705 ;
        RECT -77.400 -87.025 -77.080 -86.705 ;
        RECT -67.480 -87.025 -67.160 -86.705 ;
        RECT -57.560 -87.025 -57.240 -86.705 ;
        RECT -47.640 -87.025 -47.320 -86.705 ;
        RECT -37.720 -87.025 -37.400 -86.705 ;
        RECT -27.800 -87.025 -27.480 -86.705 ;
        RECT -17.880 -87.025 -17.560 -86.705 ;
        RECT -7.960 -87.025 -7.640 -86.705 ;
        RECT 1.960 -87.025 2.280 -86.705 ;
        RECT 11.880 -87.025 12.200 -86.705 ;
        RECT 21.800 -87.025 22.120 -86.705 ;
        RECT -278.540 -87.895 -278.220 -87.575 ;
        RECT -278.070 -87.895 -277.750 -87.575 ;
        RECT -268.620 -87.895 -268.300 -87.575 ;
        RECT -268.150 -87.895 -267.830 -87.575 ;
        RECT -258.700 -87.895 -258.380 -87.575 ;
        RECT -258.230 -87.895 -257.910 -87.575 ;
        RECT -248.780 -87.895 -248.460 -87.575 ;
        RECT -248.310 -87.895 -247.990 -87.575 ;
        RECT -238.860 -87.895 -238.540 -87.575 ;
        RECT -238.390 -87.895 -238.070 -87.575 ;
        RECT -228.940 -87.895 -228.620 -87.575 ;
        RECT -228.470 -87.895 -228.150 -87.575 ;
        RECT -219.020 -87.895 -218.700 -87.575 ;
        RECT -218.550 -87.895 -218.230 -87.575 ;
        RECT -209.100 -87.895 -208.780 -87.575 ;
        RECT -208.630 -87.895 -208.310 -87.575 ;
        RECT -199.180 -87.895 -198.860 -87.575 ;
        RECT -198.710 -87.895 -198.390 -87.575 ;
        RECT -189.260 -87.895 -188.940 -87.575 ;
        RECT -188.790 -87.895 -188.470 -87.575 ;
        RECT -179.340 -87.895 -179.020 -87.575 ;
        RECT -178.870 -87.895 -178.550 -87.575 ;
        RECT -169.420 -87.895 -169.100 -87.575 ;
        RECT -168.950 -87.895 -168.630 -87.575 ;
        RECT -159.500 -87.895 -159.180 -87.575 ;
        RECT -159.030 -87.895 -158.710 -87.575 ;
        RECT -149.580 -87.895 -149.260 -87.575 ;
        RECT -149.110 -87.895 -148.790 -87.575 ;
        RECT -139.660 -87.895 -139.340 -87.575 ;
        RECT -139.190 -87.895 -138.870 -87.575 ;
        RECT -129.740 -87.895 -129.420 -87.575 ;
        RECT -129.270 -87.895 -128.950 -87.575 ;
        RECT -119.820 -87.895 -119.500 -87.575 ;
        RECT -119.350 -87.895 -119.030 -87.575 ;
        RECT -109.900 -87.895 -109.580 -87.575 ;
        RECT -109.430 -87.895 -109.110 -87.575 ;
        RECT -99.980 -87.895 -99.660 -87.575 ;
        RECT -99.510 -87.895 -99.190 -87.575 ;
        RECT -90.060 -87.895 -89.740 -87.575 ;
        RECT -89.590 -87.895 -89.270 -87.575 ;
        RECT -80.140 -87.895 -79.820 -87.575 ;
        RECT -79.670 -87.895 -79.350 -87.575 ;
        RECT -70.220 -87.895 -69.900 -87.575 ;
        RECT -69.750 -87.895 -69.430 -87.575 ;
        RECT -60.300 -87.895 -59.980 -87.575 ;
        RECT -59.830 -87.895 -59.510 -87.575 ;
        RECT -50.380 -87.895 -50.060 -87.575 ;
        RECT -49.910 -87.895 -49.590 -87.575 ;
        RECT -40.460 -87.895 -40.140 -87.575 ;
        RECT -39.990 -87.895 -39.670 -87.575 ;
        RECT -30.540 -87.895 -30.220 -87.575 ;
        RECT -30.070 -87.895 -29.750 -87.575 ;
        RECT -20.620 -87.895 -20.300 -87.575 ;
        RECT -20.150 -87.895 -19.830 -87.575 ;
        RECT -10.700 -87.895 -10.380 -87.575 ;
        RECT -10.230 -87.895 -9.910 -87.575 ;
        RECT -0.780 -87.895 -0.460 -87.575 ;
        RECT -0.310 -87.895 0.010 -87.575 ;
        RECT 9.140 -87.895 9.460 -87.575 ;
        RECT 9.610 -87.895 9.930 -87.575 ;
        RECT 19.060 -87.895 19.380 -87.575 ;
        RECT 19.530 -87.895 19.850 -87.575 ;
        RECT -285.800 -90.615 -285.480 -90.295 ;
        RECT -285.340 -90.615 -285.020 -90.295 ;
        RECT -275.880 -90.615 -275.560 -90.295 ;
        RECT -275.420 -90.615 -275.100 -90.295 ;
        RECT -265.960 -90.615 -265.640 -90.295 ;
        RECT -265.500 -90.615 -265.180 -90.295 ;
        RECT -256.040 -90.615 -255.720 -90.295 ;
        RECT -255.580 -90.615 -255.260 -90.295 ;
        RECT -246.120 -90.615 -245.800 -90.295 ;
        RECT -245.660 -90.615 -245.340 -90.295 ;
        RECT -236.200 -90.615 -235.880 -90.295 ;
        RECT -235.740 -90.615 -235.420 -90.295 ;
        RECT -226.280 -90.615 -225.960 -90.295 ;
        RECT -225.820 -90.615 -225.500 -90.295 ;
        RECT -216.360 -90.615 -216.040 -90.295 ;
        RECT -215.900 -90.615 -215.580 -90.295 ;
        RECT -206.440 -90.615 -206.120 -90.295 ;
        RECT -205.980 -90.615 -205.660 -90.295 ;
        RECT -196.520 -90.615 -196.200 -90.295 ;
        RECT -196.060 -90.615 -195.740 -90.295 ;
        RECT -186.600 -90.615 -186.280 -90.295 ;
        RECT -186.140 -90.615 -185.820 -90.295 ;
        RECT -176.680 -90.615 -176.360 -90.295 ;
        RECT -176.220 -90.615 -175.900 -90.295 ;
        RECT -166.760 -90.615 -166.440 -90.295 ;
        RECT -166.300 -90.615 -165.980 -90.295 ;
        RECT -156.840 -90.615 -156.520 -90.295 ;
        RECT -156.380 -90.615 -156.060 -90.295 ;
        RECT -146.920 -90.615 -146.600 -90.295 ;
        RECT -146.460 -90.615 -146.140 -90.295 ;
        RECT -137.000 -90.615 -136.680 -90.295 ;
        RECT -136.540 -90.615 -136.220 -90.295 ;
        RECT -127.080 -90.615 -126.760 -90.295 ;
        RECT -126.620 -90.615 -126.300 -90.295 ;
        RECT -117.160 -90.615 -116.840 -90.295 ;
        RECT -116.700 -90.615 -116.380 -90.295 ;
        RECT -107.240 -90.615 -106.920 -90.295 ;
        RECT -106.780 -90.615 -106.460 -90.295 ;
        RECT -97.320 -90.615 -97.000 -90.295 ;
        RECT -96.860 -90.615 -96.540 -90.295 ;
        RECT -87.400 -90.615 -87.080 -90.295 ;
        RECT -86.940 -90.615 -86.620 -90.295 ;
        RECT -77.480 -90.615 -77.160 -90.295 ;
        RECT -77.020 -90.615 -76.700 -90.295 ;
        RECT -67.560 -90.615 -67.240 -90.295 ;
        RECT -67.100 -90.615 -66.780 -90.295 ;
        RECT -57.640 -90.615 -57.320 -90.295 ;
        RECT -57.180 -90.615 -56.860 -90.295 ;
        RECT -47.720 -90.615 -47.400 -90.295 ;
        RECT -47.260 -90.615 -46.940 -90.295 ;
        RECT -37.800 -90.615 -37.480 -90.295 ;
        RECT -37.340 -90.615 -37.020 -90.295 ;
        RECT -27.880 -90.615 -27.560 -90.295 ;
        RECT -27.420 -90.615 -27.100 -90.295 ;
        RECT -17.960 -90.615 -17.640 -90.295 ;
        RECT -17.500 -90.615 -17.180 -90.295 ;
        RECT -8.040 -90.615 -7.720 -90.295 ;
        RECT -7.580 -90.615 -7.260 -90.295 ;
        RECT 1.880 -90.615 2.200 -90.295 ;
        RECT 2.340 -90.615 2.660 -90.295 ;
        RECT 11.800 -90.615 12.120 -90.295 ;
        RECT 12.260 -90.615 12.580 -90.295 ;
        RECT 21.720 -90.615 22.040 -90.295 ;
        RECT 22.180 -90.615 22.500 -90.295 ;
        RECT -278.150 -91.375 -277.830 -91.055 ;
        RECT -268.230 -91.375 -267.910 -91.055 ;
        RECT -258.310 -91.375 -257.990 -91.055 ;
        RECT -248.390 -91.375 -248.070 -91.055 ;
        RECT -238.470 -91.375 -238.150 -91.055 ;
        RECT -228.550 -91.375 -228.230 -91.055 ;
        RECT -218.630 -91.375 -218.310 -91.055 ;
        RECT -208.710 -91.375 -208.390 -91.055 ;
        RECT -198.790 -91.375 -198.470 -91.055 ;
        RECT -188.870 -91.375 -188.550 -91.055 ;
        RECT -178.950 -91.375 -178.630 -91.055 ;
        RECT -169.030 -91.375 -168.710 -91.055 ;
        RECT -159.110 -91.375 -158.790 -91.055 ;
        RECT -149.190 -91.375 -148.870 -91.055 ;
        RECT -139.270 -91.375 -138.950 -91.055 ;
        RECT -129.350 -91.375 -129.030 -91.055 ;
        RECT -119.430 -91.375 -119.110 -91.055 ;
        RECT -109.510 -91.375 -109.190 -91.055 ;
        RECT -99.590 -91.375 -99.270 -91.055 ;
        RECT -89.670 -91.375 -89.350 -91.055 ;
        RECT -79.750 -91.375 -79.430 -91.055 ;
        RECT -69.830 -91.375 -69.510 -91.055 ;
        RECT -59.910 -91.375 -59.590 -91.055 ;
        RECT -49.990 -91.375 -49.670 -91.055 ;
        RECT -40.070 -91.375 -39.750 -91.055 ;
        RECT -30.150 -91.375 -29.830 -91.055 ;
        RECT -20.230 -91.375 -19.910 -91.055 ;
        RECT -10.310 -91.375 -9.990 -91.055 ;
        RECT -0.390 -91.375 -0.070 -91.055 ;
        RECT 9.530 -91.375 9.850 -91.055 ;
        RECT 19.450 -91.375 19.770 -91.055 ;
        RECT -285.470 -174.735 -285.150 -174.415 ;
        RECT -275.550 -174.735 -275.230 -174.415 ;
        RECT -265.630 -174.735 -265.310 -174.415 ;
        RECT -255.710 -174.735 -255.390 -174.415 ;
        RECT -245.790 -174.735 -245.470 -174.415 ;
        RECT -235.870 -174.735 -235.550 -174.415 ;
        RECT -225.950 -174.735 -225.630 -174.415 ;
        RECT -216.030 -174.735 -215.710 -174.415 ;
        RECT -206.110 -174.735 -205.790 -174.415 ;
        RECT -196.190 -174.735 -195.870 -174.415 ;
        RECT -186.270 -174.735 -185.950 -174.415 ;
        RECT -176.350 -174.735 -176.030 -174.415 ;
        RECT -166.430 -174.735 -166.110 -174.415 ;
        RECT -156.510 -174.735 -156.190 -174.415 ;
        RECT -146.590 -174.735 -146.270 -174.415 ;
        RECT -136.670 -174.735 -136.350 -174.415 ;
        RECT -126.750 -174.735 -126.430 -174.415 ;
        RECT -116.830 -174.735 -116.510 -174.415 ;
        RECT -106.910 -174.735 -106.590 -174.415 ;
        RECT -96.990 -174.735 -96.670 -174.415 ;
        RECT -87.070 -174.735 -86.750 -174.415 ;
        RECT -77.150 -174.735 -76.830 -174.415 ;
        RECT -67.230 -174.735 -66.910 -174.415 ;
        RECT -57.310 -174.735 -56.990 -174.415 ;
        RECT -47.390 -174.735 -47.070 -174.415 ;
        RECT -37.470 -174.735 -37.150 -174.415 ;
        RECT -27.550 -174.735 -27.230 -174.415 ;
        RECT -17.630 -174.735 -17.310 -174.415 ;
        RECT -7.710 -174.735 -7.390 -174.415 ;
        RECT 2.210 -174.735 2.530 -174.415 ;
        RECT 12.130 -174.735 12.450 -174.415 ;
        RECT 22.050 -174.735 22.370 -174.415 ;
        RECT -278.290 -175.605 -277.970 -175.285 ;
        RECT -277.820 -175.605 -277.500 -175.285 ;
        RECT -268.370 -175.605 -268.050 -175.285 ;
        RECT -267.900 -175.605 -267.580 -175.285 ;
        RECT -258.450 -175.605 -258.130 -175.285 ;
        RECT -257.980 -175.605 -257.660 -175.285 ;
        RECT -248.530 -175.605 -248.210 -175.285 ;
        RECT -248.060 -175.605 -247.740 -175.285 ;
        RECT -238.610 -175.605 -238.290 -175.285 ;
        RECT -238.140 -175.605 -237.820 -175.285 ;
        RECT -228.690 -175.605 -228.370 -175.285 ;
        RECT -228.220 -175.605 -227.900 -175.285 ;
        RECT -218.770 -175.605 -218.450 -175.285 ;
        RECT -218.300 -175.605 -217.980 -175.285 ;
        RECT -208.850 -175.605 -208.530 -175.285 ;
        RECT -208.380 -175.605 -208.060 -175.285 ;
        RECT -198.930 -175.605 -198.610 -175.285 ;
        RECT -198.460 -175.605 -198.140 -175.285 ;
        RECT -189.010 -175.605 -188.690 -175.285 ;
        RECT -188.540 -175.605 -188.220 -175.285 ;
        RECT -179.090 -175.605 -178.770 -175.285 ;
        RECT -178.620 -175.605 -178.300 -175.285 ;
        RECT -169.170 -175.605 -168.850 -175.285 ;
        RECT -168.700 -175.605 -168.380 -175.285 ;
        RECT -159.250 -175.605 -158.930 -175.285 ;
        RECT -158.780 -175.605 -158.460 -175.285 ;
        RECT -149.330 -175.605 -149.010 -175.285 ;
        RECT -148.860 -175.605 -148.540 -175.285 ;
        RECT -139.410 -175.605 -139.090 -175.285 ;
        RECT -138.940 -175.605 -138.620 -175.285 ;
        RECT -129.490 -175.605 -129.170 -175.285 ;
        RECT -129.020 -175.605 -128.700 -175.285 ;
        RECT -119.570 -175.605 -119.250 -175.285 ;
        RECT -119.100 -175.605 -118.780 -175.285 ;
        RECT -109.650 -175.605 -109.330 -175.285 ;
        RECT -109.180 -175.605 -108.860 -175.285 ;
        RECT -99.730 -175.605 -99.410 -175.285 ;
        RECT -99.260 -175.605 -98.940 -175.285 ;
        RECT -89.810 -175.605 -89.490 -175.285 ;
        RECT -89.340 -175.605 -89.020 -175.285 ;
        RECT -79.890 -175.605 -79.570 -175.285 ;
        RECT -79.420 -175.605 -79.100 -175.285 ;
        RECT -69.970 -175.605 -69.650 -175.285 ;
        RECT -69.500 -175.605 -69.180 -175.285 ;
        RECT -60.050 -175.605 -59.730 -175.285 ;
        RECT -59.580 -175.605 -59.260 -175.285 ;
        RECT -50.130 -175.605 -49.810 -175.285 ;
        RECT -49.660 -175.605 -49.340 -175.285 ;
        RECT -40.210 -175.605 -39.890 -175.285 ;
        RECT -39.740 -175.605 -39.420 -175.285 ;
        RECT -30.290 -175.605 -29.970 -175.285 ;
        RECT -29.820 -175.605 -29.500 -175.285 ;
        RECT -20.370 -175.605 -20.050 -175.285 ;
        RECT -19.900 -175.605 -19.580 -175.285 ;
        RECT -10.450 -175.605 -10.130 -175.285 ;
        RECT -9.980 -175.605 -9.660 -175.285 ;
        RECT -0.530 -175.605 -0.210 -175.285 ;
        RECT -0.060 -175.605 0.260 -175.285 ;
        RECT 9.390 -175.605 9.710 -175.285 ;
        RECT 9.860 -175.605 10.180 -175.285 ;
        RECT 19.310 -175.605 19.630 -175.285 ;
        RECT 19.780 -175.605 20.100 -175.285 ;
        RECT -285.550 -178.325 -285.230 -178.005 ;
        RECT -285.090 -178.325 -284.770 -178.005 ;
        RECT -275.630 -178.325 -275.310 -178.005 ;
        RECT -275.170 -178.325 -274.850 -178.005 ;
        RECT -265.710 -178.325 -265.390 -178.005 ;
        RECT -265.250 -178.325 -264.930 -178.005 ;
        RECT -255.790 -178.325 -255.470 -178.005 ;
        RECT -255.330 -178.325 -255.010 -178.005 ;
        RECT -245.870 -178.325 -245.550 -178.005 ;
        RECT -245.410 -178.325 -245.090 -178.005 ;
        RECT -235.950 -178.325 -235.630 -178.005 ;
        RECT -235.490 -178.325 -235.170 -178.005 ;
        RECT -226.030 -178.325 -225.710 -178.005 ;
        RECT -225.570 -178.325 -225.250 -178.005 ;
        RECT -216.110 -178.325 -215.790 -178.005 ;
        RECT -215.650 -178.325 -215.330 -178.005 ;
        RECT -206.190 -178.325 -205.870 -178.005 ;
        RECT -205.730 -178.325 -205.410 -178.005 ;
        RECT -196.270 -178.325 -195.950 -178.005 ;
        RECT -195.810 -178.325 -195.490 -178.005 ;
        RECT -186.350 -178.325 -186.030 -178.005 ;
        RECT -185.890 -178.325 -185.570 -178.005 ;
        RECT -176.430 -178.325 -176.110 -178.005 ;
        RECT -175.970 -178.325 -175.650 -178.005 ;
        RECT -166.510 -178.325 -166.190 -178.005 ;
        RECT -166.050 -178.325 -165.730 -178.005 ;
        RECT -156.590 -178.325 -156.270 -178.005 ;
        RECT -156.130 -178.325 -155.810 -178.005 ;
        RECT -146.670 -178.325 -146.350 -178.005 ;
        RECT -146.210 -178.325 -145.890 -178.005 ;
        RECT -136.750 -178.325 -136.430 -178.005 ;
        RECT -136.290 -178.325 -135.970 -178.005 ;
        RECT -126.830 -178.325 -126.510 -178.005 ;
        RECT -126.370 -178.325 -126.050 -178.005 ;
        RECT -116.910 -178.325 -116.590 -178.005 ;
        RECT -116.450 -178.325 -116.130 -178.005 ;
        RECT -106.990 -178.325 -106.670 -178.005 ;
        RECT -106.530 -178.325 -106.210 -178.005 ;
        RECT -97.070 -178.325 -96.750 -178.005 ;
        RECT -96.610 -178.325 -96.290 -178.005 ;
        RECT -87.150 -178.325 -86.830 -178.005 ;
        RECT -86.690 -178.325 -86.370 -178.005 ;
        RECT -77.230 -178.325 -76.910 -178.005 ;
        RECT -76.770 -178.325 -76.450 -178.005 ;
        RECT -67.310 -178.325 -66.990 -178.005 ;
        RECT -66.850 -178.325 -66.530 -178.005 ;
        RECT -57.390 -178.325 -57.070 -178.005 ;
        RECT -56.930 -178.325 -56.610 -178.005 ;
        RECT -47.470 -178.325 -47.150 -178.005 ;
        RECT -47.010 -178.325 -46.690 -178.005 ;
        RECT -37.550 -178.325 -37.230 -178.005 ;
        RECT -37.090 -178.325 -36.770 -178.005 ;
        RECT -27.630 -178.325 -27.310 -178.005 ;
        RECT -27.170 -178.325 -26.850 -178.005 ;
        RECT -17.710 -178.325 -17.390 -178.005 ;
        RECT -17.250 -178.325 -16.930 -178.005 ;
        RECT -7.790 -178.325 -7.470 -178.005 ;
        RECT -7.330 -178.325 -7.010 -178.005 ;
        RECT 2.130 -178.325 2.450 -178.005 ;
        RECT 2.590 -178.325 2.910 -178.005 ;
        RECT 12.050 -178.325 12.370 -178.005 ;
        RECT 12.510 -178.325 12.830 -178.005 ;
        RECT 21.970 -178.325 22.290 -178.005 ;
        RECT 22.430 -178.325 22.750 -178.005 ;
        RECT -277.900 -179.085 -277.580 -178.765 ;
        RECT -267.980 -179.085 -267.660 -178.765 ;
        RECT -258.060 -179.085 -257.740 -178.765 ;
        RECT -248.140 -179.085 -247.820 -178.765 ;
        RECT -238.220 -179.085 -237.900 -178.765 ;
        RECT -228.300 -179.085 -227.980 -178.765 ;
        RECT -218.380 -179.085 -218.060 -178.765 ;
        RECT -208.460 -179.085 -208.140 -178.765 ;
        RECT -198.540 -179.085 -198.220 -178.765 ;
        RECT -188.620 -179.085 -188.300 -178.765 ;
        RECT -178.700 -179.085 -178.380 -178.765 ;
        RECT -168.780 -179.085 -168.460 -178.765 ;
        RECT -158.860 -179.085 -158.540 -178.765 ;
        RECT -148.940 -179.085 -148.620 -178.765 ;
        RECT -139.020 -179.085 -138.700 -178.765 ;
        RECT -129.100 -179.085 -128.780 -178.765 ;
        RECT -119.180 -179.085 -118.860 -178.765 ;
        RECT -109.260 -179.085 -108.940 -178.765 ;
        RECT -99.340 -179.085 -99.020 -178.765 ;
        RECT -89.420 -179.085 -89.100 -178.765 ;
        RECT -79.500 -179.085 -79.180 -178.765 ;
        RECT -69.580 -179.085 -69.260 -178.765 ;
        RECT -59.660 -179.085 -59.340 -178.765 ;
        RECT -49.740 -179.085 -49.420 -178.765 ;
        RECT -39.820 -179.085 -39.500 -178.765 ;
        RECT -29.900 -179.085 -29.580 -178.765 ;
        RECT -19.980 -179.085 -19.660 -178.765 ;
        RECT -10.060 -179.085 -9.740 -178.765 ;
        RECT -0.140 -179.085 0.180 -178.765 ;
        RECT 9.780 -179.085 10.100 -178.765 ;
        RECT 19.700 -179.085 20.020 -178.765 ;
      LAYER met4 ;
        RECT -361.230 94.570 -353.030 94.740 ;
        RECT -361.230 94.560 -296.360 94.570 ;
        RECT -366.890 91.100 68.120 94.560 ;
        RECT -367.230 89.390 68.120 91.100 ;
        RECT -367.230 89.340 -296.360 89.390 ;
        RECT -367.230 89.330 -308.360 89.340 ;
        RECT -367.230 6.730 -353.030 89.330 ;
        RECT -300.990 6.730 68.370 6.850 ;
        RECT -367.230 1.680 68.370 6.730 ;
        RECT -367.230 1.500 -297.140 1.680 ;
        RECT -367.230 -86.450 -353.030 1.500 ;
        RECT -367.230 -86.510 -302.700 -86.450 ;
        RECT -299.230 -86.510 70.130 -86.500 ;
        RECT -367.230 -91.670 70.130 -86.510 ;
        RECT -367.230 -91.740 -294.800 -91.670 ;
        RECT -367.230 -174.010 -353.030 -91.740 ;
        RECT -367.230 -174.210 -297.960 -174.010 ;
        RECT -367.230 -179.060 70.380 -174.210 ;
        RECT -363.590 -179.240 70.380 -179.060 ;
        RECT -361.230 -179.420 -353.030 -179.240 ;
        RECT -307.960 -179.380 70.380 -179.240 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -283.195 93.570 -279.425 95.330 ;
        RECT -273.275 93.570 -269.505 95.330 ;
        RECT -263.355 93.570 -259.585 95.330 ;
        RECT -253.435 93.570 -249.665 95.330 ;
        RECT -243.515 93.570 -239.745 95.330 ;
        RECT -233.595 93.570 -229.825 95.330 ;
        RECT -223.675 93.570 -219.905 95.330 ;
        RECT -213.755 93.570 -209.985 95.330 ;
        RECT -203.835 93.570 -200.065 95.330 ;
        RECT -193.915 93.570 -190.145 95.330 ;
        RECT -183.995 93.570 -180.225 95.330 ;
        RECT -174.075 93.570 -170.305 95.330 ;
        RECT -164.155 93.570 -160.385 95.330 ;
        RECT -154.235 93.570 -150.465 95.330 ;
        RECT -144.315 93.570 -140.545 95.330 ;
        RECT -134.395 93.570 -130.625 95.330 ;
        RECT -124.475 93.570 -120.705 95.330 ;
        RECT -114.555 93.570 -110.785 95.330 ;
        RECT -104.635 93.570 -100.865 95.330 ;
        RECT -94.715 93.570 -90.945 95.330 ;
        RECT -84.795 93.570 -81.025 95.330 ;
        RECT -74.875 93.570 -71.105 95.330 ;
        RECT -64.955 93.570 -61.185 95.330 ;
        RECT -55.035 93.570 -51.265 95.330 ;
        RECT -45.115 93.570 -41.345 95.330 ;
        RECT -35.195 93.570 -31.425 95.330 ;
        RECT -25.275 93.570 -21.505 95.330 ;
        RECT -15.355 93.570 -11.585 95.330 ;
        RECT -5.435 93.570 -1.665 95.330 ;
        RECT 4.485 93.570 8.255 95.330 ;
        RECT 14.405 93.570 18.175 95.330 ;
        RECT 24.325 95.095 25.930 95.330 ;
        RECT 24.325 95.090 26.440 95.095 ;
        RECT 24.325 93.570 26.630 95.090 ;
        RECT -281.730 93.520 -280.890 93.570 ;
        RECT -288.070 91.915 -284.470 93.520 ;
        RECT -283.110 90.420 -279.510 92.025 ;
        RECT -278.150 91.915 -274.550 93.520 ;
        RECT -271.810 93.510 -270.970 93.570 ;
        RECT -261.890 93.520 -261.050 93.570 ;
        RECT -273.190 90.420 -269.590 92.025 ;
        RECT -268.230 91.915 -264.630 93.520 ;
        RECT -263.270 90.420 -259.670 92.025 ;
        RECT -258.310 91.915 -254.710 93.520 ;
        RECT -251.970 93.510 -251.130 93.570 ;
        RECT -242.050 93.520 -241.210 93.570 ;
        RECT -253.350 90.420 -249.750 92.025 ;
        RECT -248.390 91.915 -244.790 93.520 ;
        RECT -243.430 90.420 -239.830 92.025 ;
        RECT -238.470 91.915 -234.870 93.520 ;
        RECT -232.130 93.510 -231.290 93.570 ;
        RECT -222.210 93.520 -221.370 93.570 ;
        RECT -233.510 90.420 -229.910 92.025 ;
        RECT -228.550 91.915 -224.950 93.520 ;
        RECT -223.590 90.420 -219.990 92.025 ;
        RECT -218.630 91.915 -215.030 93.520 ;
        RECT -212.290 93.510 -211.450 93.570 ;
        RECT -202.370 93.520 -201.530 93.570 ;
        RECT -213.670 90.420 -210.070 92.025 ;
        RECT -208.710 91.915 -205.110 93.520 ;
        RECT -203.750 90.420 -200.150 92.025 ;
        RECT -198.790 91.915 -195.190 93.520 ;
        RECT -192.450 93.510 -191.610 93.570 ;
        RECT -182.530 93.520 -181.690 93.570 ;
        RECT -193.830 90.420 -190.230 92.025 ;
        RECT -188.870 91.915 -185.270 93.520 ;
        RECT -183.910 90.420 -180.310 92.025 ;
        RECT -178.950 91.915 -175.350 93.520 ;
        RECT -172.610 93.510 -171.770 93.570 ;
        RECT -162.690 93.520 -161.850 93.570 ;
        RECT -173.990 90.420 -170.390 92.025 ;
        RECT -169.030 91.915 -165.430 93.520 ;
        RECT -164.070 90.420 -160.470 92.025 ;
        RECT -159.110 91.915 -155.510 93.520 ;
        RECT -152.770 93.510 -151.930 93.570 ;
        RECT -142.850 93.520 -142.010 93.570 ;
        RECT -154.150 90.420 -150.550 92.025 ;
        RECT -149.190 91.915 -145.590 93.520 ;
        RECT -144.230 90.420 -140.630 92.025 ;
        RECT -139.270 91.915 -135.670 93.520 ;
        RECT -132.930 93.510 -132.090 93.570 ;
        RECT -123.010 93.520 -122.170 93.570 ;
        RECT -134.310 90.420 -130.710 92.025 ;
        RECT -129.350 91.915 -125.750 93.520 ;
        RECT -124.390 90.420 -120.790 92.025 ;
        RECT -119.430 91.915 -115.830 93.520 ;
        RECT -113.090 93.510 -112.250 93.570 ;
        RECT -103.170 93.520 -102.330 93.570 ;
        RECT -114.470 90.420 -110.870 92.025 ;
        RECT -109.510 91.915 -105.910 93.520 ;
        RECT -104.550 90.420 -100.950 92.025 ;
        RECT -99.590 91.915 -95.990 93.520 ;
        RECT -93.250 93.510 -92.410 93.570 ;
        RECT -83.330 93.520 -82.490 93.570 ;
        RECT -94.630 90.420 -91.030 92.025 ;
        RECT -89.670 91.915 -86.070 93.520 ;
        RECT -84.710 90.420 -81.110 92.025 ;
        RECT -79.750 91.915 -76.150 93.520 ;
        RECT -73.410 93.510 -72.570 93.570 ;
        RECT -63.490 93.520 -62.650 93.570 ;
        RECT -74.790 90.420 -71.190 92.025 ;
        RECT -69.830 91.915 -66.230 93.520 ;
        RECT -64.870 90.420 -61.270 92.025 ;
        RECT -59.910 91.915 -56.310 93.520 ;
        RECT -53.570 93.510 -52.730 93.570 ;
        RECT -43.650 93.520 -42.810 93.570 ;
        RECT -54.950 90.420 -51.350 92.025 ;
        RECT -49.990 91.915 -46.390 93.520 ;
        RECT -45.030 90.420 -41.430 92.025 ;
        RECT -40.070 91.915 -36.470 93.520 ;
        RECT -33.730 93.510 -32.890 93.570 ;
        RECT -23.810 93.520 -22.970 93.570 ;
        RECT -35.110 90.420 -31.510 92.025 ;
        RECT -30.150 91.915 -26.550 93.520 ;
        RECT -25.190 90.420 -21.590 92.025 ;
        RECT -20.230 91.915 -16.630 93.520 ;
        RECT -13.890 93.510 -13.050 93.570 ;
        RECT -3.970 93.520 -3.130 93.570 ;
        RECT -15.270 90.420 -11.670 92.025 ;
        RECT -10.310 91.915 -6.710 93.520 ;
        RECT -5.350 90.420 -1.750 92.025 ;
        RECT -0.390 91.915 3.210 93.520 ;
        RECT 5.950 93.510 6.790 93.570 ;
        RECT 15.870 93.520 16.710 93.570 ;
        RECT 25.790 93.520 26.630 93.570 ;
        RECT 4.570 90.420 8.170 92.025 ;
        RECT 9.530 91.915 13.130 93.520 ;
        RECT 14.490 90.420 18.090 92.025 ;
        RECT 19.450 91.915 23.050 93.520 ;
        RECT 24.410 90.420 26.630 92.025 ;
        RECT -288.155 88.610 -284.385 90.370 ;
        RECT -278.235 88.610 -274.465 90.370 ;
        RECT -268.315 88.610 -264.545 90.370 ;
        RECT -258.395 88.610 -254.625 90.370 ;
        RECT -248.475 88.610 -244.705 90.370 ;
        RECT -238.555 88.610 -234.785 90.370 ;
        RECT -228.635 88.610 -224.865 90.370 ;
        RECT -218.715 88.610 -214.945 90.370 ;
        RECT -208.795 88.610 -205.025 90.370 ;
        RECT -198.875 88.610 -195.105 90.370 ;
        RECT -188.955 88.610 -185.185 90.370 ;
        RECT -179.035 88.610 -175.265 90.370 ;
        RECT -169.115 88.610 -165.345 90.370 ;
        RECT -159.195 88.610 -155.425 90.370 ;
        RECT -149.275 88.610 -145.505 90.370 ;
        RECT -139.355 88.610 -135.585 90.370 ;
        RECT -129.435 88.610 -125.665 90.370 ;
        RECT -119.515 88.610 -115.745 90.370 ;
        RECT -109.595 88.610 -105.825 90.370 ;
        RECT -99.675 88.610 -95.905 90.370 ;
        RECT -89.755 88.610 -85.985 90.370 ;
        RECT -79.835 88.610 -76.065 90.370 ;
        RECT -69.915 88.610 -66.145 90.370 ;
        RECT -59.995 88.610 -56.225 90.370 ;
        RECT -50.075 88.610 -46.305 90.370 ;
        RECT -40.155 88.610 -36.385 90.370 ;
        RECT -30.235 88.610 -26.465 90.370 ;
        RECT -20.315 88.610 -16.545 90.370 ;
        RECT -10.395 88.610 -6.625 90.370 ;
        RECT -0.475 88.610 3.295 90.370 ;
        RECT 9.445 88.610 13.215 90.370 ;
        RECT 19.365 88.610 23.135 90.370 ;
        RECT -282.945 5.860 -279.175 7.620 ;
        RECT -273.025 5.860 -269.255 7.620 ;
        RECT -263.105 5.860 -259.335 7.620 ;
        RECT -253.185 5.860 -249.415 7.620 ;
        RECT -243.265 5.860 -239.495 7.620 ;
        RECT -233.345 5.860 -229.575 7.620 ;
        RECT -223.425 5.860 -219.655 7.620 ;
        RECT -213.505 5.860 -209.735 7.620 ;
        RECT -203.585 5.860 -199.815 7.620 ;
        RECT -193.665 5.860 -189.895 7.620 ;
        RECT -183.745 5.860 -179.975 7.620 ;
        RECT -173.825 5.860 -170.055 7.620 ;
        RECT -163.905 5.860 -160.135 7.620 ;
        RECT -153.985 5.860 -150.215 7.620 ;
        RECT -144.065 5.860 -140.295 7.620 ;
        RECT -134.145 5.860 -130.375 7.620 ;
        RECT -124.225 5.860 -120.455 7.620 ;
        RECT -114.305 5.860 -110.535 7.620 ;
        RECT -104.385 5.860 -100.615 7.620 ;
        RECT -94.465 5.860 -90.695 7.620 ;
        RECT -84.545 5.860 -80.775 7.620 ;
        RECT -74.625 5.860 -70.855 7.620 ;
        RECT -64.705 5.860 -60.935 7.620 ;
        RECT -54.785 5.860 -51.015 7.620 ;
        RECT -44.865 5.860 -41.095 7.620 ;
        RECT -34.945 5.860 -31.175 7.620 ;
        RECT -25.025 5.860 -21.255 7.620 ;
        RECT -15.105 5.860 -11.335 7.620 ;
        RECT -5.185 5.860 -1.415 7.620 ;
        RECT 4.735 5.860 8.505 7.620 ;
        RECT 14.655 5.860 18.425 7.620 ;
        RECT 24.575 7.385 26.180 7.620 ;
        RECT 24.575 7.380 26.690 7.385 ;
        RECT 24.575 5.860 26.880 7.380 ;
        RECT -281.480 5.810 -280.640 5.860 ;
        RECT -287.820 4.205 -284.220 5.810 ;
        RECT -282.860 2.710 -279.260 4.315 ;
        RECT -277.900 4.205 -274.300 5.810 ;
        RECT -271.560 5.800 -270.720 5.860 ;
        RECT -261.640 5.810 -260.800 5.860 ;
        RECT -272.940 2.710 -269.340 4.315 ;
        RECT -267.980 4.205 -264.380 5.810 ;
        RECT -263.020 2.710 -259.420 4.315 ;
        RECT -258.060 4.205 -254.460 5.810 ;
        RECT -251.720 5.800 -250.880 5.860 ;
        RECT -241.800 5.810 -240.960 5.860 ;
        RECT -253.100 2.710 -249.500 4.315 ;
        RECT -248.140 4.205 -244.540 5.810 ;
        RECT -243.180 2.710 -239.580 4.315 ;
        RECT -238.220 4.205 -234.620 5.810 ;
        RECT -231.880 5.800 -231.040 5.860 ;
        RECT -221.960 5.810 -221.120 5.860 ;
        RECT -233.260 2.710 -229.660 4.315 ;
        RECT -228.300 4.205 -224.700 5.810 ;
        RECT -223.340 2.710 -219.740 4.315 ;
        RECT -218.380 4.205 -214.780 5.810 ;
        RECT -212.040 5.800 -211.200 5.860 ;
        RECT -202.120 5.810 -201.280 5.860 ;
        RECT -213.420 2.710 -209.820 4.315 ;
        RECT -208.460 4.205 -204.860 5.810 ;
        RECT -203.500 2.710 -199.900 4.315 ;
        RECT -198.540 4.205 -194.940 5.810 ;
        RECT -192.200 5.800 -191.360 5.860 ;
        RECT -182.280 5.810 -181.440 5.860 ;
        RECT -193.580 2.710 -189.980 4.315 ;
        RECT -188.620 4.205 -185.020 5.810 ;
        RECT -183.660 2.710 -180.060 4.315 ;
        RECT -178.700 4.205 -175.100 5.810 ;
        RECT -172.360 5.800 -171.520 5.860 ;
        RECT -162.440 5.810 -161.600 5.860 ;
        RECT -173.740 2.710 -170.140 4.315 ;
        RECT -168.780 4.205 -165.180 5.810 ;
        RECT -163.820 2.710 -160.220 4.315 ;
        RECT -158.860 4.205 -155.260 5.810 ;
        RECT -152.520 5.800 -151.680 5.860 ;
        RECT -142.600 5.810 -141.760 5.860 ;
        RECT -153.900 2.710 -150.300 4.315 ;
        RECT -148.940 4.205 -145.340 5.810 ;
        RECT -143.980 2.710 -140.380 4.315 ;
        RECT -139.020 4.205 -135.420 5.810 ;
        RECT -132.680 5.800 -131.840 5.860 ;
        RECT -122.760 5.810 -121.920 5.860 ;
        RECT -134.060 2.710 -130.460 4.315 ;
        RECT -129.100 4.205 -125.500 5.810 ;
        RECT -124.140 2.710 -120.540 4.315 ;
        RECT -119.180 4.205 -115.580 5.810 ;
        RECT -112.840 5.800 -112.000 5.860 ;
        RECT -102.920 5.810 -102.080 5.860 ;
        RECT -114.220 2.710 -110.620 4.315 ;
        RECT -109.260 4.205 -105.660 5.810 ;
        RECT -104.300 2.710 -100.700 4.315 ;
        RECT -99.340 4.205 -95.740 5.810 ;
        RECT -93.000 5.800 -92.160 5.860 ;
        RECT -83.080 5.810 -82.240 5.860 ;
        RECT -94.380 2.710 -90.780 4.315 ;
        RECT -89.420 4.205 -85.820 5.810 ;
        RECT -84.460 2.710 -80.860 4.315 ;
        RECT -79.500 4.205 -75.900 5.810 ;
        RECT -73.160 5.800 -72.320 5.860 ;
        RECT -63.240 5.810 -62.400 5.860 ;
        RECT -74.540 2.710 -70.940 4.315 ;
        RECT -69.580 4.205 -65.980 5.810 ;
        RECT -64.620 2.710 -61.020 4.315 ;
        RECT -59.660 4.205 -56.060 5.810 ;
        RECT -53.320 5.800 -52.480 5.860 ;
        RECT -43.400 5.810 -42.560 5.860 ;
        RECT -54.700 2.710 -51.100 4.315 ;
        RECT -49.740 4.205 -46.140 5.810 ;
        RECT -44.780 2.710 -41.180 4.315 ;
        RECT -39.820 4.205 -36.220 5.810 ;
        RECT -33.480 5.800 -32.640 5.860 ;
        RECT -23.560 5.810 -22.720 5.860 ;
        RECT -34.860 2.710 -31.260 4.315 ;
        RECT -29.900 4.205 -26.300 5.810 ;
        RECT -24.940 2.710 -21.340 4.315 ;
        RECT -19.980 4.205 -16.380 5.810 ;
        RECT -13.640 5.800 -12.800 5.860 ;
        RECT -3.720 5.810 -2.880 5.860 ;
        RECT -15.020 2.710 -11.420 4.315 ;
        RECT -10.060 4.205 -6.460 5.810 ;
        RECT -5.100 2.710 -1.500 4.315 ;
        RECT -0.140 4.205 3.460 5.810 ;
        RECT 6.200 5.800 7.040 5.860 ;
        RECT 16.120 5.810 16.960 5.860 ;
        RECT 26.040 5.810 26.880 5.860 ;
        RECT 4.820 2.710 8.420 4.315 ;
        RECT 9.780 4.205 13.380 5.810 ;
        RECT 14.740 2.710 18.340 4.315 ;
        RECT 19.700 4.205 23.300 5.810 ;
        RECT 24.660 2.710 26.880 4.315 ;
        RECT -287.905 0.900 -284.135 2.660 ;
        RECT -277.985 0.900 -274.215 2.660 ;
        RECT -268.065 0.900 -264.295 2.660 ;
        RECT -258.145 0.900 -254.375 2.660 ;
        RECT -248.225 0.900 -244.455 2.660 ;
        RECT -238.305 0.900 -234.535 2.660 ;
        RECT -228.385 0.900 -224.615 2.660 ;
        RECT -218.465 0.900 -214.695 2.660 ;
        RECT -208.545 0.900 -204.775 2.660 ;
        RECT -198.625 0.900 -194.855 2.660 ;
        RECT -188.705 0.900 -184.935 2.660 ;
        RECT -178.785 0.900 -175.015 2.660 ;
        RECT -168.865 0.900 -165.095 2.660 ;
        RECT -158.945 0.900 -155.175 2.660 ;
        RECT -149.025 0.900 -145.255 2.660 ;
        RECT -139.105 0.900 -135.335 2.660 ;
        RECT -129.185 0.900 -125.415 2.660 ;
        RECT -119.265 0.900 -115.495 2.660 ;
        RECT -109.345 0.900 -105.575 2.660 ;
        RECT -99.425 0.900 -95.655 2.660 ;
        RECT -89.505 0.900 -85.735 2.660 ;
        RECT -79.585 0.900 -75.815 2.660 ;
        RECT -69.665 0.900 -65.895 2.660 ;
        RECT -59.745 0.900 -55.975 2.660 ;
        RECT -49.825 0.900 -46.055 2.660 ;
        RECT -39.905 0.900 -36.135 2.660 ;
        RECT -29.985 0.900 -26.215 2.660 ;
        RECT -20.065 0.900 -16.295 2.660 ;
        RECT -10.145 0.900 -6.375 2.660 ;
        RECT -0.225 0.900 3.545 2.660 ;
        RECT 9.695 0.900 13.465 2.660 ;
        RECT 19.615 0.900 23.385 2.660 ;
        RECT -281.185 -87.490 -277.415 -85.730 ;
        RECT -271.265 -87.490 -267.495 -85.730 ;
        RECT -261.345 -87.490 -257.575 -85.730 ;
        RECT -251.425 -87.490 -247.655 -85.730 ;
        RECT -241.505 -87.490 -237.735 -85.730 ;
        RECT -231.585 -87.490 -227.815 -85.730 ;
        RECT -221.665 -87.490 -217.895 -85.730 ;
        RECT -211.745 -87.490 -207.975 -85.730 ;
        RECT -201.825 -87.490 -198.055 -85.730 ;
        RECT -191.905 -87.490 -188.135 -85.730 ;
        RECT -181.985 -87.490 -178.215 -85.730 ;
        RECT -172.065 -87.490 -168.295 -85.730 ;
        RECT -162.145 -87.490 -158.375 -85.730 ;
        RECT -152.225 -87.490 -148.455 -85.730 ;
        RECT -142.305 -87.490 -138.535 -85.730 ;
        RECT -132.385 -87.490 -128.615 -85.730 ;
        RECT -122.465 -87.490 -118.695 -85.730 ;
        RECT -112.545 -87.490 -108.775 -85.730 ;
        RECT -102.625 -87.490 -98.855 -85.730 ;
        RECT -92.705 -87.490 -88.935 -85.730 ;
        RECT -82.785 -87.490 -79.015 -85.730 ;
        RECT -72.865 -87.490 -69.095 -85.730 ;
        RECT -62.945 -87.490 -59.175 -85.730 ;
        RECT -53.025 -87.490 -49.255 -85.730 ;
        RECT -43.105 -87.490 -39.335 -85.730 ;
        RECT -33.185 -87.490 -29.415 -85.730 ;
        RECT -23.265 -87.490 -19.495 -85.730 ;
        RECT -13.345 -87.490 -9.575 -85.730 ;
        RECT -3.425 -87.490 0.345 -85.730 ;
        RECT 6.495 -87.490 10.265 -85.730 ;
        RECT 16.415 -87.490 20.185 -85.730 ;
        RECT 26.335 -85.965 27.940 -85.730 ;
        RECT 26.335 -85.970 28.450 -85.965 ;
        RECT 26.335 -87.490 28.640 -85.970 ;
        RECT -279.720 -87.540 -278.880 -87.490 ;
        RECT -286.060 -89.145 -282.460 -87.540 ;
        RECT -281.100 -90.640 -277.500 -89.035 ;
        RECT -276.140 -89.145 -272.540 -87.540 ;
        RECT -269.800 -87.550 -268.960 -87.490 ;
        RECT -259.880 -87.540 -259.040 -87.490 ;
        RECT -271.180 -90.640 -267.580 -89.035 ;
        RECT -266.220 -89.145 -262.620 -87.540 ;
        RECT -261.260 -90.640 -257.660 -89.035 ;
        RECT -256.300 -89.145 -252.700 -87.540 ;
        RECT -249.960 -87.550 -249.120 -87.490 ;
        RECT -240.040 -87.540 -239.200 -87.490 ;
        RECT -251.340 -90.640 -247.740 -89.035 ;
        RECT -246.380 -89.145 -242.780 -87.540 ;
        RECT -241.420 -90.640 -237.820 -89.035 ;
        RECT -236.460 -89.145 -232.860 -87.540 ;
        RECT -230.120 -87.550 -229.280 -87.490 ;
        RECT -220.200 -87.540 -219.360 -87.490 ;
        RECT -231.500 -90.640 -227.900 -89.035 ;
        RECT -226.540 -89.145 -222.940 -87.540 ;
        RECT -221.580 -90.640 -217.980 -89.035 ;
        RECT -216.620 -89.145 -213.020 -87.540 ;
        RECT -210.280 -87.550 -209.440 -87.490 ;
        RECT -200.360 -87.540 -199.520 -87.490 ;
        RECT -211.660 -90.640 -208.060 -89.035 ;
        RECT -206.700 -89.145 -203.100 -87.540 ;
        RECT -201.740 -90.640 -198.140 -89.035 ;
        RECT -196.780 -89.145 -193.180 -87.540 ;
        RECT -190.440 -87.550 -189.600 -87.490 ;
        RECT -180.520 -87.540 -179.680 -87.490 ;
        RECT -191.820 -90.640 -188.220 -89.035 ;
        RECT -186.860 -89.145 -183.260 -87.540 ;
        RECT -181.900 -90.640 -178.300 -89.035 ;
        RECT -176.940 -89.145 -173.340 -87.540 ;
        RECT -170.600 -87.550 -169.760 -87.490 ;
        RECT -160.680 -87.540 -159.840 -87.490 ;
        RECT -171.980 -90.640 -168.380 -89.035 ;
        RECT -167.020 -89.145 -163.420 -87.540 ;
        RECT -162.060 -90.640 -158.460 -89.035 ;
        RECT -157.100 -89.145 -153.500 -87.540 ;
        RECT -150.760 -87.550 -149.920 -87.490 ;
        RECT -140.840 -87.540 -140.000 -87.490 ;
        RECT -152.140 -90.640 -148.540 -89.035 ;
        RECT -147.180 -89.145 -143.580 -87.540 ;
        RECT -142.220 -90.640 -138.620 -89.035 ;
        RECT -137.260 -89.145 -133.660 -87.540 ;
        RECT -130.920 -87.550 -130.080 -87.490 ;
        RECT -121.000 -87.540 -120.160 -87.490 ;
        RECT -132.300 -90.640 -128.700 -89.035 ;
        RECT -127.340 -89.145 -123.740 -87.540 ;
        RECT -122.380 -90.640 -118.780 -89.035 ;
        RECT -117.420 -89.145 -113.820 -87.540 ;
        RECT -111.080 -87.550 -110.240 -87.490 ;
        RECT -101.160 -87.540 -100.320 -87.490 ;
        RECT -112.460 -90.640 -108.860 -89.035 ;
        RECT -107.500 -89.145 -103.900 -87.540 ;
        RECT -102.540 -90.640 -98.940 -89.035 ;
        RECT -97.580 -89.145 -93.980 -87.540 ;
        RECT -91.240 -87.550 -90.400 -87.490 ;
        RECT -81.320 -87.540 -80.480 -87.490 ;
        RECT -92.620 -90.640 -89.020 -89.035 ;
        RECT -87.660 -89.145 -84.060 -87.540 ;
        RECT -82.700 -90.640 -79.100 -89.035 ;
        RECT -77.740 -89.145 -74.140 -87.540 ;
        RECT -71.400 -87.550 -70.560 -87.490 ;
        RECT -61.480 -87.540 -60.640 -87.490 ;
        RECT -72.780 -90.640 -69.180 -89.035 ;
        RECT -67.820 -89.145 -64.220 -87.540 ;
        RECT -62.860 -90.640 -59.260 -89.035 ;
        RECT -57.900 -89.145 -54.300 -87.540 ;
        RECT -51.560 -87.550 -50.720 -87.490 ;
        RECT -41.640 -87.540 -40.800 -87.490 ;
        RECT -52.940 -90.640 -49.340 -89.035 ;
        RECT -47.980 -89.145 -44.380 -87.540 ;
        RECT -43.020 -90.640 -39.420 -89.035 ;
        RECT -38.060 -89.145 -34.460 -87.540 ;
        RECT -31.720 -87.550 -30.880 -87.490 ;
        RECT -21.800 -87.540 -20.960 -87.490 ;
        RECT -33.100 -90.640 -29.500 -89.035 ;
        RECT -28.140 -89.145 -24.540 -87.540 ;
        RECT -23.180 -90.640 -19.580 -89.035 ;
        RECT -18.220 -89.145 -14.620 -87.540 ;
        RECT -11.880 -87.550 -11.040 -87.490 ;
        RECT -1.960 -87.540 -1.120 -87.490 ;
        RECT -13.260 -90.640 -9.660 -89.035 ;
        RECT -8.300 -89.145 -4.700 -87.540 ;
        RECT -3.340 -90.640 0.260 -89.035 ;
        RECT 1.620 -89.145 5.220 -87.540 ;
        RECT 7.960 -87.550 8.800 -87.490 ;
        RECT 17.880 -87.540 18.720 -87.490 ;
        RECT 27.800 -87.540 28.640 -87.490 ;
        RECT 6.580 -90.640 10.180 -89.035 ;
        RECT 11.540 -89.145 15.140 -87.540 ;
        RECT 16.500 -90.640 20.100 -89.035 ;
        RECT 21.460 -89.145 25.060 -87.540 ;
        RECT 26.420 -90.640 28.640 -89.035 ;
        RECT -286.145 -92.450 -282.375 -90.690 ;
        RECT -276.225 -92.450 -272.455 -90.690 ;
        RECT -266.305 -92.450 -262.535 -90.690 ;
        RECT -256.385 -92.450 -252.615 -90.690 ;
        RECT -246.465 -92.450 -242.695 -90.690 ;
        RECT -236.545 -92.450 -232.775 -90.690 ;
        RECT -226.625 -92.450 -222.855 -90.690 ;
        RECT -216.705 -92.450 -212.935 -90.690 ;
        RECT -206.785 -92.450 -203.015 -90.690 ;
        RECT -196.865 -92.450 -193.095 -90.690 ;
        RECT -186.945 -92.450 -183.175 -90.690 ;
        RECT -177.025 -92.450 -173.255 -90.690 ;
        RECT -167.105 -92.450 -163.335 -90.690 ;
        RECT -157.185 -92.450 -153.415 -90.690 ;
        RECT -147.265 -92.450 -143.495 -90.690 ;
        RECT -137.345 -92.450 -133.575 -90.690 ;
        RECT -127.425 -92.450 -123.655 -90.690 ;
        RECT -117.505 -92.450 -113.735 -90.690 ;
        RECT -107.585 -92.450 -103.815 -90.690 ;
        RECT -97.665 -92.450 -93.895 -90.690 ;
        RECT -87.745 -92.450 -83.975 -90.690 ;
        RECT -77.825 -92.450 -74.055 -90.690 ;
        RECT -67.905 -92.450 -64.135 -90.690 ;
        RECT -57.985 -92.450 -54.215 -90.690 ;
        RECT -48.065 -92.450 -44.295 -90.690 ;
        RECT -38.145 -92.450 -34.375 -90.690 ;
        RECT -28.225 -92.450 -24.455 -90.690 ;
        RECT -18.305 -92.450 -14.535 -90.690 ;
        RECT -8.385 -92.450 -4.615 -90.690 ;
        RECT 1.535 -92.450 5.305 -90.690 ;
        RECT 11.455 -92.450 15.225 -90.690 ;
        RECT 21.375 -92.450 25.145 -90.690 ;
        RECT -280.935 -175.200 -277.165 -173.440 ;
        RECT -271.015 -175.200 -267.245 -173.440 ;
        RECT -261.095 -175.200 -257.325 -173.440 ;
        RECT -251.175 -175.200 -247.405 -173.440 ;
        RECT -241.255 -175.200 -237.485 -173.440 ;
        RECT -231.335 -175.200 -227.565 -173.440 ;
        RECT -221.415 -175.200 -217.645 -173.440 ;
        RECT -211.495 -175.200 -207.725 -173.440 ;
        RECT -201.575 -175.200 -197.805 -173.440 ;
        RECT -191.655 -175.200 -187.885 -173.440 ;
        RECT -181.735 -175.200 -177.965 -173.440 ;
        RECT -171.815 -175.200 -168.045 -173.440 ;
        RECT -161.895 -175.200 -158.125 -173.440 ;
        RECT -151.975 -175.200 -148.205 -173.440 ;
        RECT -142.055 -175.200 -138.285 -173.440 ;
        RECT -132.135 -175.200 -128.365 -173.440 ;
        RECT -122.215 -175.200 -118.445 -173.440 ;
        RECT -112.295 -175.200 -108.525 -173.440 ;
        RECT -102.375 -175.200 -98.605 -173.440 ;
        RECT -92.455 -175.200 -88.685 -173.440 ;
        RECT -82.535 -175.200 -78.765 -173.440 ;
        RECT -72.615 -175.200 -68.845 -173.440 ;
        RECT -62.695 -175.200 -58.925 -173.440 ;
        RECT -52.775 -175.200 -49.005 -173.440 ;
        RECT -42.855 -175.200 -39.085 -173.440 ;
        RECT -32.935 -175.200 -29.165 -173.440 ;
        RECT -23.015 -175.200 -19.245 -173.440 ;
        RECT -13.095 -175.200 -9.325 -173.440 ;
        RECT -3.175 -175.200 0.595 -173.440 ;
        RECT 6.745 -175.200 10.515 -173.440 ;
        RECT 16.665 -175.200 20.435 -173.440 ;
        RECT 26.585 -173.675 28.190 -173.440 ;
        RECT 26.585 -173.680 28.700 -173.675 ;
        RECT 26.585 -175.200 28.890 -173.680 ;
        RECT -279.470 -175.250 -278.630 -175.200 ;
        RECT -285.810 -176.855 -282.210 -175.250 ;
        RECT -280.850 -178.350 -277.250 -176.745 ;
        RECT -275.890 -176.855 -272.290 -175.250 ;
        RECT -269.550 -175.260 -268.710 -175.200 ;
        RECT -259.630 -175.250 -258.790 -175.200 ;
        RECT -270.930 -178.350 -267.330 -176.745 ;
        RECT -265.970 -176.855 -262.370 -175.250 ;
        RECT -261.010 -178.350 -257.410 -176.745 ;
        RECT -256.050 -176.855 -252.450 -175.250 ;
        RECT -249.710 -175.260 -248.870 -175.200 ;
        RECT -239.790 -175.250 -238.950 -175.200 ;
        RECT -251.090 -178.350 -247.490 -176.745 ;
        RECT -246.130 -176.855 -242.530 -175.250 ;
        RECT -241.170 -178.350 -237.570 -176.745 ;
        RECT -236.210 -176.855 -232.610 -175.250 ;
        RECT -229.870 -175.260 -229.030 -175.200 ;
        RECT -219.950 -175.250 -219.110 -175.200 ;
        RECT -231.250 -178.350 -227.650 -176.745 ;
        RECT -226.290 -176.855 -222.690 -175.250 ;
        RECT -221.330 -178.350 -217.730 -176.745 ;
        RECT -216.370 -176.855 -212.770 -175.250 ;
        RECT -210.030 -175.260 -209.190 -175.200 ;
        RECT -200.110 -175.250 -199.270 -175.200 ;
        RECT -211.410 -178.350 -207.810 -176.745 ;
        RECT -206.450 -176.855 -202.850 -175.250 ;
        RECT -201.490 -178.350 -197.890 -176.745 ;
        RECT -196.530 -176.855 -192.930 -175.250 ;
        RECT -190.190 -175.260 -189.350 -175.200 ;
        RECT -180.270 -175.250 -179.430 -175.200 ;
        RECT -191.570 -178.350 -187.970 -176.745 ;
        RECT -186.610 -176.855 -183.010 -175.250 ;
        RECT -181.650 -178.350 -178.050 -176.745 ;
        RECT -176.690 -176.855 -173.090 -175.250 ;
        RECT -170.350 -175.260 -169.510 -175.200 ;
        RECT -160.430 -175.250 -159.590 -175.200 ;
        RECT -171.730 -178.350 -168.130 -176.745 ;
        RECT -166.770 -176.855 -163.170 -175.250 ;
        RECT -161.810 -178.350 -158.210 -176.745 ;
        RECT -156.850 -176.855 -153.250 -175.250 ;
        RECT -150.510 -175.260 -149.670 -175.200 ;
        RECT -140.590 -175.250 -139.750 -175.200 ;
        RECT -151.890 -178.350 -148.290 -176.745 ;
        RECT -146.930 -176.855 -143.330 -175.250 ;
        RECT -141.970 -178.350 -138.370 -176.745 ;
        RECT -137.010 -176.855 -133.410 -175.250 ;
        RECT -130.670 -175.260 -129.830 -175.200 ;
        RECT -120.750 -175.250 -119.910 -175.200 ;
        RECT -132.050 -178.350 -128.450 -176.745 ;
        RECT -127.090 -176.855 -123.490 -175.250 ;
        RECT -122.130 -178.350 -118.530 -176.745 ;
        RECT -117.170 -176.855 -113.570 -175.250 ;
        RECT -110.830 -175.260 -109.990 -175.200 ;
        RECT -100.910 -175.250 -100.070 -175.200 ;
        RECT -112.210 -178.350 -108.610 -176.745 ;
        RECT -107.250 -176.855 -103.650 -175.250 ;
        RECT -102.290 -178.350 -98.690 -176.745 ;
        RECT -97.330 -176.855 -93.730 -175.250 ;
        RECT -90.990 -175.260 -90.150 -175.200 ;
        RECT -81.070 -175.250 -80.230 -175.200 ;
        RECT -92.370 -178.350 -88.770 -176.745 ;
        RECT -87.410 -176.855 -83.810 -175.250 ;
        RECT -82.450 -178.350 -78.850 -176.745 ;
        RECT -77.490 -176.855 -73.890 -175.250 ;
        RECT -71.150 -175.260 -70.310 -175.200 ;
        RECT -61.230 -175.250 -60.390 -175.200 ;
        RECT -72.530 -178.350 -68.930 -176.745 ;
        RECT -67.570 -176.855 -63.970 -175.250 ;
        RECT -62.610 -178.350 -59.010 -176.745 ;
        RECT -57.650 -176.855 -54.050 -175.250 ;
        RECT -51.310 -175.260 -50.470 -175.200 ;
        RECT -41.390 -175.250 -40.550 -175.200 ;
        RECT -52.690 -178.350 -49.090 -176.745 ;
        RECT -47.730 -176.855 -44.130 -175.250 ;
        RECT -42.770 -178.350 -39.170 -176.745 ;
        RECT -37.810 -176.855 -34.210 -175.250 ;
        RECT -31.470 -175.260 -30.630 -175.200 ;
        RECT -21.550 -175.250 -20.710 -175.200 ;
        RECT -32.850 -178.350 -29.250 -176.745 ;
        RECT -27.890 -176.855 -24.290 -175.250 ;
        RECT -22.930 -178.350 -19.330 -176.745 ;
        RECT -17.970 -176.855 -14.370 -175.250 ;
        RECT -11.630 -175.260 -10.790 -175.200 ;
        RECT -1.710 -175.250 -0.870 -175.200 ;
        RECT -13.010 -178.350 -9.410 -176.745 ;
        RECT -8.050 -176.855 -4.450 -175.250 ;
        RECT -3.090 -178.350 0.510 -176.745 ;
        RECT 1.870 -176.855 5.470 -175.250 ;
        RECT 8.210 -175.260 9.050 -175.200 ;
        RECT 18.130 -175.250 18.970 -175.200 ;
        RECT 28.050 -175.250 28.890 -175.200 ;
        RECT 6.830 -178.350 10.430 -176.745 ;
        RECT 11.790 -176.855 15.390 -175.250 ;
        RECT 16.750 -178.350 20.350 -176.745 ;
        RECT 21.710 -176.855 25.310 -175.250 ;
        RECT 26.670 -178.350 28.890 -176.745 ;
        RECT -285.895 -180.160 -282.125 -178.400 ;
        RECT -275.975 -180.160 -272.205 -178.400 ;
        RECT -266.055 -180.160 -262.285 -178.400 ;
        RECT -256.135 -180.160 -252.365 -178.400 ;
        RECT -246.215 -180.160 -242.445 -178.400 ;
        RECT -236.295 -180.160 -232.525 -178.400 ;
        RECT -226.375 -180.160 -222.605 -178.400 ;
        RECT -216.455 -180.160 -212.685 -178.400 ;
        RECT -206.535 -180.160 -202.765 -178.400 ;
        RECT -196.615 -180.160 -192.845 -178.400 ;
        RECT -186.695 -180.160 -182.925 -178.400 ;
        RECT -176.775 -180.160 -173.005 -178.400 ;
        RECT -166.855 -180.160 -163.085 -178.400 ;
        RECT -156.935 -180.160 -153.165 -178.400 ;
        RECT -147.015 -180.160 -143.245 -178.400 ;
        RECT -137.095 -180.160 -133.325 -178.400 ;
        RECT -127.175 -180.160 -123.405 -178.400 ;
        RECT -117.255 -180.160 -113.485 -178.400 ;
        RECT -107.335 -180.160 -103.565 -178.400 ;
        RECT -97.415 -180.160 -93.645 -178.400 ;
        RECT -87.495 -180.160 -83.725 -178.400 ;
        RECT -77.575 -180.160 -73.805 -178.400 ;
        RECT -67.655 -180.160 -63.885 -178.400 ;
        RECT -57.735 -180.160 -53.965 -178.400 ;
        RECT -47.815 -180.160 -44.045 -178.400 ;
        RECT -37.895 -180.160 -34.125 -178.400 ;
        RECT -27.975 -180.160 -24.205 -178.400 ;
        RECT -18.055 -180.160 -14.285 -178.400 ;
        RECT -8.135 -180.160 -4.365 -178.400 ;
        RECT 1.785 -180.160 5.555 -178.400 ;
        RECT 11.705 -180.160 15.475 -178.400 ;
        RECT 21.625 -180.160 25.395 -178.400 ;
      LAYER li1 ;
        RECT -281.865 94.990 -281.695 95.140 ;
        RECT -280.925 94.990 -280.755 95.140 ;
        RECT -281.865 94.820 -280.755 94.990 ;
        RECT -281.865 94.615 -281.695 94.820 ;
        RECT -282.625 94.285 -281.695 94.615 ;
        RECT -281.865 93.760 -281.695 94.285 ;
        RECT -281.455 93.655 -281.165 94.820 ;
        RECT -280.925 94.615 -280.755 94.820 ;
        RECT -271.945 94.990 -271.775 95.140 ;
        RECT -271.005 94.990 -270.835 95.140 ;
        RECT -271.945 94.820 -270.835 94.990 ;
        RECT -271.945 94.615 -271.775 94.820 ;
        RECT -280.925 94.285 -279.995 94.615 ;
        RECT -272.705 94.285 -271.775 94.615 ;
        RECT -280.925 93.760 -280.755 94.285 ;
        RECT -271.945 93.760 -271.775 94.285 ;
        RECT -271.535 93.655 -271.245 94.820 ;
        RECT -271.005 94.615 -270.835 94.820 ;
        RECT -262.025 94.990 -261.855 95.140 ;
        RECT -261.085 94.990 -260.915 95.140 ;
        RECT -262.025 94.820 -260.915 94.990 ;
        RECT -262.025 94.615 -261.855 94.820 ;
        RECT -271.005 94.285 -270.075 94.615 ;
        RECT -262.785 94.285 -261.855 94.615 ;
        RECT -271.005 93.760 -270.835 94.285 ;
        RECT -262.025 93.760 -261.855 94.285 ;
        RECT -261.615 93.655 -261.325 94.820 ;
        RECT -261.085 94.615 -260.915 94.820 ;
        RECT -252.105 94.990 -251.935 95.140 ;
        RECT -251.165 94.990 -250.995 95.140 ;
        RECT -252.105 94.820 -250.995 94.990 ;
        RECT -252.105 94.615 -251.935 94.820 ;
        RECT -261.085 94.285 -260.155 94.615 ;
        RECT -252.865 94.285 -251.935 94.615 ;
        RECT -261.085 93.760 -260.915 94.285 ;
        RECT -252.105 93.760 -251.935 94.285 ;
        RECT -251.695 93.655 -251.405 94.820 ;
        RECT -251.165 94.615 -250.995 94.820 ;
        RECT -242.185 94.990 -242.015 95.140 ;
        RECT -241.245 94.990 -241.075 95.140 ;
        RECT -242.185 94.820 -241.075 94.990 ;
        RECT -242.185 94.615 -242.015 94.820 ;
        RECT -251.165 94.285 -250.235 94.615 ;
        RECT -242.945 94.285 -242.015 94.615 ;
        RECT -251.165 93.760 -250.995 94.285 ;
        RECT -242.185 93.760 -242.015 94.285 ;
        RECT -241.775 93.655 -241.485 94.820 ;
        RECT -241.245 94.615 -241.075 94.820 ;
        RECT -232.265 94.990 -232.095 95.140 ;
        RECT -231.325 94.990 -231.155 95.140 ;
        RECT -232.265 94.820 -231.155 94.990 ;
        RECT -232.265 94.615 -232.095 94.820 ;
        RECT -241.245 94.285 -240.315 94.615 ;
        RECT -233.025 94.285 -232.095 94.615 ;
        RECT -241.245 93.760 -241.075 94.285 ;
        RECT -232.265 93.760 -232.095 94.285 ;
        RECT -231.855 93.655 -231.565 94.820 ;
        RECT -231.325 94.615 -231.155 94.820 ;
        RECT -222.345 94.990 -222.175 95.140 ;
        RECT -221.405 94.990 -221.235 95.140 ;
        RECT -222.345 94.820 -221.235 94.990 ;
        RECT -222.345 94.615 -222.175 94.820 ;
        RECT -231.325 94.285 -230.395 94.615 ;
        RECT -223.105 94.285 -222.175 94.615 ;
        RECT -231.325 93.760 -231.155 94.285 ;
        RECT -222.345 93.760 -222.175 94.285 ;
        RECT -221.935 93.655 -221.645 94.820 ;
        RECT -221.405 94.615 -221.235 94.820 ;
        RECT -212.425 94.990 -212.255 95.140 ;
        RECT -211.485 94.990 -211.315 95.140 ;
        RECT -212.425 94.820 -211.315 94.990 ;
        RECT -212.425 94.615 -212.255 94.820 ;
        RECT -221.405 94.285 -220.475 94.615 ;
        RECT -213.185 94.285 -212.255 94.615 ;
        RECT -221.405 93.760 -221.235 94.285 ;
        RECT -212.425 93.760 -212.255 94.285 ;
        RECT -212.015 93.655 -211.725 94.820 ;
        RECT -211.485 94.615 -211.315 94.820 ;
        RECT -202.505 94.990 -202.335 95.140 ;
        RECT -201.565 94.990 -201.395 95.140 ;
        RECT -202.505 94.820 -201.395 94.990 ;
        RECT -202.505 94.615 -202.335 94.820 ;
        RECT -211.485 94.285 -210.555 94.615 ;
        RECT -203.265 94.285 -202.335 94.615 ;
        RECT -211.485 93.760 -211.315 94.285 ;
        RECT -202.505 93.760 -202.335 94.285 ;
        RECT -202.095 93.655 -201.805 94.820 ;
        RECT -201.565 94.615 -201.395 94.820 ;
        RECT -192.585 94.990 -192.415 95.140 ;
        RECT -191.645 94.990 -191.475 95.140 ;
        RECT -192.585 94.820 -191.475 94.990 ;
        RECT -192.585 94.615 -192.415 94.820 ;
        RECT -201.565 94.285 -200.635 94.615 ;
        RECT -193.345 94.285 -192.415 94.615 ;
        RECT -201.565 93.760 -201.395 94.285 ;
        RECT -192.585 93.760 -192.415 94.285 ;
        RECT -192.175 93.655 -191.885 94.820 ;
        RECT -191.645 94.615 -191.475 94.820 ;
        RECT -182.665 94.990 -182.495 95.140 ;
        RECT -181.725 94.990 -181.555 95.140 ;
        RECT -182.665 94.820 -181.555 94.990 ;
        RECT -182.665 94.615 -182.495 94.820 ;
        RECT -191.645 94.285 -190.715 94.615 ;
        RECT -183.425 94.285 -182.495 94.615 ;
        RECT -191.645 93.760 -191.475 94.285 ;
        RECT -182.665 93.760 -182.495 94.285 ;
        RECT -182.255 93.655 -181.965 94.820 ;
        RECT -181.725 94.615 -181.555 94.820 ;
        RECT -172.745 94.990 -172.575 95.140 ;
        RECT -171.805 94.990 -171.635 95.140 ;
        RECT -172.745 94.820 -171.635 94.990 ;
        RECT -172.745 94.615 -172.575 94.820 ;
        RECT -181.725 94.285 -180.795 94.615 ;
        RECT -173.505 94.285 -172.575 94.615 ;
        RECT -181.725 93.760 -181.555 94.285 ;
        RECT -172.745 93.760 -172.575 94.285 ;
        RECT -172.335 93.655 -172.045 94.820 ;
        RECT -171.805 94.615 -171.635 94.820 ;
        RECT -162.825 94.990 -162.655 95.140 ;
        RECT -161.885 94.990 -161.715 95.140 ;
        RECT -162.825 94.820 -161.715 94.990 ;
        RECT -162.825 94.615 -162.655 94.820 ;
        RECT -171.805 94.285 -170.875 94.615 ;
        RECT -163.585 94.285 -162.655 94.615 ;
        RECT -171.805 93.760 -171.635 94.285 ;
        RECT -162.825 93.760 -162.655 94.285 ;
        RECT -162.415 93.655 -162.125 94.820 ;
        RECT -161.885 94.615 -161.715 94.820 ;
        RECT -152.905 94.990 -152.735 95.140 ;
        RECT -151.965 94.990 -151.795 95.140 ;
        RECT -152.905 94.820 -151.795 94.990 ;
        RECT -152.905 94.615 -152.735 94.820 ;
        RECT -161.885 94.285 -160.955 94.615 ;
        RECT -153.665 94.285 -152.735 94.615 ;
        RECT -161.885 93.760 -161.715 94.285 ;
        RECT -152.905 93.760 -152.735 94.285 ;
        RECT -152.495 93.655 -152.205 94.820 ;
        RECT -151.965 94.615 -151.795 94.820 ;
        RECT -142.985 94.990 -142.815 95.140 ;
        RECT -142.045 94.990 -141.875 95.140 ;
        RECT -142.985 94.820 -141.875 94.990 ;
        RECT -142.985 94.615 -142.815 94.820 ;
        RECT -151.965 94.285 -151.035 94.615 ;
        RECT -143.745 94.285 -142.815 94.615 ;
        RECT -151.965 93.760 -151.795 94.285 ;
        RECT -142.985 93.760 -142.815 94.285 ;
        RECT -142.575 93.655 -142.285 94.820 ;
        RECT -142.045 94.615 -141.875 94.820 ;
        RECT -133.065 94.990 -132.895 95.140 ;
        RECT -132.125 94.990 -131.955 95.140 ;
        RECT -133.065 94.820 -131.955 94.990 ;
        RECT -133.065 94.615 -132.895 94.820 ;
        RECT -142.045 94.285 -141.115 94.615 ;
        RECT -133.825 94.285 -132.895 94.615 ;
        RECT -142.045 93.760 -141.875 94.285 ;
        RECT -133.065 93.760 -132.895 94.285 ;
        RECT -132.655 93.655 -132.365 94.820 ;
        RECT -132.125 94.615 -131.955 94.820 ;
        RECT -123.145 94.990 -122.975 95.140 ;
        RECT -122.205 94.990 -122.035 95.140 ;
        RECT -123.145 94.820 -122.035 94.990 ;
        RECT -123.145 94.615 -122.975 94.820 ;
        RECT -132.125 94.285 -131.195 94.615 ;
        RECT -123.905 94.285 -122.975 94.615 ;
        RECT -132.125 93.760 -131.955 94.285 ;
        RECT -123.145 93.760 -122.975 94.285 ;
        RECT -122.735 93.655 -122.445 94.820 ;
        RECT -122.205 94.615 -122.035 94.820 ;
        RECT -113.225 94.990 -113.055 95.140 ;
        RECT -112.285 94.990 -112.115 95.140 ;
        RECT -113.225 94.820 -112.115 94.990 ;
        RECT -113.225 94.615 -113.055 94.820 ;
        RECT -122.205 94.285 -121.275 94.615 ;
        RECT -113.985 94.285 -113.055 94.615 ;
        RECT -122.205 93.760 -122.035 94.285 ;
        RECT -113.225 93.760 -113.055 94.285 ;
        RECT -112.815 93.655 -112.525 94.820 ;
        RECT -112.285 94.615 -112.115 94.820 ;
        RECT -103.305 94.990 -103.135 95.140 ;
        RECT -102.365 94.990 -102.195 95.140 ;
        RECT -103.305 94.820 -102.195 94.990 ;
        RECT -103.305 94.615 -103.135 94.820 ;
        RECT -112.285 94.285 -111.355 94.615 ;
        RECT -104.065 94.285 -103.135 94.615 ;
        RECT -112.285 93.760 -112.115 94.285 ;
        RECT -103.305 93.760 -103.135 94.285 ;
        RECT -102.895 93.655 -102.605 94.820 ;
        RECT -102.365 94.615 -102.195 94.820 ;
        RECT -93.385 94.990 -93.215 95.140 ;
        RECT -92.445 94.990 -92.275 95.140 ;
        RECT -93.385 94.820 -92.275 94.990 ;
        RECT -93.385 94.615 -93.215 94.820 ;
        RECT -102.365 94.285 -101.435 94.615 ;
        RECT -94.145 94.285 -93.215 94.615 ;
        RECT -102.365 93.760 -102.195 94.285 ;
        RECT -93.385 93.760 -93.215 94.285 ;
        RECT -92.975 93.655 -92.685 94.820 ;
        RECT -92.445 94.615 -92.275 94.820 ;
        RECT -83.465 94.990 -83.295 95.140 ;
        RECT -82.525 94.990 -82.355 95.140 ;
        RECT -83.465 94.820 -82.355 94.990 ;
        RECT -83.465 94.615 -83.295 94.820 ;
        RECT -92.445 94.285 -91.515 94.615 ;
        RECT -84.225 94.285 -83.295 94.615 ;
        RECT -92.445 93.760 -92.275 94.285 ;
        RECT -83.465 93.760 -83.295 94.285 ;
        RECT -83.055 93.655 -82.765 94.820 ;
        RECT -82.525 94.615 -82.355 94.820 ;
        RECT -73.545 94.990 -73.375 95.140 ;
        RECT -72.605 94.990 -72.435 95.140 ;
        RECT -73.545 94.820 -72.435 94.990 ;
        RECT -73.545 94.615 -73.375 94.820 ;
        RECT -82.525 94.285 -81.595 94.615 ;
        RECT -74.305 94.285 -73.375 94.615 ;
        RECT -82.525 93.760 -82.355 94.285 ;
        RECT -73.545 93.760 -73.375 94.285 ;
        RECT -73.135 93.655 -72.845 94.820 ;
        RECT -72.605 94.615 -72.435 94.820 ;
        RECT -63.625 94.990 -63.455 95.140 ;
        RECT -62.685 94.990 -62.515 95.140 ;
        RECT -63.625 94.820 -62.515 94.990 ;
        RECT -63.625 94.615 -63.455 94.820 ;
        RECT -72.605 94.285 -71.675 94.615 ;
        RECT -64.385 94.285 -63.455 94.615 ;
        RECT -72.605 93.760 -72.435 94.285 ;
        RECT -63.625 93.760 -63.455 94.285 ;
        RECT -63.215 93.655 -62.925 94.820 ;
        RECT -62.685 94.615 -62.515 94.820 ;
        RECT -53.705 94.990 -53.535 95.140 ;
        RECT -52.765 94.990 -52.595 95.140 ;
        RECT -53.705 94.820 -52.595 94.990 ;
        RECT -53.705 94.615 -53.535 94.820 ;
        RECT -62.685 94.285 -61.755 94.615 ;
        RECT -54.465 94.285 -53.535 94.615 ;
        RECT -62.685 93.760 -62.515 94.285 ;
        RECT -53.705 93.760 -53.535 94.285 ;
        RECT -53.295 93.655 -53.005 94.820 ;
        RECT -52.765 94.615 -52.595 94.820 ;
        RECT -43.785 94.990 -43.615 95.140 ;
        RECT -42.845 94.990 -42.675 95.140 ;
        RECT -43.785 94.820 -42.675 94.990 ;
        RECT -43.785 94.615 -43.615 94.820 ;
        RECT -52.765 94.285 -51.835 94.615 ;
        RECT -44.545 94.285 -43.615 94.615 ;
        RECT -52.765 93.760 -52.595 94.285 ;
        RECT -43.785 93.760 -43.615 94.285 ;
        RECT -43.375 93.655 -43.085 94.820 ;
        RECT -42.845 94.615 -42.675 94.820 ;
        RECT -33.865 94.990 -33.695 95.140 ;
        RECT -32.925 94.990 -32.755 95.140 ;
        RECT -33.865 94.820 -32.755 94.990 ;
        RECT -33.865 94.615 -33.695 94.820 ;
        RECT -42.845 94.285 -41.915 94.615 ;
        RECT -34.625 94.285 -33.695 94.615 ;
        RECT -42.845 93.760 -42.675 94.285 ;
        RECT -33.865 93.760 -33.695 94.285 ;
        RECT -33.455 93.655 -33.165 94.820 ;
        RECT -32.925 94.615 -32.755 94.820 ;
        RECT -23.945 94.990 -23.775 95.140 ;
        RECT -23.005 94.990 -22.835 95.140 ;
        RECT -23.945 94.820 -22.835 94.990 ;
        RECT -23.945 94.615 -23.775 94.820 ;
        RECT -32.925 94.285 -31.995 94.615 ;
        RECT -24.705 94.285 -23.775 94.615 ;
        RECT -32.925 93.760 -32.755 94.285 ;
        RECT -23.945 93.760 -23.775 94.285 ;
        RECT -23.535 93.655 -23.245 94.820 ;
        RECT -23.005 94.615 -22.835 94.820 ;
        RECT -14.025 94.990 -13.855 95.140 ;
        RECT -13.085 94.990 -12.915 95.140 ;
        RECT -14.025 94.820 -12.915 94.990 ;
        RECT -14.025 94.615 -13.855 94.820 ;
        RECT -23.005 94.285 -22.075 94.615 ;
        RECT -14.785 94.285 -13.855 94.615 ;
        RECT -23.005 93.760 -22.835 94.285 ;
        RECT -14.025 93.760 -13.855 94.285 ;
        RECT -13.615 93.655 -13.325 94.820 ;
        RECT -13.085 94.615 -12.915 94.820 ;
        RECT -4.105 94.990 -3.935 95.140 ;
        RECT -3.165 94.990 -2.995 95.140 ;
        RECT -4.105 94.820 -2.995 94.990 ;
        RECT -4.105 94.615 -3.935 94.820 ;
        RECT -13.085 94.285 -12.155 94.615 ;
        RECT -4.865 94.285 -3.935 94.615 ;
        RECT -13.085 93.760 -12.915 94.285 ;
        RECT -4.105 93.760 -3.935 94.285 ;
        RECT -3.695 93.655 -3.405 94.820 ;
        RECT -3.165 94.615 -2.995 94.820 ;
        RECT 5.815 94.990 5.985 95.140 ;
        RECT 6.755 94.990 6.925 95.140 ;
        RECT 5.815 94.820 6.925 94.990 ;
        RECT 5.815 94.615 5.985 94.820 ;
        RECT -3.165 94.285 -2.235 94.615 ;
        RECT 5.055 94.285 5.985 94.615 ;
        RECT -3.165 93.760 -2.995 94.285 ;
        RECT 5.815 93.760 5.985 94.285 ;
        RECT 6.225 93.655 6.515 94.820 ;
        RECT 6.755 94.615 6.925 94.820 ;
        RECT 15.735 94.990 15.905 95.140 ;
        RECT 16.675 94.990 16.845 95.140 ;
        RECT 15.735 94.820 16.845 94.990 ;
        RECT 15.735 94.615 15.905 94.820 ;
        RECT 6.755 94.285 7.685 94.615 ;
        RECT 14.975 94.285 15.905 94.615 ;
        RECT 6.755 93.760 6.925 94.285 ;
        RECT 15.735 93.760 15.905 94.285 ;
        RECT 16.145 93.655 16.435 94.820 ;
        RECT 16.675 94.615 16.845 94.820 ;
        RECT 25.655 94.990 25.825 95.140 ;
        RECT 25.655 94.820 26.440 94.990 ;
        RECT 25.655 94.615 25.825 94.820 ;
        RECT 16.675 94.285 17.605 94.615 ;
        RECT 24.895 94.285 25.825 94.615 ;
        RECT 16.675 93.760 16.845 94.285 ;
        RECT 25.655 93.760 25.825 94.285 ;
        RECT 26.065 93.655 26.355 94.820 ;
        RECT -287.880 93.245 -284.660 93.415 ;
        RECT -277.960 93.245 -274.740 93.415 ;
        RECT -268.040 93.245 -264.820 93.415 ;
        RECT -258.120 93.245 -254.900 93.415 ;
        RECT -248.200 93.245 -244.980 93.415 ;
        RECT -238.280 93.245 -235.060 93.415 ;
        RECT -228.360 93.245 -225.140 93.415 ;
        RECT -218.440 93.245 -215.220 93.415 ;
        RECT -208.520 93.245 -205.300 93.415 ;
        RECT -198.600 93.245 -195.380 93.415 ;
        RECT -188.680 93.245 -185.460 93.415 ;
        RECT -178.760 93.245 -175.540 93.415 ;
        RECT -168.840 93.245 -165.620 93.415 ;
        RECT -158.920 93.245 -155.700 93.415 ;
        RECT -149.000 93.245 -145.780 93.415 ;
        RECT -139.080 93.245 -135.860 93.415 ;
        RECT -129.160 93.245 -125.940 93.415 ;
        RECT -119.240 93.245 -116.020 93.415 ;
        RECT -109.320 93.245 -106.100 93.415 ;
        RECT -99.400 93.245 -96.180 93.415 ;
        RECT -89.480 93.245 -86.260 93.415 ;
        RECT -79.560 93.245 -76.340 93.415 ;
        RECT -69.640 93.245 -66.420 93.415 ;
        RECT -59.720 93.245 -56.500 93.415 ;
        RECT -49.800 93.245 -46.580 93.415 ;
        RECT -39.880 93.245 -36.660 93.415 ;
        RECT -29.960 93.245 -26.740 93.415 ;
        RECT -20.040 93.245 -16.820 93.415 ;
        RECT -10.120 93.245 -6.900 93.415 ;
        RECT -0.200 93.245 3.020 93.415 ;
        RECT 9.720 93.245 12.940 93.415 ;
        RECT 19.640 93.245 22.860 93.415 ;
        RECT -287.795 92.105 -287.535 93.245 ;
        RECT -286.865 92.105 -286.585 93.245 ;
        RECT -286.415 92.080 -286.125 93.245 ;
        RECT -285.955 92.105 -285.675 93.245 ;
        RECT -285.005 92.105 -284.745 93.245 ;
        RECT -277.875 92.105 -277.615 93.245 ;
        RECT -276.945 92.105 -276.665 93.245 ;
        RECT -276.495 92.080 -276.205 93.245 ;
        RECT -276.035 92.105 -275.755 93.245 ;
        RECT -275.085 92.105 -274.825 93.245 ;
        RECT -267.955 92.105 -267.695 93.245 ;
        RECT -267.025 92.105 -266.745 93.245 ;
        RECT -266.575 92.080 -266.285 93.245 ;
        RECT -266.115 92.105 -265.835 93.245 ;
        RECT -265.165 92.105 -264.905 93.245 ;
        RECT -258.035 92.105 -257.775 93.245 ;
        RECT -257.105 92.105 -256.825 93.245 ;
        RECT -256.655 92.080 -256.365 93.245 ;
        RECT -256.195 92.105 -255.915 93.245 ;
        RECT -255.245 92.105 -254.985 93.245 ;
        RECT -248.115 92.105 -247.855 93.245 ;
        RECT -247.185 92.105 -246.905 93.245 ;
        RECT -246.735 92.080 -246.445 93.245 ;
        RECT -246.275 92.105 -245.995 93.245 ;
        RECT -245.325 92.105 -245.065 93.245 ;
        RECT -238.195 92.105 -237.935 93.245 ;
        RECT -237.265 92.105 -236.985 93.245 ;
        RECT -236.815 92.080 -236.525 93.245 ;
        RECT -236.355 92.105 -236.075 93.245 ;
        RECT -235.405 92.105 -235.145 93.245 ;
        RECT -228.275 92.105 -228.015 93.245 ;
        RECT -227.345 92.105 -227.065 93.245 ;
        RECT -226.895 92.080 -226.605 93.245 ;
        RECT -226.435 92.105 -226.155 93.245 ;
        RECT -225.485 92.105 -225.225 93.245 ;
        RECT -218.355 92.105 -218.095 93.245 ;
        RECT -217.425 92.105 -217.145 93.245 ;
        RECT -216.975 92.080 -216.685 93.245 ;
        RECT -216.515 92.105 -216.235 93.245 ;
        RECT -215.565 92.105 -215.305 93.245 ;
        RECT -208.435 92.105 -208.175 93.245 ;
        RECT -207.505 92.105 -207.225 93.245 ;
        RECT -207.055 92.080 -206.765 93.245 ;
        RECT -206.595 92.105 -206.315 93.245 ;
        RECT -205.645 92.105 -205.385 93.245 ;
        RECT -198.515 92.105 -198.255 93.245 ;
        RECT -197.585 92.105 -197.305 93.245 ;
        RECT -197.135 92.080 -196.845 93.245 ;
        RECT -196.675 92.105 -196.395 93.245 ;
        RECT -195.725 92.105 -195.465 93.245 ;
        RECT -188.595 92.105 -188.335 93.245 ;
        RECT -187.665 92.105 -187.385 93.245 ;
        RECT -187.215 92.080 -186.925 93.245 ;
        RECT -186.755 92.105 -186.475 93.245 ;
        RECT -185.805 92.105 -185.545 93.245 ;
        RECT -178.675 92.105 -178.415 93.245 ;
        RECT -177.745 92.105 -177.465 93.245 ;
        RECT -177.295 92.080 -177.005 93.245 ;
        RECT -176.835 92.105 -176.555 93.245 ;
        RECT -175.885 92.105 -175.625 93.245 ;
        RECT -168.755 92.105 -168.495 93.245 ;
        RECT -167.825 92.105 -167.545 93.245 ;
        RECT -167.375 92.080 -167.085 93.245 ;
        RECT -166.915 92.105 -166.635 93.245 ;
        RECT -165.965 92.105 -165.705 93.245 ;
        RECT -158.835 92.105 -158.575 93.245 ;
        RECT -157.905 92.105 -157.625 93.245 ;
        RECT -157.455 92.080 -157.165 93.245 ;
        RECT -156.995 92.105 -156.715 93.245 ;
        RECT -156.045 92.105 -155.785 93.245 ;
        RECT -148.915 92.105 -148.655 93.245 ;
        RECT -147.985 92.105 -147.705 93.245 ;
        RECT -147.535 92.080 -147.245 93.245 ;
        RECT -147.075 92.105 -146.795 93.245 ;
        RECT -146.125 92.105 -145.865 93.245 ;
        RECT -138.995 92.105 -138.735 93.245 ;
        RECT -138.065 92.105 -137.785 93.245 ;
        RECT -137.615 92.080 -137.325 93.245 ;
        RECT -137.155 92.105 -136.875 93.245 ;
        RECT -136.205 92.105 -135.945 93.245 ;
        RECT -129.075 92.105 -128.815 93.245 ;
        RECT -128.145 92.105 -127.865 93.245 ;
        RECT -127.695 92.080 -127.405 93.245 ;
        RECT -127.235 92.105 -126.955 93.245 ;
        RECT -126.285 92.105 -126.025 93.245 ;
        RECT -119.155 92.105 -118.895 93.245 ;
        RECT -118.225 92.105 -117.945 93.245 ;
        RECT -117.775 92.080 -117.485 93.245 ;
        RECT -117.315 92.105 -117.035 93.245 ;
        RECT -116.365 92.105 -116.105 93.245 ;
        RECT -109.235 92.105 -108.975 93.245 ;
        RECT -108.305 92.105 -108.025 93.245 ;
        RECT -107.855 92.080 -107.565 93.245 ;
        RECT -107.395 92.105 -107.115 93.245 ;
        RECT -106.445 92.105 -106.185 93.245 ;
        RECT -99.315 92.105 -99.055 93.245 ;
        RECT -98.385 92.105 -98.105 93.245 ;
        RECT -97.935 92.080 -97.645 93.245 ;
        RECT -97.475 92.105 -97.195 93.245 ;
        RECT -96.525 92.105 -96.265 93.245 ;
        RECT -89.395 92.105 -89.135 93.245 ;
        RECT -88.465 92.105 -88.185 93.245 ;
        RECT -88.015 92.080 -87.725 93.245 ;
        RECT -87.555 92.105 -87.275 93.245 ;
        RECT -86.605 92.105 -86.345 93.245 ;
        RECT -79.475 92.105 -79.215 93.245 ;
        RECT -78.545 92.105 -78.265 93.245 ;
        RECT -78.095 92.080 -77.805 93.245 ;
        RECT -77.635 92.105 -77.355 93.245 ;
        RECT -76.685 92.105 -76.425 93.245 ;
        RECT -69.555 92.105 -69.295 93.245 ;
        RECT -68.625 92.105 -68.345 93.245 ;
        RECT -68.175 92.080 -67.885 93.245 ;
        RECT -67.715 92.105 -67.435 93.245 ;
        RECT -66.765 92.105 -66.505 93.245 ;
        RECT -59.635 92.105 -59.375 93.245 ;
        RECT -58.705 92.105 -58.425 93.245 ;
        RECT -58.255 92.080 -57.965 93.245 ;
        RECT -57.795 92.105 -57.515 93.245 ;
        RECT -56.845 92.105 -56.585 93.245 ;
        RECT -49.715 92.105 -49.455 93.245 ;
        RECT -48.785 92.105 -48.505 93.245 ;
        RECT -48.335 92.080 -48.045 93.245 ;
        RECT -47.875 92.105 -47.595 93.245 ;
        RECT -46.925 92.105 -46.665 93.245 ;
        RECT -39.795 92.105 -39.535 93.245 ;
        RECT -38.865 92.105 -38.585 93.245 ;
        RECT -38.415 92.080 -38.125 93.245 ;
        RECT -37.955 92.105 -37.675 93.245 ;
        RECT -37.005 92.105 -36.745 93.245 ;
        RECT -29.875 92.105 -29.615 93.245 ;
        RECT -28.945 92.105 -28.665 93.245 ;
        RECT -28.495 92.080 -28.205 93.245 ;
        RECT -28.035 92.105 -27.755 93.245 ;
        RECT -27.085 92.105 -26.825 93.245 ;
        RECT -19.955 92.105 -19.695 93.245 ;
        RECT -19.025 92.105 -18.745 93.245 ;
        RECT -18.575 92.080 -18.285 93.245 ;
        RECT -18.115 92.105 -17.835 93.245 ;
        RECT -17.165 92.105 -16.905 93.245 ;
        RECT -10.035 92.105 -9.775 93.245 ;
        RECT -9.105 92.105 -8.825 93.245 ;
        RECT -8.655 92.080 -8.365 93.245 ;
        RECT -8.195 92.105 -7.915 93.245 ;
        RECT -7.245 92.105 -6.985 93.245 ;
        RECT -0.115 92.105 0.145 93.245 ;
        RECT 0.815 92.105 1.095 93.245 ;
        RECT 1.265 92.080 1.555 93.245 ;
        RECT 1.725 92.105 2.005 93.245 ;
        RECT 2.675 92.105 2.935 93.245 ;
        RECT 9.805 92.105 10.065 93.245 ;
        RECT 10.735 92.105 11.015 93.245 ;
        RECT 11.185 92.080 11.475 93.245 ;
        RECT 11.645 92.105 11.925 93.245 ;
        RECT 12.595 92.105 12.855 93.245 ;
        RECT 19.725 92.105 19.985 93.245 ;
        RECT 20.655 92.105 20.935 93.245 ;
        RECT 21.105 92.080 21.395 93.245 ;
        RECT 21.565 92.105 21.845 93.245 ;
        RECT 22.515 92.105 22.775 93.245 ;
        RECT -282.835 90.695 -282.575 91.835 ;
        RECT -281.905 90.695 -281.625 91.835 ;
        RECT -281.455 90.695 -281.165 91.860 ;
        RECT -280.995 90.695 -280.715 91.835 ;
        RECT -280.045 90.695 -279.785 91.835 ;
        RECT -272.915 90.695 -272.655 91.835 ;
        RECT -271.985 90.695 -271.705 91.835 ;
        RECT -271.535 90.695 -271.245 91.860 ;
        RECT -271.075 90.695 -270.795 91.835 ;
        RECT -270.125 90.695 -269.865 91.835 ;
        RECT -262.995 90.695 -262.735 91.835 ;
        RECT -262.065 90.695 -261.785 91.835 ;
        RECT -261.615 90.695 -261.325 91.860 ;
        RECT -261.155 90.695 -260.875 91.835 ;
        RECT -260.205 90.695 -259.945 91.835 ;
        RECT -253.075 90.695 -252.815 91.835 ;
        RECT -252.145 90.695 -251.865 91.835 ;
        RECT -251.695 90.695 -251.405 91.860 ;
        RECT -251.235 90.695 -250.955 91.835 ;
        RECT -250.285 90.695 -250.025 91.835 ;
        RECT -243.155 90.695 -242.895 91.835 ;
        RECT -242.225 90.695 -241.945 91.835 ;
        RECT -241.775 90.695 -241.485 91.860 ;
        RECT -241.315 90.695 -241.035 91.835 ;
        RECT -240.365 90.695 -240.105 91.835 ;
        RECT -233.235 90.695 -232.975 91.835 ;
        RECT -232.305 90.695 -232.025 91.835 ;
        RECT -231.855 90.695 -231.565 91.860 ;
        RECT -231.395 90.695 -231.115 91.835 ;
        RECT -230.445 90.695 -230.185 91.835 ;
        RECT -223.315 90.695 -223.055 91.835 ;
        RECT -222.385 90.695 -222.105 91.835 ;
        RECT -221.935 90.695 -221.645 91.860 ;
        RECT -221.475 90.695 -221.195 91.835 ;
        RECT -220.525 90.695 -220.265 91.835 ;
        RECT -213.395 90.695 -213.135 91.835 ;
        RECT -212.465 90.695 -212.185 91.835 ;
        RECT -212.015 90.695 -211.725 91.860 ;
        RECT -211.555 90.695 -211.275 91.835 ;
        RECT -210.605 90.695 -210.345 91.835 ;
        RECT -203.475 90.695 -203.215 91.835 ;
        RECT -202.545 90.695 -202.265 91.835 ;
        RECT -202.095 90.695 -201.805 91.860 ;
        RECT -201.635 90.695 -201.355 91.835 ;
        RECT -200.685 90.695 -200.425 91.835 ;
        RECT -193.555 90.695 -193.295 91.835 ;
        RECT -192.625 90.695 -192.345 91.835 ;
        RECT -192.175 90.695 -191.885 91.860 ;
        RECT -191.715 90.695 -191.435 91.835 ;
        RECT -190.765 90.695 -190.505 91.835 ;
        RECT -183.635 90.695 -183.375 91.835 ;
        RECT -182.705 90.695 -182.425 91.835 ;
        RECT -182.255 90.695 -181.965 91.860 ;
        RECT -181.795 90.695 -181.515 91.835 ;
        RECT -180.845 90.695 -180.585 91.835 ;
        RECT -173.715 90.695 -173.455 91.835 ;
        RECT -172.785 90.695 -172.505 91.835 ;
        RECT -172.335 90.695 -172.045 91.860 ;
        RECT -171.875 90.695 -171.595 91.835 ;
        RECT -170.925 90.695 -170.665 91.835 ;
        RECT -163.795 90.695 -163.535 91.835 ;
        RECT -162.865 90.695 -162.585 91.835 ;
        RECT -162.415 90.695 -162.125 91.860 ;
        RECT -161.955 90.695 -161.675 91.835 ;
        RECT -161.005 90.695 -160.745 91.835 ;
        RECT -153.875 90.695 -153.615 91.835 ;
        RECT -152.945 90.695 -152.665 91.835 ;
        RECT -152.495 90.695 -152.205 91.860 ;
        RECT -152.035 90.695 -151.755 91.835 ;
        RECT -151.085 90.695 -150.825 91.835 ;
        RECT -143.955 90.695 -143.695 91.835 ;
        RECT -143.025 90.695 -142.745 91.835 ;
        RECT -142.575 90.695 -142.285 91.860 ;
        RECT -142.115 90.695 -141.835 91.835 ;
        RECT -141.165 90.695 -140.905 91.835 ;
        RECT -134.035 90.695 -133.775 91.835 ;
        RECT -133.105 90.695 -132.825 91.835 ;
        RECT -132.655 90.695 -132.365 91.860 ;
        RECT -132.195 90.695 -131.915 91.835 ;
        RECT -131.245 90.695 -130.985 91.835 ;
        RECT -124.115 90.695 -123.855 91.835 ;
        RECT -123.185 90.695 -122.905 91.835 ;
        RECT -122.735 90.695 -122.445 91.860 ;
        RECT -122.275 90.695 -121.995 91.835 ;
        RECT -121.325 90.695 -121.065 91.835 ;
        RECT -114.195 90.695 -113.935 91.835 ;
        RECT -113.265 90.695 -112.985 91.835 ;
        RECT -112.815 90.695 -112.525 91.860 ;
        RECT -112.355 90.695 -112.075 91.835 ;
        RECT -111.405 90.695 -111.145 91.835 ;
        RECT -104.275 90.695 -104.015 91.835 ;
        RECT -103.345 90.695 -103.065 91.835 ;
        RECT -102.895 90.695 -102.605 91.860 ;
        RECT -102.435 90.695 -102.155 91.835 ;
        RECT -101.485 90.695 -101.225 91.835 ;
        RECT -94.355 90.695 -94.095 91.835 ;
        RECT -93.425 90.695 -93.145 91.835 ;
        RECT -92.975 90.695 -92.685 91.860 ;
        RECT -92.515 90.695 -92.235 91.835 ;
        RECT -91.565 90.695 -91.305 91.835 ;
        RECT -84.435 90.695 -84.175 91.835 ;
        RECT -83.505 90.695 -83.225 91.835 ;
        RECT -83.055 90.695 -82.765 91.860 ;
        RECT -82.595 90.695 -82.315 91.835 ;
        RECT -81.645 90.695 -81.385 91.835 ;
        RECT -74.515 90.695 -74.255 91.835 ;
        RECT -73.585 90.695 -73.305 91.835 ;
        RECT -73.135 90.695 -72.845 91.860 ;
        RECT -72.675 90.695 -72.395 91.835 ;
        RECT -71.725 90.695 -71.465 91.835 ;
        RECT -64.595 90.695 -64.335 91.835 ;
        RECT -63.665 90.695 -63.385 91.835 ;
        RECT -63.215 90.695 -62.925 91.860 ;
        RECT -62.755 90.695 -62.475 91.835 ;
        RECT -61.805 90.695 -61.545 91.835 ;
        RECT -54.675 90.695 -54.415 91.835 ;
        RECT -53.745 90.695 -53.465 91.835 ;
        RECT -53.295 90.695 -53.005 91.860 ;
        RECT -52.835 90.695 -52.555 91.835 ;
        RECT -51.885 90.695 -51.625 91.835 ;
        RECT -44.755 90.695 -44.495 91.835 ;
        RECT -43.825 90.695 -43.545 91.835 ;
        RECT -43.375 90.695 -43.085 91.860 ;
        RECT -42.915 90.695 -42.635 91.835 ;
        RECT -41.965 90.695 -41.705 91.835 ;
        RECT -34.835 90.695 -34.575 91.835 ;
        RECT -33.905 90.695 -33.625 91.835 ;
        RECT -33.455 90.695 -33.165 91.860 ;
        RECT -32.995 90.695 -32.715 91.835 ;
        RECT -32.045 90.695 -31.785 91.835 ;
        RECT -24.915 90.695 -24.655 91.835 ;
        RECT -23.985 90.695 -23.705 91.835 ;
        RECT -23.535 90.695 -23.245 91.860 ;
        RECT -23.075 90.695 -22.795 91.835 ;
        RECT -22.125 90.695 -21.865 91.835 ;
        RECT -14.995 90.695 -14.735 91.835 ;
        RECT -14.065 90.695 -13.785 91.835 ;
        RECT -13.615 90.695 -13.325 91.860 ;
        RECT -13.155 90.695 -12.875 91.835 ;
        RECT -12.205 90.695 -11.945 91.835 ;
        RECT -5.075 90.695 -4.815 91.835 ;
        RECT -4.145 90.695 -3.865 91.835 ;
        RECT -3.695 90.695 -3.405 91.860 ;
        RECT -3.235 90.695 -2.955 91.835 ;
        RECT -2.285 90.695 -2.025 91.835 ;
        RECT 4.845 90.695 5.105 91.835 ;
        RECT 5.775 90.695 6.055 91.835 ;
        RECT 6.225 90.695 6.515 91.860 ;
        RECT 6.685 90.695 6.965 91.835 ;
        RECT 7.635 90.695 7.895 91.835 ;
        RECT 14.765 90.695 15.025 91.835 ;
        RECT 15.695 90.695 15.975 91.835 ;
        RECT 16.145 90.695 16.435 91.860 ;
        RECT 16.605 90.695 16.885 91.835 ;
        RECT 17.555 90.695 17.815 91.835 ;
        RECT 24.685 90.695 24.945 91.835 ;
        RECT 25.615 90.695 25.895 91.835 ;
        RECT 26.065 90.695 26.355 91.860 ;
        RECT -282.920 90.525 -279.700 90.695 ;
        RECT -273.000 90.525 -269.780 90.695 ;
        RECT -263.080 90.525 -259.860 90.695 ;
        RECT -253.160 90.525 -249.940 90.695 ;
        RECT -243.240 90.525 -240.020 90.695 ;
        RECT -233.320 90.525 -230.100 90.695 ;
        RECT -223.400 90.525 -220.180 90.695 ;
        RECT -213.480 90.525 -210.260 90.695 ;
        RECT -203.560 90.525 -200.340 90.695 ;
        RECT -193.640 90.525 -190.420 90.695 ;
        RECT -183.720 90.525 -180.500 90.695 ;
        RECT -173.800 90.525 -170.580 90.695 ;
        RECT -163.880 90.525 -160.660 90.695 ;
        RECT -153.960 90.525 -150.740 90.695 ;
        RECT -144.040 90.525 -140.820 90.695 ;
        RECT -134.120 90.525 -130.900 90.695 ;
        RECT -124.200 90.525 -120.980 90.695 ;
        RECT -114.280 90.525 -111.060 90.695 ;
        RECT -104.360 90.525 -101.140 90.695 ;
        RECT -94.440 90.525 -91.220 90.695 ;
        RECT -84.520 90.525 -81.300 90.695 ;
        RECT -74.600 90.525 -71.380 90.695 ;
        RECT -64.680 90.525 -61.460 90.695 ;
        RECT -54.760 90.525 -51.540 90.695 ;
        RECT -44.840 90.525 -41.620 90.695 ;
        RECT -34.920 90.525 -31.700 90.695 ;
        RECT -25.000 90.525 -21.780 90.695 ;
        RECT -15.080 90.525 -11.860 90.695 ;
        RECT -5.160 90.525 -1.940 90.695 ;
        RECT 4.760 90.525 7.980 90.695 ;
        RECT 14.680 90.525 17.900 90.695 ;
        RECT 24.600 90.525 26.440 90.695 ;
        RECT -286.825 90.110 -286.655 90.180 ;
        RECT -285.885 90.110 -285.715 90.180 ;
        RECT -286.825 89.940 -285.715 90.110 ;
        RECT -286.825 89.655 -286.655 89.940 ;
        RECT -287.585 89.325 -286.655 89.655 ;
        RECT -286.825 88.800 -286.655 89.325 ;
        RECT -286.415 88.775 -286.125 89.940 ;
        RECT -285.885 89.655 -285.715 89.940 ;
        RECT -276.905 90.110 -276.735 90.180 ;
        RECT -275.965 90.110 -275.795 90.180 ;
        RECT -276.905 89.940 -275.795 90.110 ;
        RECT -276.905 89.655 -276.735 89.940 ;
        RECT -285.885 89.325 -284.955 89.655 ;
        RECT -277.665 89.325 -276.735 89.655 ;
        RECT -285.885 88.800 -285.715 89.325 ;
        RECT -276.905 88.800 -276.735 89.325 ;
        RECT -276.495 88.775 -276.205 89.940 ;
        RECT -275.965 89.655 -275.795 89.940 ;
        RECT -266.985 90.110 -266.815 90.180 ;
        RECT -266.045 90.110 -265.875 90.180 ;
        RECT -266.985 89.940 -265.875 90.110 ;
        RECT -266.985 89.655 -266.815 89.940 ;
        RECT -275.965 89.325 -275.035 89.655 ;
        RECT -267.745 89.325 -266.815 89.655 ;
        RECT -275.965 88.800 -275.795 89.325 ;
        RECT -266.985 88.800 -266.815 89.325 ;
        RECT -266.575 88.775 -266.285 89.940 ;
        RECT -266.045 89.655 -265.875 89.940 ;
        RECT -257.065 90.110 -256.895 90.180 ;
        RECT -256.125 90.110 -255.955 90.180 ;
        RECT -257.065 89.940 -255.955 90.110 ;
        RECT -257.065 89.655 -256.895 89.940 ;
        RECT -266.045 89.325 -265.115 89.655 ;
        RECT -257.825 89.325 -256.895 89.655 ;
        RECT -266.045 88.800 -265.875 89.325 ;
        RECT -257.065 88.800 -256.895 89.325 ;
        RECT -256.655 88.775 -256.365 89.940 ;
        RECT -256.125 89.655 -255.955 89.940 ;
        RECT -247.145 90.110 -246.975 90.180 ;
        RECT -246.205 90.110 -246.035 90.180 ;
        RECT -247.145 89.940 -246.035 90.110 ;
        RECT -247.145 89.655 -246.975 89.940 ;
        RECT -256.125 89.325 -255.195 89.655 ;
        RECT -247.905 89.325 -246.975 89.655 ;
        RECT -256.125 88.800 -255.955 89.325 ;
        RECT -247.145 88.800 -246.975 89.325 ;
        RECT -246.735 88.775 -246.445 89.940 ;
        RECT -246.205 89.655 -246.035 89.940 ;
        RECT -237.225 90.110 -237.055 90.180 ;
        RECT -236.285 90.110 -236.115 90.180 ;
        RECT -237.225 89.940 -236.115 90.110 ;
        RECT -237.225 89.655 -237.055 89.940 ;
        RECT -246.205 89.325 -245.275 89.655 ;
        RECT -237.985 89.325 -237.055 89.655 ;
        RECT -246.205 88.800 -246.035 89.325 ;
        RECT -237.225 88.800 -237.055 89.325 ;
        RECT -236.815 88.775 -236.525 89.940 ;
        RECT -236.285 89.655 -236.115 89.940 ;
        RECT -227.305 90.110 -227.135 90.180 ;
        RECT -226.365 90.110 -226.195 90.180 ;
        RECT -227.305 89.940 -226.195 90.110 ;
        RECT -227.305 89.655 -227.135 89.940 ;
        RECT -236.285 89.325 -235.355 89.655 ;
        RECT -228.065 89.325 -227.135 89.655 ;
        RECT -236.285 88.800 -236.115 89.325 ;
        RECT -227.305 88.800 -227.135 89.325 ;
        RECT -226.895 88.775 -226.605 89.940 ;
        RECT -226.365 89.655 -226.195 89.940 ;
        RECT -217.385 90.110 -217.215 90.180 ;
        RECT -216.445 90.110 -216.275 90.180 ;
        RECT -217.385 89.940 -216.275 90.110 ;
        RECT -217.385 89.655 -217.215 89.940 ;
        RECT -226.365 89.325 -225.435 89.655 ;
        RECT -218.145 89.325 -217.215 89.655 ;
        RECT -226.365 88.800 -226.195 89.325 ;
        RECT -217.385 88.800 -217.215 89.325 ;
        RECT -216.975 88.775 -216.685 89.940 ;
        RECT -216.445 89.655 -216.275 89.940 ;
        RECT -207.465 90.110 -207.295 90.180 ;
        RECT -206.525 90.110 -206.355 90.180 ;
        RECT -207.465 89.940 -206.355 90.110 ;
        RECT -207.465 89.655 -207.295 89.940 ;
        RECT -216.445 89.325 -215.515 89.655 ;
        RECT -208.225 89.325 -207.295 89.655 ;
        RECT -216.445 88.800 -216.275 89.325 ;
        RECT -207.465 88.800 -207.295 89.325 ;
        RECT -207.055 88.775 -206.765 89.940 ;
        RECT -206.525 89.655 -206.355 89.940 ;
        RECT -197.545 90.110 -197.375 90.180 ;
        RECT -196.605 90.110 -196.435 90.180 ;
        RECT -197.545 89.940 -196.435 90.110 ;
        RECT -197.545 89.655 -197.375 89.940 ;
        RECT -206.525 89.325 -205.595 89.655 ;
        RECT -198.305 89.325 -197.375 89.655 ;
        RECT -206.525 88.800 -206.355 89.325 ;
        RECT -197.545 88.800 -197.375 89.325 ;
        RECT -197.135 88.775 -196.845 89.940 ;
        RECT -196.605 89.655 -196.435 89.940 ;
        RECT -187.625 90.110 -187.455 90.180 ;
        RECT -186.685 90.110 -186.515 90.180 ;
        RECT -187.625 89.940 -186.515 90.110 ;
        RECT -187.625 89.655 -187.455 89.940 ;
        RECT -196.605 89.325 -195.675 89.655 ;
        RECT -188.385 89.325 -187.455 89.655 ;
        RECT -196.605 88.800 -196.435 89.325 ;
        RECT -187.625 88.800 -187.455 89.325 ;
        RECT -187.215 88.775 -186.925 89.940 ;
        RECT -186.685 89.655 -186.515 89.940 ;
        RECT -177.705 90.110 -177.535 90.180 ;
        RECT -176.765 90.110 -176.595 90.180 ;
        RECT -177.705 89.940 -176.595 90.110 ;
        RECT -177.705 89.655 -177.535 89.940 ;
        RECT -186.685 89.325 -185.755 89.655 ;
        RECT -178.465 89.325 -177.535 89.655 ;
        RECT -186.685 88.800 -186.515 89.325 ;
        RECT -177.705 88.800 -177.535 89.325 ;
        RECT -177.295 88.775 -177.005 89.940 ;
        RECT -176.765 89.655 -176.595 89.940 ;
        RECT -167.785 90.110 -167.615 90.180 ;
        RECT -166.845 90.110 -166.675 90.180 ;
        RECT -167.785 89.940 -166.675 90.110 ;
        RECT -167.785 89.655 -167.615 89.940 ;
        RECT -176.765 89.325 -175.835 89.655 ;
        RECT -168.545 89.325 -167.615 89.655 ;
        RECT -176.765 88.800 -176.595 89.325 ;
        RECT -167.785 88.800 -167.615 89.325 ;
        RECT -167.375 88.775 -167.085 89.940 ;
        RECT -166.845 89.655 -166.675 89.940 ;
        RECT -157.865 90.110 -157.695 90.180 ;
        RECT -156.925 90.110 -156.755 90.180 ;
        RECT -157.865 89.940 -156.755 90.110 ;
        RECT -157.865 89.655 -157.695 89.940 ;
        RECT -166.845 89.325 -165.915 89.655 ;
        RECT -158.625 89.325 -157.695 89.655 ;
        RECT -166.845 88.800 -166.675 89.325 ;
        RECT -157.865 88.800 -157.695 89.325 ;
        RECT -157.455 88.775 -157.165 89.940 ;
        RECT -156.925 89.655 -156.755 89.940 ;
        RECT -147.945 90.110 -147.775 90.180 ;
        RECT -147.005 90.110 -146.835 90.180 ;
        RECT -147.945 89.940 -146.835 90.110 ;
        RECT -147.945 89.655 -147.775 89.940 ;
        RECT -156.925 89.325 -155.995 89.655 ;
        RECT -148.705 89.325 -147.775 89.655 ;
        RECT -156.925 88.800 -156.755 89.325 ;
        RECT -147.945 88.800 -147.775 89.325 ;
        RECT -147.535 88.775 -147.245 89.940 ;
        RECT -147.005 89.655 -146.835 89.940 ;
        RECT -138.025 90.110 -137.855 90.180 ;
        RECT -137.085 90.110 -136.915 90.180 ;
        RECT -138.025 89.940 -136.915 90.110 ;
        RECT -138.025 89.655 -137.855 89.940 ;
        RECT -147.005 89.325 -146.075 89.655 ;
        RECT -138.785 89.325 -137.855 89.655 ;
        RECT -147.005 88.800 -146.835 89.325 ;
        RECT -138.025 88.800 -137.855 89.325 ;
        RECT -137.615 88.775 -137.325 89.940 ;
        RECT -137.085 89.655 -136.915 89.940 ;
        RECT -128.105 90.110 -127.935 90.180 ;
        RECT -127.165 90.110 -126.995 90.180 ;
        RECT -128.105 89.940 -126.995 90.110 ;
        RECT -128.105 89.655 -127.935 89.940 ;
        RECT -137.085 89.325 -136.155 89.655 ;
        RECT -128.865 89.325 -127.935 89.655 ;
        RECT -137.085 88.800 -136.915 89.325 ;
        RECT -128.105 88.800 -127.935 89.325 ;
        RECT -127.695 88.775 -127.405 89.940 ;
        RECT -127.165 89.655 -126.995 89.940 ;
        RECT -118.185 90.110 -118.015 90.180 ;
        RECT -117.245 90.110 -117.075 90.180 ;
        RECT -118.185 89.940 -117.075 90.110 ;
        RECT -118.185 89.655 -118.015 89.940 ;
        RECT -127.165 89.325 -126.235 89.655 ;
        RECT -118.945 89.325 -118.015 89.655 ;
        RECT -127.165 88.800 -126.995 89.325 ;
        RECT -118.185 88.800 -118.015 89.325 ;
        RECT -117.775 88.775 -117.485 89.940 ;
        RECT -117.245 89.655 -117.075 89.940 ;
        RECT -108.265 90.110 -108.095 90.180 ;
        RECT -107.325 90.110 -107.155 90.180 ;
        RECT -108.265 89.940 -107.155 90.110 ;
        RECT -108.265 89.655 -108.095 89.940 ;
        RECT -117.245 89.325 -116.315 89.655 ;
        RECT -109.025 89.325 -108.095 89.655 ;
        RECT -117.245 88.800 -117.075 89.325 ;
        RECT -108.265 88.800 -108.095 89.325 ;
        RECT -107.855 88.775 -107.565 89.940 ;
        RECT -107.325 89.655 -107.155 89.940 ;
        RECT -98.345 90.110 -98.175 90.180 ;
        RECT -97.405 90.110 -97.235 90.180 ;
        RECT -98.345 89.940 -97.235 90.110 ;
        RECT -98.345 89.655 -98.175 89.940 ;
        RECT -107.325 89.325 -106.395 89.655 ;
        RECT -99.105 89.325 -98.175 89.655 ;
        RECT -107.325 88.800 -107.155 89.325 ;
        RECT -98.345 88.800 -98.175 89.325 ;
        RECT -97.935 88.775 -97.645 89.940 ;
        RECT -97.405 89.655 -97.235 89.940 ;
        RECT -88.425 90.110 -88.255 90.180 ;
        RECT -87.485 90.110 -87.315 90.180 ;
        RECT -88.425 89.940 -87.315 90.110 ;
        RECT -88.425 89.655 -88.255 89.940 ;
        RECT -97.405 89.325 -96.475 89.655 ;
        RECT -89.185 89.325 -88.255 89.655 ;
        RECT -97.405 88.800 -97.235 89.325 ;
        RECT -88.425 88.800 -88.255 89.325 ;
        RECT -88.015 88.775 -87.725 89.940 ;
        RECT -87.485 89.655 -87.315 89.940 ;
        RECT -78.505 90.110 -78.335 90.180 ;
        RECT -77.565 90.110 -77.395 90.180 ;
        RECT -78.505 89.940 -77.395 90.110 ;
        RECT -78.505 89.655 -78.335 89.940 ;
        RECT -87.485 89.325 -86.555 89.655 ;
        RECT -79.265 89.325 -78.335 89.655 ;
        RECT -87.485 88.800 -87.315 89.325 ;
        RECT -78.505 88.800 -78.335 89.325 ;
        RECT -78.095 88.775 -77.805 89.940 ;
        RECT -77.565 89.655 -77.395 89.940 ;
        RECT -68.585 90.110 -68.415 90.180 ;
        RECT -67.645 90.110 -67.475 90.180 ;
        RECT -68.585 89.940 -67.475 90.110 ;
        RECT -68.585 89.655 -68.415 89.940 ;
        RECT -77.565 89.325 -76.635 89.655 ;
        RECT -69.345 89.325 -68.415 89.655 ;
        RECT -77.565 88.800 -77.395 89.325 ;
        RECT -68.585 88.800 -68.415 89.325 ;
        RECT -68.175 88.775 -67.885 89.940 ;
        RECT -67.645 89.655 -67.475 89.940 ;
        RECT -58.665 90.110 -58.495 90.180 ;
        RECT -57.725 90.110 -57.555 90.180 ;
        RECT -58.665 89.940 -57.555 90.110 ;
        RECT -58.665 89.655 -58.495 89.940 ;
        RECT -67.645 89.325 -66.715 89.655 ;
        RECT -59.425 89.325 -58.495 89.655 ;
        RECT -67.645 88.800 -67.475 89.325 ;
        RECT -58.665 88.800 -58.495 89.325 ;
        RECT -58.255 88.775 -57.965 89.940 ;
        RECT -57.725 89.655 -57.555 89.940 ;
        RECT -48.745 90.110 -48.575 90.180 ;
        RECT -47.805 90.110 -47.635 90.180 ;
        RECT -48.745 89.940 -47.635 90.110 ;
        RECT -48.745 89.655 -48.575 89.940 ;
        RECT -57.725 89.325 -56.795 89.655 ;
        RECT -49.505 89.325 -48.575 89.655 ;
        RECT -57.725 88.800 -57.555 89.325 ;
        RECT -48.745 88.800 -48.575 89.325 ;
        RECT -48.335 88.775 -48.045 89.940 ;
        RECT -47.805 89.655 -47.635 89.940 ;
        RECT -38.825 90.110 -38.655 90.180 ;
        RECT -37.885 90.110 -37.715 90.180 ;
        RECT -38.825 89.940 -37.715 90.110 ;
        RECT -38.825 89.655 -38.655 89.940 ;
        RECT -47.805 89.325 -46.875 89.655 ;
        RECT -39.585 89.325 -38.655 89.655 ;
        RECT -47.805 88.800 -47.635 89.325 ;
        RECT -38.825 88.800 -38.655 89.325 ;
        RECT -38.415 88.775 -38.125 89.940 ;
        RECT -37.885 89.655 -37.715 89.940 ;
        RECT -28.905 90.110 -28.735 90.180 ;
        RECT -27.965 90.110 -27.795 90.180 ;
        RECT -28.905 89.940 -27.795 90.110 ;
        RECT -28.905 89.655 -28.735 89.940 ;
        RECT -37.885 89.325 -36.955 89.655 ;
        RECT -29.665 89.325 -28.735 89.655 ;
        RECT -37.885 88.800 -37.715 89.325 ;
        RECT -28.905 88.800 -28.735 89.325 ;
        RECT -28.495 88.775 -28.205 89.940 ;
        RECT -27.965 89.655 -27.795 89.940 ;
        RECT -18.985 90.110 -18.815 90.180 ;
        RECT -18.045 90.110 -17.875 90.180 ;
        RECT -18.985 89.940 -17.875 90.110 ;
        RECT -18.985 89.655 -18.815 89.940 ;
        RECT -27.965 89.325 -27.035 89.655 ;
        RECT -19.745 89.325 -18.815 89.655 ;
        RECT -27.965 88.800 -27.795 89.325 ;
        RECT -18.985 88.800 -18.815 89.325 ;
        RECT -18.575 88.775 -18.285 89.940 ;
        RECT -18.045 89.655 -17.875 89.940 ;
        RECT -9.065 90.110 -8.895 90.180 ;
        RECT -8.125 90.110 -7.955 90.180 ;
        RECT -9.065 89.940 -7.955 90.110 ;
        RECT -9.065 89.655 -8.895 89.940 ;
        RECT -18.045 89.325 -17.115 89.655 ;
        RECT -9.825 89.325 -8.895 89.655 ;
        RECT -18.045 88.800 -17.875 89.325 ;
        RECT -9.065 88.800 -8.895 89.325 ;
        RECT -8.655 88.775 -8.365 89.940 ;
        RECT -8.125 89.655 -7.955 89.940 ;
        RECT 0.855 90.110 1.025 90.180 ;
        RECT 1.795 90.110 1.965 90.180 ;
        RECT 0.855 89.940 1.965 90.110 ;
        RECT 0.855 89.655 1.025 89.940 ;
        RECT -8.125 89.325 -7.195 89.655 ;
        RECT 0.095 89.325 1.025 89.655 ;
        RECT -8.125 88.800 -7.955 89.325 ;
        RECT 0.855 88.800 1.025 89.325 ;
        RECT 1.265 88.775 1.555 89.940 ;
        RECT 1.795 89.655 1.965 89.940 ;
        RECT 10.775 90.110 10.945 90.180 ;
        RECT 11.715 90.110 11.885 90.180 ;
        RECT 10.775 89.940 11.885 90.110 ;
        RECT 10.775 89.655 10.945 89.940 ;
        RECT 1.795 89.325 2.725 89.655 ;
        RECT 10.015 89.325 10.945 89.655 ;
        RECT 1.795 88.800 1.965 89.325 ;
        RECT 10.775 88.800 10.945 89.325 ;
        RECT 11.185 88.775 11.475 89.940 ;
        RECT 11.715 89.655 11.885 89.940 ;
        RECT 20.695 90.110 20.865 90.180 ;
        RECT 21.635 90.110 21.805 90.180 ;
        RECT 20.695 89.940 21.805 90.110 ;
        RECT 20.695 89.655 20.865 89.940 ;
        RECT 11.715 89.325 12.645 89.655 ;
        RECT 19.935 89.325 20.865 89.655 ;
        RECT 11.715 88.800 11.885 89.325 ;
        RECT 20.695 88.800 20.865 89.325 ;
        RECT 21.105 88.775 21.395 89.940 ;
        RECT 21.635 89.655 21.805 89.940 ;
        RECT 21.635 89.325 22.565 89.655 ;
        RECT 21.635 88.800 21.805 89.325 ;
        RECT -281.615 7.280 -281.445 7.430 ;
        RECT -280.675 7.280 -280.505 7.430 ;
        RECT -281.615 7.110 -280.505 7.280 ;
        RECT -281.615 6.905 -281.445 7.110 ;
        RECT -282.375 6.575 -281.445 6.905 ;
        RECT -281.615 6.050 -281.445 6.575 ;
        RECT -281.205 5.945 -280.915 7.110 ;
        RECT -280.675 6.905 -280.505 7.110 ;
        RECT -271.695 7.280 -271.525 7.430 ;
        RECT -270.755 7.280 -270.585 7.430 ;
        RECT -271.695 7.110 -270.585 7.280 ;
        RECT -271.695 6.905 -271.525 7.110 ;
        RECT -280.675 6.575 -279.745 6.905 ;
        RECT -272.455 6.575 -271.525 6.905 ;
        RECT -280.675 6.050 -280.505 6.575 ;
        RECT -271.695 6.050 -271.525 6.575 ;
        RECT -271.285 5.945 -270.995 7.110 ;
        RECT -270.755 6.905 -270.585 7.110 ;
        RECT -261.775 7.280 -261.605 7.430 ;
        RECT -260.835 7.280 -260.665 7.430 ;
        RECT -261.775 7.110 -260.665 7.280 ;
        RECT -261.775 6.905 -261.605 7.110 ;
        RECT -270.755 6.575 -269.825 6.905 ;
        RECT -262.535 6.575 -261.605 6.905 ;
        RECT -270.755 6.050 -270.585 6.575 ;
        RECT -261.775 6.050 -261.605 6.575 ;
        RECT -261.365 5.945 -261.075 7.110 ;
        RECT -260.835 6.905 -260.665 7.110 ;
        RECT -251.855 7.280 -251.685 7.430 ;
        RECT -250.915 7.280 -250.745 7.430 ;
        RECT -251.855 7.110 -250.745 7.280 ;
        RECT -251.855 6.905 -251.685 7.110 ;
        RECT -260.835 6.575 -259.905 6.905 ;
        RECT -252.615 6.575 -251.685 6.905 ;
        RECT -260.835 6.050 -260.665 6.575 ;
        RECT -251.855 6.050 -251.685 6.575 ;
        RECT -251.445 5.945 -251.155 7.110 ;
        RECT -250.915 6.905 -250.745 7.110 ;
        RECT -241.935 7.280 -241.765 7.430 ;
        RECT -240.995 7.280 -240.825 7.430 ;
        RECT -241.935 7.110 -240.825 7.280 ;
        RECT -241.935 6.905 -241.765 7.110 ;
        RECT -250.915 6.575 -249.985 6.905 ;
        RECT -242.695 6.575 -241.765 6.905 ;
        RECT -250.915 6.050 -250.745 6.575 ;
        RECT -241.935 6.050 -241.765 6.575 ;
        RECT -241.525 5.945 -241.235 7.110 ;
        RECT -240.995 6.905 -240.825 7.110 ;
        RECT -232.015 7.280 -231.845 7.430 ;
        RECT -231.075 7.280 -230.905 7.430 ;
        RECT -232.015 7.110 -230.905 7.280 ;
        RECT -232.015 6.905 -231.845 7.110 ;
        RECT -240.995 6.575 -240.065 6.905 ;
        RECT -232.775 6.575 -231.845 6.905 ;
        RECT -240.995 6.050 -240.825 6.575 ;
        RECT -232.015 6.050 -231.845 6.575 ;
        RECT -231.605 5.945 -231.315 7.110 ;
        RECT -231.075 6.905 -230.905 7.110 ;
        RECT -222.095 7.280 -221.925 7.430 ;
        RECT -221.155 7.280 -220.985 7.430 ;
        RECT -222.095 7.110 -220.985 7.280 ;
        RECT -222.095 6.905 -221.925 7.110 ;
        RECT -231.075 6.575 -230.145 6.905 ;
        RECT -222.855 6.575 -221.925 6.905 ;
        RECT -231.075 6.050 -230.905 6.575 ;
        RECT -222.095 6.050 -221.925 6.575 ;
        RECT -221.685 5.945 -221.395 7.110 ;
        RECT -221.155 6.905 -220.985 7.110 ;
        RECT -212.175 7.280 -212.005 7.430 ;
        RECT -211.235 7.280 -211.065 7.430 ;
        RECT -212.175 7.110 -211.065 7.280 ;
        RECT -212.175 6.905 -212.005 7.110 ;
        RECT -221.155 6.575 -220.225 6.905 ;
        RECT -212.935 6.575 -212.005 6.905 ;
        RECT -221.155 6.050 -220.985 6.575 ;
        RECT -212.175 6.050 -212.005 6.575 ;
        RECT -211.765 5.945 -211.475 7.110 ;
        RECT -211.235 6.905 -211.065 7.110 ;
        RECT -202.255 7.280 -202.085 7.430 ;
        RECT -201.315 7.280 -201.145 7.430 ;
        RECT -202.255 7.110 -201.145 7.280 ;
        RECT -202.255 6.905 -202.085 7.110 ;
        RECT -211.235 6.575 -210.305 6.905 ;
        RECT -203.015 6.575 -202.085 6.905 ;
        RECT -211.235 6.050 -211.065 6.575 ;
        RECT -202.255 6.050 -202.085 6.575 ;
        RECT -201.845 5.945 -201.555 7.110 ;
        RECT -201.315 6.905 -201.145 7.110 ;
        RECT -192.335 7.280 -192.165 7.430 ;
        RECT -191.395 7.280 -191.225 7.430 ;
        RECT -192.335 7.110 -191.225 7.280 ;
        RECT -192.335 6.905 -192.165 7.110 ;
        RECT -201.315 6.575 -200.385 6.905 ;
        RECT -193.095 6.575 -192.165 6.905 ;
        RECT -201.315 6.050 -201.145 6.575 ;
        RECT -192.335 6.050 -192.165 6.575 ;
        RECT -191.925 5.945 -191.635 7.110 ;
        RECT -191.395 6.905 -191.225 7.110 ;
        RECT -182.415 7.280 -182.245 7.430 ;
        RECT -181.475 7.280 -181.305 7.430 ;
        RECT -182.415 7.110 -181.305 7.280 ;
        RECT -182.415 6.905 -182.245 7.110 ;
        RECT -191.395 6.575 -190.465 6.905 ;
        RECT -183.175 6.575 -182.245 6.905 ;
        RECT -191.395 6.050 -191.225 6.575 ;
        RECT -182.415 6.050 -182.245 6.575 ;
        RECT -182.005 5.945 -181.715 7.110 ;
        RECT -181.475 6.905 -181.305 7.110 ;
        RECT -172.495 7.280 -172.325 7.430 ;
        RECT -171.555 7.280 -171.385 7.430 ;
        RECT -172.495 7.110 -171.385 7.280 ;
        RECT -172.495 6.905 -172.325 7.110 ;
        RECT -181.475 6.575 -180.545 6.905 ;
        RECT -173.255 6.575 -172.325 6.905 ;
        RECT -181.475 6.050 -181.305 6.575 ;
        RECT -172.495 6.050 -172.325 6.575 ;
        RECT -172.085 5.945 -171.795 7.110 ;
        RECT -171.555 6.905 -171.385 7.110 ;
        RECT -162.575 7.280 -162.405 7.430 ;
        RECT -161.635 7.280 -161.465 7.430 ;
        RECT -162.575 7.110 -161.465 7.280 ;
        RECT -162.575 6.905 -162.405 7.110 ;
        RECT -171.555 6.575 -170.625 6.905 ;
        RECT -163.335 6.575 -162.405 6.905 ;
        RECT -171.555 6.050 -171.385 6.575 ;
        RECT -162.575 6.050 -162.405 6.575 ;
        RECT -162.165 5.945 -161.875 7.110 ;
        RECT -161.635 6.905 -161.465 7.110 ;
        RECT -152.655 7.280 -152.485 7.430 ;
        RECT -151.715 7.280 -151.545 7.430 ;
        RECT -152.655 7.110 -151.545 7.280 ;
        RECT -152.655 6.905 -152.485 7.110 ;
        RECT -161.635 6.575 -160.705 6.905 ;
        RECT -153.415 6.575 -152.485 6.905 ;
        RECT -161.635 6.050 -161.465 6.575 ;
        RECT -152.655 6.050 -152.485 6.575 ;
        RECT -152.245 5.945 -151.955 7.110 ;
        RECT -151.715 6.905 -151.545 7.110 ;
        RECT -142.735 7.280 -142.565 7.430 ;
        RECT -141.795 7.280 -141.625 7.430 ;
        RECT -142.735 7.110 -141.625 7.280 ;
        RECT -142.735 6.905 -142.565 7.110 ;
        RECT -151.715 6.575 -150.785 6.905 ;
        RECT -143.495 6.575 -142.565 6.905 ;
        RECT -151.715 6.050 -151.545 6.575 ;
        RECT -142.735 6.050 -142.565 6.575 ;
        RECT -142.325 5.945 -142.035 7.110 ;
        RECT -141.795 6.905 -141.625 7.110 ;
        RECT -132.815 7.280 -132.645 7.430 ;
        RECT -131.875 7.280 -131.705 7.430 ;
        RECT -132.815 7.110 -131.705 7.280 ;
        RECT -132.815 6.905 -132.645 7.110 ;
        RECT -141.795 6.575 -140.865 6.905 ;
        RECT -133.575 6.575 -132.645 6.905 ;
        RECT -141.795 6.050 -141.625 6.575 ;
        RECT -132.815 6.050 -132.645 6.575 ;
        RECT -132.405 5.945 -132.115 7.110 ;
        RECT -131.875 6.905 -131.705 7.110 ;
        RECT -122.895 7.280 -122.725 7.430 ;
        RECT -121.955 7.280 -121.785 7.430 ;
        RECT -122.895 7.110 -121.785 7.280 ;
        RECT -122.895 6.905 -122.725 7.110 ;
        RECT -131.875 6.575 -130.945 6.905 ;
        RECT -123.655 6.575 -122.725 6.905 ;
        RECT -131.875 6.050 -131.705 6.575 ;
        RECT -122.895 6.050 -122.725 6.575 ;
        RECT -122.485 5.945 -122.195 7.110 ;
        RECT -121.955 6.905 -121.785 7.110 ;
        RECT -112.975 7.280 -112.805 7.430 ;
        RECT -112.035 7.280 -111.865 7.430 ;
        RECT -112.975 7.110 -111.865 7.280 ;
        RECT -112.975 6.905 -112.805 7.110 ;
        RECT -121.955 6.575 -121.025 6.905 ;
        RECT -113.735 6.575 -112.805 6.905 ;
        RECT -121.955 6.050 -121.785 6.575 ;
        RECT -112.975 6.050 -112.805 6.575 ;
        RECT -112.565 5.945 -112.275 7.110 ;
        RECT -112.035 6.905 -111.865 7.110 ;
        RECT -103.055 7.280 -102.885 7.430 ;
        RECT -102.115 7.280 -101.945 7.430 ;
        RECT -103.055 7.110 -101.945 7.280 ;
        RECT -103.055 6.905 -102.885 7.110 ;
        RECT -112.035 6.575 -111.105 6.905 ;
        RECT -103.815 6.575 -102.885 6.905 ;
        RECT -112.035 6.050 -111.865 6.575 ;
        RECT -103.055 6.050 -102.885 6.575 ;
        RECT -102.645 5.945 -102.355 7.110 ;
        RECT -102.115 6.905 -101.945 7.110 ;
        RECT -93.135 7.280 -92.965 7.430 ;
        RECT -92.195 7.280 -92.025 7.430 ;
        RECT -93.135 7.110 -92.025 7.280 ;
        RECT -93.135 6.905 -92.965 7.110 ;
        RECT -102.115 6.575 -101.185 6.905 ;
        RECT -93.895 6.575 -92.965 6.905 ;
        RECT -102.115 6.050 -101.945 6.575 ;
        RECT -93.135 6.050 -92.965 6.575 ;
        RECT -92.725 5.945 -92.435 7.110 ;
        RECT -92.195 6.905 -92.025 7.110 ;
        RECT -83.215 7.280 -83.045 7.430 ;
        RECT -82.275 7.280 -82.105 7.430 ;
        RECT -83.215 7.110 -82.105 7.280 ;
        RECT -83.215 6.905 -83.045 7.110 ;
        RECT -92.195 6.575 -91.265 6.905 ;
        RECT -83.975 6.575 -83.045 6.905 ;
        RECT -92.195 6.050 -92.025 6.575 ;
        RECT -83.215 6.050 -83.045 6.575 ;
        RECT -82.805 5.945 -82.515 7.110 ;
        RECT -82.275 6.905 -82.105 7.110 ;
        RECT -73.295 7.280 -73.125 7.430 ;
        RECT -72.355 7.280 -72.185 7.430 ;
        RECT -73.295 7.110 -72.185 7.280 ;
        RECT -73.295 6.905 -73.125 7.110 ;
        RECT -82.275 6.575 -81.345 6.905 ;
        RECT -74.055 6.575 -73.125 6.905 ;
        RECT -82.275 6.050 -82.105 6.575 ;
        RECT -73.295 6.050 -73.125 6.575 ;
        RECT -72.885 5.945 -72.595 7.110 ;
        RECT -72.355 6.905 -72.185 7.110 ;
        RECT -63.375 7.280 -63.205 7.430 ;
        RECT -62.435 7.280 -62.265 7.430 ;
        RECT -63.375 7.110 -62.265 7.280 ;
        RECT -63.375 6.905 -63.205 7.110 ;
        RECT -72.355 6.575 -71.425 6.905 ;
        RECT -64.135 6.575 -63.205 6.905 ;
        RECT -72.355 6.050 -72.185 6.575 ;
        RECT -63.375 6.050 -63.205 6.575 ;
        RECT -62.965 5.945 -62.675 7.110 ;
        RECT -62.435 6.905 -62.265 7.110 ;
        RECT -53.455 7.280 -53.285 7.430 ;
        RECT -52.515 7.280 -52.345 7.430 ;
        RECT -53.455 7.110 -52.345 7.280 ;
        RECT -53.455 6.905 -53.285 7.110 ;
        RECT -62.435 6.575 -61.505 6.905 ;
        RECT -54.215 6.575 -53.285 6.905 ;
        RECT -62.435 6.050 -62.265 6.575 ;
        RECT -53.455 6.050 -53.285 6.575 ;
        RECT -53.045 5.945 -52.755 7.110 ;
        RECT -52.515 6.905 -52.345 7.110 ;
        RECT -43.535 7.280 -43.365 7.430 ;
        RECT -42.595 7.280 -42.425 7.430 ;
        RECT -43.535 7.110 -42.425 7.280 ;
        RECT -43.535 6.905 -43.365 7.110 ;
        RECT -52.515 6.575 -51.585 6.905 ;
        RECT -44.295 6.575 -43.365 6.905 ;
        RECT -52.515 6.050 -52.345 6.575 ;
        RECT -43.535 6.050 -43.365 6.575 ;
        RECT -43.125 5.945 -42.835 7.110 ;
        RECT -42.595 6.905 -42.425 7.110 ;
        RECT -33.615 7.280 -33.445 7.430 ;
        RECT -32.675 7.280 -32.505 7.430 ;
        RECT -33.615 7.110 -32.505 7.280 ;
        RECT -33.615 6.905 -33.445 7.110 ;
        RECT -42.595 6.575 -41.665 6.905 ;
        RECT -34.375 6.575 -33.445 6.905 ;
        RECT -42.595 6.050 -42.425 6.575 ;
        RECT -33.615 6.050 -33.445 6.575 ;
        RECT -33.205 5.945 -32.915 7.110 ;
        RECT -32.675 6.905 -32.505 7.110 ;
        RECT -23.695 7.280 -23.525 7.430 ;
        RECT -22.755 7.280 -22.585 7.430 ;
        RECT -23.695 7.110 -22.585 7.280 ;
        RECT -23.695 6.905 -23.525 7.110 ;
        RECT -32.675 6.575 -31.745 6.905 ;
        RECT -24.455 6.575 -23.525 6.905 ;
        RECT -32.675 6.050 -32.505 6.575 ;
        RECT -23.695 6.050 -23.525 6.575 ;
        RECT -23.285 5.945 -22.995 7.110 ;
        RECT -22.755 6.905 -22.585 7.110 ;
        RECT -13.775 7.280 -13.605 7.430 ;
        RECT -12.835 7.280 -12.665 7.430 ;
        RECT -13.775 7.110 -12.665 7.280 ;
        RECT -13.775 6.905 -13.605 7.110 ;
        RECT -22.755 6.575 -21.825 6.905 ;
        RECT -14.535 6.575 -13.605 6.905 ;
        RECT -22.755 6.050 -22.585 6.575 ;
        RECT -13.775 6.050 -13.605 6.575 ;
        RECT -13.365 5.945 -13.075 7.110 ;
        RECT -12.835 6.905 -12.665 7.110 ;
        RECT -3.855 7.280 -3.685 7.430 ;
        RECT -2.915 7.280 -2.745 7.430 ;
        RECT -3.855 7.110 -2.745 7.280 ;
        RECT -3.855 6.905 -3.685 7.110 ;
        RECT -12.835 6.575 -11.905 6.905 ;
        RECT -4.615 6.575 -3.685 6.905 ;
        RECT -12.835 6.050 -12.665 6.575 ;
        RECT -3.855 6.050 -3.685 6.575 ;
        RECT -3.445 5.945 -3.155 7.110 ;
        RECT -2.915 6.905 -2.745 7.110 ;
        RECT 6.065 7.280 6.235 7.430 ;
        RECT 7.005 7.280 7.175 7.430 ;
        RECT 6.065 7.110 7.175 7.280 ;
        RECT 6.065 6.905 6.235 7.110 ;
        RECT -2.915 6.575 -1.985 6.905 ;
        RECT 5.305 6.575 6.235 6.905 ;
        RECT -2.915 6.050 -2.745 6.575 ;
        RECT 6.065 6.050 6.235 6.575 ;
        RECT 6.475 5.945 6.765 7.110 ;
        RECT 7.005 6.905 7.175 7.110 ;
        RECT 15.985 7.280 16.155 7.430 ;
        RECT 16.925 7.280 17.095 7.430 ;
        RECT 15.985 7.110 17.095 7.280 ;
        RECT 15.985 6.905 16.155 7.110 ;
        RECT 7.005 6.575 7.935 6.905 ;
        RECT 15.225 6.575 16.155 6.905 ;
        RECT 7.005 6.050 7.175 6.575 ;
        RECT 15.985 6.050 16.155 6.575 ;
        RECT 16.395 5.945 16.685 7.110 ;
        RECT 16.925 6.905 17.095 7.110 ;
        RECT 25.905 7.280 26.075 7.430 ;
        RECT 25.905 7.110 26.690 7.280 ;
        RECT 25.905 6.905 26.075 7.110 ;
        RECT 16.925 6.575 17.855 6.905 ;
        RECT 25.145 6.575 26.075 6.905 ;
        RECT 16.925 6.050 17.095 6.575 ;
        RECT 25.905 6.050 26.075 6.575 ;
        RECT 26.315 5.945 26.605 7.110 ;
        RECT -287.630 5.535 -284.410 5.705 ;
        RECT -277.710 5.535 -274.490 5.705 ;
        RECT -267.790 5.535 -264.570 5.705 ;
        RECT -257.870 5.535 -254.650 5.705 ;
        RECT -247.950 5.535 -244.730 5.705 ;
        RECT -238.030 5.535 -234.810 5.705 ;
        RECT -228.110 5.535 -224.890 5.705 ;
        RECT -218.190 5.535 -214.970 5.705 ;
        RECT -208.270 5.535 -205.050 5.705 ;
        RECT -198.350 5.535 -195.130 5.705 ;
        RECT -188.430 5.535 -185.210 5.705 ;
        RECT -178.510 5.535 -175.290 5.705 ;
        RECT -168.590 5.535 -165.370 5.705 ;
        RECT -158.670 5.535 -155.450 5.705 ;
        RECT -148.750 5.535 -145.530 5.705 ;
        RECT -138.830 5.535 -135.610 5.705 ;
        RECT -128.910 5.535 -125.690 5.705 ;
        RECT -118.990 5.535 -115.770 5.705 ;
        RECT -109.070 5.535 -105.850 5.705 ;
        RECT -99.150 5.535 -95.930 5.705 ;
        RECT -89.230 5.535 -86.010 5.705 ;
        RECT -79.310 5.535 -76.090 5.705 ;
        RECT -69.390 5.535 -66.170 5.705 ;
        RECT -59.470 5.535 -56.250 5.705 ;
        RECT -49.550 5.535 -46.330 5.705 ;
        RECT -39.630 5.535 -36.410 5.705 ;
        RECT -29.710 5.535 -26.490 5.705 ;
        RECT -19.790 5.535 -16.570 5.705 ;
        RECT -9.870 5.535 -6.650 5.705 ;
        RECT 0.050 5.535 3.270 5.705 ;
        RECT 9.970 5.535 13.190 5.705 ;
        RECT 19.890 5.535 23.110 5.705 ;
        RECT -287.545 4.395 -287.285 5.535 ;
        RECT -286.615 4.395 -286.335 5.535 ;
        RECT -286.165 4.370 -285.875 5.535 ;
        RECT -285.705 4.395 -285.425 5.535 ;
        RECT -284.755 4.395 -284.495 5.535 ;
        RECT -277.625 4.395 -277.365 5.535 ;
        RECT -276.695 4.395 -276.415 5.535 ;
        RECT -276.245 4.370 -275.955 5.535 ;
        RECT -275.785 4.395 -275.505 5.535 ;
        RECT -274.835 4.395 -274.575 5.535 ;
        RECT -267.705 4.395 -267.445 5.535 ;
        RECT -266.775 4.395 -266.495 5.535 ;
        RECT -266.325 4.370 -266.035 5.535 ;
        RECT -265.865 4.395 -265.585 5.535 ;
        RECT -264.915 4.395 -264.655 5.535 ;
        RECT -257.785 4.395 -257.525 5.535 ;
        RECT -256.855 4.395 -256.575 5.535 ;
        RECT -256.405 4.370 -256.115 5.535 ;
        RECT -255.945 4.395 -255.665 5.535 ;
        RECT -254.995 4.395 -254.735 5.535 ;
        RECT -247.865 4.395 -247.605 5.535 ;
        RECT -246.935 4.395 -246.655 5.535 ;
        RECT -246.485 4.370 -246.195 5.535 ;
        RECT -246.025 4.395 -245.745 5.535 ;
        RECT -245.075 4.395 -244.815 5.535 ;
        RECT -237.945 4.395 -237.685 5.535 ;
        RECT -237.015 4.395 -236.735 5.535 ;
        RECT -236.565 4.370 -236.275 5.535 ;
        RECT -236.105 4.395 -235.825 5.535 ;
        RECT -235.155 4.395 -234.895 5.535 ;
        RECT -228.025 4.395 -227.765 5.535 ;
        RECT -227.095 4.395 -226.815 5.535 ;
        RECT -226.645 4.370 -226.355 5.535 ;
        RECT -226.185 4.395 -225.905 5.535 ;
        RECT -225.235 4.395 -224.975 5.535 ;
        RECT -218.105 4.395 -217.845 5.535 ;
        RECT -217.175 4.395 -216.895 5.535 ;
        RECT -216.725 4.370 -216.435 5.535 ;
        RECT -216.265 4.395 -215.985 5.535 ;
        RECT -215.315 4.395 -215.055 5.535 ;
        RECT -208.185 4.395 -207.925 5.535 ;
        RECT -207.255 4.395 -206.975 5.535 ;
        RECT -206.805 4.370 -206.515 5.535 ;
        RECT -206.345 4.395 -206.065 5.535 ;
        RECT -205.395 4.395 -205.135 5.535 ;
        RECT -198.265 4.395 -198.005 5.535 ;
        RECT -197.335 4.395 -197.055 5.535 ;
        RECT -196.885 4.370 -196.595 5.535 ;
        RECT -196.425 4.395 -196.145 5.535 ;
        RECT -195.475 4.395 -195.215 5.535 ;
        RECT -188.345 4.395 -188.085 5.535 ;
        RECT -187.415 4.395 -187.135 5.535 ;
        RECT -186.965 4.370 -186.675 5.535 ;
        RECT -186.505 4.395 -186.225 5.535 ;
        RECT -185.555 4.395 -185.295 5.535 ;
        RECT -178.425 4.395 -178.165 5.535 ;
        RECT -177.495 4.395 -177.215 5.535 ;
        RECT -177.045 4.370 -176.755 5.535 ;
        RECT -176.585 4.395 -176.305 5.535 ;
        RECT -175.635 4.395 -175.375 5.535 ;
        RECT -168.505 4.395 -168.245 5.535 ;
        RECT -167.575 4.395 -167.295 5.535 ;
        RECT -167.125 4.370 -166.835 5.535 ;
        RECT -166.665 4.395 -166.385 5.535 ;
        RECT -165.715 4.395 -165.455 5.535 ;
        RECT -158.585 4.395 -158.325 5.535 ;
        RECT -157.655 4.395 -157.375 5.535 ;
        RECT -157.205 4.370 -156.915 5.535 ;
        RECT -156.745 4.395 -156.465 5.535 ;
        RECT -155.795 4.395 -155.535 5.535 ;
        RECT -148.665 4.395 -148.405 5.535 ;
        RECT -147.735 4.395 -147.455 5.535 ;
        RECT -147.285 4.370 -146.995 5.535 ;
        RECT -146.825 4.395 -146.545 5.535 ;
        RECT -145.875 4.395 -145.615 5.535 ;
        RECT -138.745 4.395 -138.485 5.535 ;
        RECT -137.815 4.395 -137.535 5.535 ;
        RECT -137.365 4.370 -137.075 5.535 ;
        RECT -136.905 4.395 -136.625 5.535 ;
        RECT -135.955 4.395 -135.695 5.535 ;
        RECT -128.825 4.395 -128.565 5.535 ;
        RECT -127.895 4.395 -127.615 5.535 ;
        RECT -127.445 4.370 -127.155 5.535 ;
        RECT -126.985 4.395 -126.705 5.535 ;
        RECT -126.035 4.395 -125.775 5.535 ;
        RECT -118.905 4.395 -118.645 5.535 ;
        RECT -117.975 4.395 -117.695 5.535 ;
        RECT -117.525 4.370 -117.235 5.535 ;
        RECT -117.065 4.395 -116.785 5.535 ;
        RECT -116.115 4.395 -115.855 5.535 ;
        RECT -108.985 4.395 -108.725 5.535 ;
        RECT -108.055 4.395 -107.775 5.535 ;
        RECT -107.605 4.370 -107.315 5.535 ;
        RECT -107.145 4.395 -106.865 5.535 ;
        RECT -106.195 4.395 -105.935 5.535 ;
        RECT -99.065 4.395 -98.805 5.535 ;
        RECT -98.135 4.395 -97.855 5.535 ;
        RECT -97.685 4.370 -97.395 5.535 ;
        RECT -97.225 4.395 -96.945 5.535 ;
        RECT -96.275 4.395 -96.015 5.535 ;
        RECT -89.145 4.395 -88.885 5.535 ;
        RECT -88.215 4.395 -87.935 5.535 ;
        RECT -87.765 4.370 -87.475 5.535 ;
        RECT -87.305 4.395 -87.025 5.535 ;
        RECT -86.355 4.395 -86.095 5.535 ;
        RECT -79.225 4.395 -78.965 5.535 ;
        RECT -78.295 4.395 -78.015 5.535 ;
        RECT -77.845 4.370 -77.555 5.535 ;
        RECT -77.385 4.395 -77.105 5.535 ;
        RECT -76.435 4.395 -76.175 5.535 ;
        RECT -69.305 4.395 -69.045 5.535 ;
        RECT -68.375 4.395 -68.095 5.535 ;
        RECT -67.925 4.370 -67.635 5.535 ;
        RECT -67.465 4.395 -67.185 5.535 ;
        RECT -66.515 4.395 -66.255 5.535 ;
        RECT -59.385 4.395 -59.125 5.535 ;
        RECT -58.455 4.395 -58.175 5.535 ;
        RECT -58.005 4.370 -57.715 5.535 ;
        RECT -57.545 4.395 -57.265 5.535 ;
        RECT -56.595 4.395 -56.335 5.535 ;
        RECT -49.465 4.395 -49.205 5.535 ;
        RECT -48.535 4.395 -48.255 5.535 ;
        RECT -48.085 4.370 -47.795 5.535 ;
        RECT -47.625 4.395 -47.345 5.535 ;
        RECT -46.675 4.395 -46.415 5.535 ;
        RECT -39.545 4.395 -39.285 5.535 ;
        RECT -38.615 4.395 -38.335 5.535 ;
        RECT -38.165 4.370 -37.875 5.535 ;
        RECT -37.705 4.395 -37.425 5.535 ;
        RECT -36.755 4.395 -36.495 5.535 ;
        RECT -29.625 4.395 -29.365 5.535 ;
        RECT -28.695 4.395 -28.415 5.535 ;
        RECT -28.245 4.370 -27.955 5.535 ;
        RECT -27.785 4.395 -27.505 5.535 ;
        RECT -26.835 4.395 -26.575 5.535 ;
        RECT -19.705 4.395 -19.445 5.535 ;
        RECT -18.775 4.395 -18.495 5.535 ;
        RECT -18.325 4.370 -18.035 5.535 ;
        RECT -17.865 4.395 -17.585 5.535 ;
        RECT -16.915 4.395 -16.655 5.535 ;
        RECT -9.785 4.395 -9.525 5.535 ;
        RECT -8.855 4.395 -8.575 5.535 ;
        RECT -8.405 4.370 -8.115 5.535 ;
        RECT -7.945 4.395 -7.665 5.535 ;
        RECT -6.995 4.395 -6.735 5.535 ;
        RECT 0.135 4.395 0.395 5.535 ;
        RECT 1.065 4.395 1.345 5.535 ;
        RECT 1.515 4.370 1.805 5.535 ;
        RECT 1.975 4.395 2.255 5.535 ;
        RECT 2.925 4.395 3.185 5.535 ;
        RECT 10.055 4.395 10.315 5.535 ;
        RECT 10.985 4.395 11.265 5.535 ;
        RECT 11.435 4.370 11.725 5.535 ;
        RECT 11.895 4.395 12.175 5.535 ;
        RECT 12.845 4.395 13.105 5.535 ;
        RECT 19.975 4.395 20.235 5.535 ;
        RECT 20.905 4.395 21.185 5.535 ;
        RECT 21.355 4.370 21.645 5.535 ;
        RECT 21.815 4.395 22.095 5.535 ;
        RECT 22.765 4.395 23.025 5.535 ;
        RECT -282.585 2.985 -282.325 4.125 ;
        RECT -281.655 2.985 -281.375 4.125 ;
        RECT -281.205 2.985 -280.915 4.150 ;
        RECT -280.745 2.985 -280.465 4.125 ;
        RECT -279.795 2.985 -279.535 4.125 ;
        RECT -272.665 2.985 -272.405 4.125 ;
        RECT -271.735 2.985 -271.455 4.125 ;
        RECT -271.285 2.985 -270.995 4.150 ;
        RECT -270.825 2.985 -270.545 4.125 ;
        RECT -269.875 2.985 -269.615 4.125 ;
        RECT -262.745 2.985 -262.485 4.125 ;
        RECT -261.815 2.985 -261.535 4.125 ;
        RECT -261.365 2.985 -261.075 4.150 ;
        RECT -260.905 2.985 -260.625 4.125 ;
        RECT -259.955 2.985 -259.695 4.125 ;
        RECT -252.825 2.985 -252.565 4.125 ;
        RECT -251.895 2.985 -251.615 4.125 ;
        RECT -251.445 2.985 -251.155 4.150 ;
        RECT -250.985 2.985 -250.705 4.125 ;
        RECT -250.035 2.985 -249.775 4.125 ;
        RECT -242.905 2.985 -242.645 4.125 ;
        RECT -241.975 2.985 -241.695 4.125 ;
        RECT -241.525 2.985 -241.235 4.150 ;
        RECT -241.065 2.985 -240.785 4.125 ;
        RECT -240.115 2.985 -239.855 4.125 ;
        RECT -232.985 2.985 -232.725 4.125 ;
        RECT -232.055 2.985 -231.775 4.125 ;
        RECT -231.605 2.985 -231.315 4.150 ;
        RECT -231.145 2.985 -230.865 4.125 ;
        RECT -230.195 2.985 -229.935 4.125 ;
        RECT -223.065 2.985 -222.805 4.125 ;
        RECT -222.135 2.985 -221.855 4.125 ;
        RECT -221.685 2.985 -221.395 4.150 ;
        RECT -221.225 2.985 -220.945 4.125 ;
        RECT -220.275 2.985 -220.015 4.125 ;
        RECT -213.145 2.985 -212.885 4.125 ;
        RECT -212.215 2.985 -211.935 4.125 ;
        RECT -211.765 2.985 -211.475 4.150 ;
        RECT -211.305 2.985 -211.025 4.125 ;
        RECT -210.355 2.985 -210.095 4.125 ;
        RECT -203.225 2.985 -202.965 4.125 ;
        RECT -202.295 2.985 -202.015 4.125 ;
        RECT -201.845 2.985 -201.555 4.150 ;
        RECT -201.385 2.985 -201.105 4.125 ;
        RECT -200.435 2.985 -200.175 4.125 ;
        RECT -193.305 2.985 -193.045 4.125 ;
        RECT -192.375 2.985 -192.095 4.125 ;
        RECT -191.925 2.985 -191.635 4.150 ;
        RECT -191.465 2.985 -191.185 4.125 ;
        RECT -190.515 2.985 -190.255 4.125 ;
        RECT -183.385 2.985 -183.125 4.125 ;
        RECT -182.455 2.985 -182.175 4.125 ;
        RECT -182.005 2.985 -181.715 4.150 ;
        RECT -181.545 2.985 -181.265 4.125 ;
        RECT -180.595 2.985 -180.335 4.125 ;
        RECT -173.465 2.985 -173.205 4.125 ;
        RECT -172.535 2.985 -172.255 4.125 ;
        RECT -172.085 2.985 -171.795 4.150 ;
        RECT -171.625 2.985 -171.345 4.125 ;
        RECT -170.675 2.985 -170.415 4.125 ;
        RECT -163.545 2.985 -163.285 4.125 ;
        RECT -162.615 2.985 -162.335 4.125 ;
        RECT -162.165 2.985 -161.875 4.150 ;
        RECT -161.705 2.985 -161.425 4.125 ;
        RECT -160.755 2.985 -160.495 4.125 ;
        RECT -153.625 2.985 -153.365 4.125 ;
        RECT -152.695 2.985 -152.415 4.125 ;
        RECT -152.245 2.985 -151.955 4.150 ;
        RECT -151.785 2.985 -151.505 4.125 ;
        RECT -150.835 2.985 -150.575 4.125 ;
        RECT -143.705 2.985 -143.445 4.125 ;
        RECT -142.775 2.985 -142.495 4.125 ;
        RECT -142.325 2.985 -142.035 4.150 ;
        RECT -141.865 2.985 -141.585 4.125 ;
        RECT -140.915 2.985 -140.655 4.125 ;
        RECT -133.785 2.985 -133.525 4.125 ;
        RECT -132.855 2.985 -132.575 4.125 ;
        RECT -132.405 2.985 -132.115 4.150 ;
        RECT -131.945 2.985 -131.665 4.125 ;
        RECT -130.995 2.985 -130.735 4.125 ;
        RECT -123.865 2.985 -123.605 4.125 ;
        RECT -122.935 2.985 -122.655 4.125 ;
        RECT -122.485 2.985 -122.195 4.150 ;
        RECT -122.025 2.985 -121.745 4.125 ;
        RECT -121.075 2.985 -120.815 4.125 ;
        RECT -113.945 2.985 -113.685 4.125 ;
        RECT -113.015 2.985 -112.735 4.125 ;
        RECT -112.565 2.985 -112.275 4.150 ;
        RECT -112.105 2.985 -111.825 4.125 ;
        RECT -111.155 2.985 -110.895 4.125 ;
        RECT -104.025 2.985 -103.765 4.125 ;
        RECT -103.095 2.985 -102.815 4.125 ;
        RECT -102.645 2.985 -102.355 4.150 ;
        RECT -102.185 2.985 -101.905 4.125 ;
        RECT -101.235 2.985 -100.975 4.125 ;
        RECT -94.105 2.985 -93.845 4.125 ;
        RECT -93.175 2.985 -92.895 4.125 ;
        RECT -92.725 2.985 -92.435 4.150 ;
        RECT -92.265 2.985 -91.985 4.125 ;
        RECT -91.315 2.985 -91.055 4.125 ;
        RECT -84.185 2.985 -83.925 4.125 ;
        RECT -83.255 2.985 -82.975 4.125 ;
        RECT -82.805 2.985 -82.515 4.150 ;
        RECT -82.345 2.985 -82.065 4.125 ;
        RECT -81.395 2.985 -81.135 4.125 ;
        RECT -74.265 2.985 -74.005 4.125 ;
        RECT -73.335 2.985 -73.055 4.125 ;
        RECT -72.885 2.985 -72.595 4.150 ;
        RECT -72.425 2.985 -72.145 4.125 ;
        RECT -71.475 2.985 -71.215 4.125 ;
        RECT -64.345 2.985 -64.085 4.125 ;
        RECT -63.415 2.985 -63.135 4.125 ;
        RECT -62.965 2.985 -62.675 4.150 ;
        RECT -62.505 2.985 -62.225 4.125 ;
        RECT -61.555 2.985 -61.295 4.125 ;
        RECT -54.425 2.985 -54.165 4.125 ;
        RECT -53.495 2.985 -53.215 4.125 ;
        RECT -53.045 2.985 -52.755 4.150 ;
        RECT -52.585 2.985 -52.305 4.125 ;
        RECT -51.635 2.985 -51.375 4.125 ;
        RECT -44.505 2.985 -44.245 4.125 ;
        RECT -43.575 2.985 -43.295 4.125 ;
        RECT -43.125 2.985 -42.835 4.150 ;
        RECT -42.665 2.985 -42.385 4.125 ;
        RECT -41.715 2.985 -41.455 4.125 ;
        RECT -34.585 2.985 -34.325 4.125 ;
        RECT -33.655 2.985 -33.375 4.125 ;
        RECT -33.205 2.985 -32.915 4.150 ;
        RECT -32.745 2.985 -32.465 4.125 ;
        RECT -31.795 2.985 -31.535 4.125 ;
        RECT -24.665 2.985 -24.405 4.125 ;
        RECT -23.735 2.985 -23.455 4.125 ;
        RECT -23.285 2.985 -22.995 4.150 ;
        RECT -22.825 2.985 -22.545 4.125 ;
        RECT -21.875 2.985 -21.615 4.125 ;
        RECT -14.745 2.985 -14.485 4.125 ;
        RECT -13.815 2.985 -13.535 4.125 ;
        RECT -13.365 2.985 -13.075 4.150 ;
        RECT -12.905 2.985 -12.625 4.125 ;
        RECT -11.955 2.985 -11.695 4.125 ;
        RECT -4.825 2.985 -4.565 4.125 ;
        RECT -3.895 2.985 -3.615 4.125 ;
        RECT -3.445 2.985 -3.155 4.150 ;
        RECT -2.985 2.985 -2.705 4.125 ;
        RECT -2.035 2.985 -1.775 4.125 ;
        RECT 5.095 2.985 5.355 4.125 ;
        RECT 6.025 2.985 6.305 4.125 ;
        RECT 6.475 2.985 6.765 4.150 ;
        RECT 6.935 2.985 7.215 4.125 ;
        RECT 7.885 2.985 8.145 4.125 ;
        RECT 15.015 2.985 15.275 4.125 ;
        RECT 15.945 2.985 16.225 4.125 ;
        RECT 16.395 2.985 16.685 4.150 ;
        RECT 16.855 2.985 17.135 4.125 ;
        RECT 17.805 2.985 18.065 4.125 ;
        RECT 24.935 2.985 25.195 4.125 ;
        RECT 25.865 2.985 26.145 4.125 ;
        RECT 26.315 2.985 26.605 4.150 ;
        RECT -282.670 2.815 -279.450 2.985 ;
        RECT -272.750 2.815 -269.530 2.985 ;
        RECT -262.830 2.815 -259.610 2.985 ;
        RECT -252.910 2.815 -249.690 2.985 ;
        RECT -242.990 2.815 -239.770 2.985 ;
        RECT -233.070 2.815 -229.850 2.985 ;
        RECT -223.150 2.815 -219.930 2.985 ;
        RECT -213.230 2.815 -210.010 2.985 ;
        RECT -203.310 2.815 -200.090 2.985 ;
        RECT -193.390 2.815 -190.170 2.985 ;
        RECT -183.470 2.815 -180.250 2.985 ;
        RECT -173.550 2.815 -170.330 2.985 ;
        RECT -163.630 2.815 -160.410 2.985 ;
        RECT -153.710 2.815 -150.490 2.985 ;
        RECT -143.790 2.815 -140.570 2.985 ;
        RECT -133.870 2.815 -130.650 2.985 ;
        RECT -123.950 2.815 -120.730 2.985 ;
        RECT -114.030 2.815 -110.810 2.985 ;
        RECT -104.110 2.815 -100.890 2.985 ;
        RECT -94.190 2.815 -90.970 2.985 ;
        RECT -84.270 2.815 -81.050 2.985 ;
        RECT -74.350 2.815 -71.130 2.985 ;
        RECT -64.430 2.815 -61.210 2.985 ;
        RECT -54.510 2.815 -51.290 2.985 ;
        RECT -44.590 2.815 -41.370 2.985 ;
        RECT -34.670 2.815 -31.450 2.985 ;
        RECT -24.750 2.815 -21.530 2.985 ;
        RECT -14.830 2.815 -11.610 2.985 ;
        RECT -4.910 2.815 -1.690 2.985 ;
        RECT 5.010 2.815 8.230 2.985 ;
        RECT 14.930 2.815 18.150 2.985 ;
        RECT 24.850 2.815 26.690 2.985 ;
        RECT -286.575 2.400 -286.405 2.470 ;
        RECT -285.635 2.400 -285.465 2.470 ;
        RECT -286.575 2.230 -285.465 2.400 ;
        RECT -286.575 1.945 -286.405 2.230 ;
        RECT -287.335 1.615 -286.405 1.945 ;
        RECT -286.575 1.090 -286.405 1.615 ;
        RECT -286.165 1.065 -285.875 2.230 ;
        RECT -285.635 1.945 -285.465 2.230 ;
        RECT -276.655 2.400 -276.485 2.470 ;
        RECT -275.715 2.400 -275.545 2.470 ;
        RECT -276.655 2.230 -275.545 2.400 ;
        RECT -276.655 1.945 -276.485 2.230 ;
        RECT -285.635 1.615 -284.705 1.945 ;
        RECT -277.415 1.615 -276.485 1.945 ;
        RECT -285.635 1.090 -285.465 1.615 ;
        RECT -276.655 1.090 -276.485 1.615 ;
        RECT -276.245 1.065 -275.955 2.230 ;
        RECT -275.715 1.945 -275.545 2.230 ;
        RECT -266.735 2.400 -266.565 2.470 ;
        RECT -265.795 2.400 -265.625 2.470 ;
        RECT -266.735 2.230 -265.625 2.400 ;
        RECT -266.735 1.945 -266.565 2.230 ;
        RECT -275.715 1.615 -274.785 1.945 ;
        RECT -267.495 1.615 -266.565 1.945 ;
        RECT -275.715 1.090 -275.545 1.615 ;
        RECT -266.735 1.090 -266.565 1.615 ;
        RECT -266.325 1.065 -266.035 2.230 ;
        RECT -265.795 1.945 -265.625 2.230 ;
        RECT -256.815 2.400 -256.645 2.470 ;
        RECT -255.875 2.400 -255.705 2.470 ;
        RECT -256.815 2.230 -255.705 2.400 ;
        RECT -256.815 1.945 -256.645 2.230 ;
        RECT -265.795 1.615 -264.865 1.945 ;
        RECT -257.575 1.615 -256.645 1.945 ;
        RECT -265.795 1.090 -265.625 1.615 ;
        RECT -256.815 1.090 -256.645 1.615 ;
        RECT -256.405 1.065 -256.115 2.230 ;
        RECT -255.875 1.945 -255.705 2.230 ;
        RECT -246.895 2.400 -246.725 2.470 ;
        RECT -245.955 2.400 -245.785 2.470 ;
        RECT -246.895 2.230 -245.785 2.400 ;
        RECT -246.895 1.945 -246.725 2.230 ;
        RECT -255.875 1.615 -254.945 1.945 ;
        RECT -247.655 1.615 -246.725 1.945 ;
        RECT -255.875 1.090 -255.705 1.615 ;
        RECT -246.895 1.090 -246.725 1.615 ;
        RECT -246.485 1.065 -246.195 2.230 ;
        RECT -245.955 1.945 -245.785 2.230 ;
        RECT -236.975 2.400 -236.805 2.470 ;
        RECT -236.035 2.400 -235.865 2.470 ;
        RECT -236.975 2.230 -235.865 2.400 ;
        RECT -236.975 1.945 -236.805 2.230 ;
        RECT -245.955 1.615 -245.025 1.945 ;
        RECT -237.735 1.615 -236.805 1.945 ;
        RECT -245.955 1.090 -245.785 1.615 ;
        RECT -236.975 1.090 -236.805 1.615 ;
        RECT -236.565 1.065 -236.275 2.230 ;
        RECT -236.035 1.945 -235.865 2.230 ;
        RECT -227.055 2.400 -226.885 2.470 ;
        RECT -226.115 2.400 -225.945 2.470 ;
        RECT -227.055 2.230 -225.945 2.400 ;
        RECT -227.055 1.945 -226.885 2.230 ;
        RECT -236.035 1.615 -235.105 1.945 ;
        RECT -227.815 1.615 -226.885 1.945 ;
        RECT -236.035 1.090 -235.865 1.615 ;
        RECT -227.055 1.090 -226.885 1.615 ;
        RECT -226.645 1.065 -226.355 2.230 ;
        RECT -226.115 1.945 -225.945 2.230 ;
        RECT -217.135 2.400 -216.965 2.470 ;
        RECT -216.195 2.400 -216.025 2.470 ;
        RECT -217.135 2.230 -216.025 2.400 ;
        RECT -217.135 1.945 -216.965 2.230 ;
        RECT -226.115 1.615 -225.185 1.945 ;
        RECT -217.895 1.615 -216.965 1.945 ;
        RECT -226.115 1.090 -225.945 1.615 ;
        RECT -217.135 1.090 -216.965 1.615 ;
        RECT -216.725 1.065 -216.435 2.230 ;
        RECT -216.195 1.945 -216.025 2.230 ;
        RECT -207.215 2.400 -207.045 2.470 ;
        RECT -206.275 2.400 -206.105 2.470 ;
        RECT -207.215 2.230 -206.105 2.400 ;
        RECT -207.215 1.945 -207.045 2.230 ;
        RECT -216.195 1.615 -215.265 1.945 ;
        RECT -207.975 1.615 -207.045 1.945 ;
        RECT -216.195 1.090 -216.025 1.615 ;
        RECT -207.215 1.090 -207.045 1.615 ;
        RECT -206.805 1.065 -206.515 2.230 ;
        RECT -206.275 1.945 -206.105 2.230 ;
        RECT -197.295 2.400 -197.125 2.470 ;
        RECT -196.355 2.400 -196.185 2.470 ;
        RECT -197.295 2.230 -196.185 2.400 ;
        RECT -197.295 1.945 -197.125 2.230 ;
        RECT -206.275 1.615 -205.345 1.945 ;
        RECT -198.055 1.615 -197.125 1.945 ;
        RECT -206.275 1.090 -206.105 1.615 ;
        RECT -197.295 1.090 -197.125 1.615 ;
        RECT -196.885 1.065 -196.595 2.230 ;
        RECT -196.355 1.945 -196.185 2.230 ;
        RECT -187.375 2.400 -187.205 2.470 ;
        RECT -186.435 2.400 -186.265 2.470 ;
        RECT -187.375 2.230 -186.265 2.400 ;
        RECT -187.375 1.945 -187.205 2.230 ;
        RECT -196.355 1.615 -195.425 1.945 ;
        RECT -188.135 1.615 -187.205 1.945 ;
        RECT -196.355 1.090 -196.185 1.615 ;
        RECT -187.375 1.090 -187.205 1.615 ;
        RECT -186.965 1.065 -186.675 2.230 ;
        RECT -186.435 1.945 -186.265 2.230 ;
        RECT -177.455 2.400 -177.285 2.470 ;
        RECT -176.515 2.400 -176.345 2.470 ;
        RECT -177.455 2.230 -176.345 2.400 ;
        RECT -177.455 1.945 -177.285 2.230 ;
        RECT -186.435 1.615 -185.505 1.945 ;
        RECT -178.215 1.615 -177.285 1.945 ;
        RECT -186.435 1.090 -186.265 1.615 ;
        RECT -177.455 1.090 -177.285 1.615 ;
        RECT -177.045 1.065 -176.755 2.230 ;
        RECT -176.515 1.945 -176.345 2.230 ;
        RECT -167.535 2.400 -167.365 2.470 ;
        RECT -166.595 2.400 -166.425 2.470 ;
        RECT -167.535 2.230 -166.425 2.400 ;
        RECT -167.535 1.945 -167.365 2.230 ;
        RECT -176.515 1.615 -175.585 1.945 ;
        RECT -168.295 1.615 -167.365 1.945 ;
        RECT -176.515 1.090 -176.345 1.615 ;
        RECT -167.535 1.090 -167.365 1.615 ;
        RECT -167.125 1.065 -166.835 2.230 ;
        RECT -166.595 1.945 -166.425 2.230 ;
        RECT -157.615 2.400 -157.445 2.470 ;
        RECT -156.675 2.400 -156.505 2.470 ;
        RECT -157.615 2.230 -156.505 2.400 ;
        RECT -157.615 1.945 -157.445 2.230 ;
        RECT -166.595 1.615 -165.665 1.945 ;
        RECT -158.375 1.615 -157.445 1.945 ;
        RECT -166.595 1.090 -166.425 1.615 ;
        RECT -157.615 1.090 -157.445 1.615 ;
        RECT -157.205 1.065 -156.915 2.230 ;
        RECT -156.675 1.945 -156.505 2.230 ;
        RECT -147.695 2.400 -147.525 2.470 ;
        RECT -146.755 2.400 -146.585 2.470 ;
        RECT -147.695 2.230 -146.585 2.400 ;
        RECT -147.695 1.945 -147.525 2.230 ;
        RECT -156.675 1.615 -155.745 1.945 ;
        RECT -148.455 1.615 -147.525 1.945 ;
        RECT -156.675 1.090 -156.505 1.615 ;
        RECT -147.695 1.090 -147.525 1.615 ;
        RECT -147.285 1.065 -146.995 2.230 ;
        RECT -146.755 1.945 -146.585 2.230 ;
        RECT -137.775 2.400 -137.605 2.470 ;
        RECT -136.835 2.400 -136.665 2.470 ;
        RECT -137.775 2.230 -136.665 2.400 ;
        RECT -137.775 1.945 -137.605 2.230 ;
        RECT -146.755 1.615 -145.825 1.945 ;
        RECT -138.535 1.615 -137.605 1.945 ;
        RECT -146.755 1.090 -146.585 1.615 ;
        RECT -137.775 1.090 -137.605 1.615 ;
        RECT -137.365 1.065 -137.075 2.230 ;
        RECT -136.835 1.945 -136.665 2.230 ;
        RECT -127.855 2.400 -127.685 2.470 ;
        RECT -126.915 2.400 -126.745 2.470 ;
        RECT -127.855 2.230 -126.745 2.400 ;
        RECT -127.855 1.945 -127.685 2.230 ;
        RECT -136.835 1.615 -135.905 1.945 ;
        RECT -128.615 1.615 -127.685 1.945 ;
        RECT -136.835 1.090 -136.665 1.615 ;
        RECT -127.855 1.090 -127.685 1.615 ;
        RECT -127.445 1.065 -127.155 2.230 ;
        RECT -126.915 1.945 -126.745 2.230 ;
        RECT -117.935 2.400 -117.765 2.470 ;
        RECT -116.995 2.400 -116.825 2.470 ;
        RECT -117.935 2.230 -116.825 2.400 ;
        RECT -117.935 1.945 -117.765 2.230 ;
        RECT -126.915 1.615 -125.985 1.945 ;
        RECT -118.695 1.615 -117.765 1.945 ;
        RECT -126.915 1.090 -126.745 1.615 ;
        RECT -117.935 1.090 -117.765 1.615 ;
        RECT -117.525 1.065 -117.235 2.230 ;
        RECT -116.995 1.945 -116.825 2.230 ;
        RECT -108.015 2.400 -107.845 2.470 ;
        RECT -107.075 2.400 -106.905 2.470 ;
        RECT -108.015 2.230 -106.905 2.400 ;
        RECT -108.015 1.945 -107.845 2.230 ;
        RECT -116.995 1.615 -116.065 1.945 ;
        RECT -108.775 1.615 -107.845 1.945 ;
        RECT -116.995 1.090 -116.825 1.615 ;
        RECT -108.015 1.090 -107.845 1.615 ;
        RECT -107.605 1.065 -107.315 2.230 ;
        RECT -107.075 1.945 -106.905 2.230 ;
        RECT -98.095 2.400 -97.925 2.470 ;
        RECT -97.155 2.400 -96.985 2.470 ;
        RECT -98.095 2.230 -96.985 2.400 ;
        RECT -98.095 1.945 -97.925 2.230 ;
        RECT -107.075 1.615 -106.145 1.945 ;
        RECT -98.855 1.615 -97.925 1.945 ;
        RECT -107.075 1.090 -106.905 1.615 ;
        RECT -98.095 1.090 -97.925 1.615 ;
        RECT -97.685 1.065 -97.395 2.230 ;
        RECT -97.155 1.945 -96.985 2.230 ;
        RECT -88.175 2.400 -88.005 2.470 ;
        RECT -87.235 2.400 -87.065 2.470 ;
        RECT -88.175 2.230 -87.065 2.400 ;
        RECT -88.175 1.945 -88.005 2.230 ;
        RECT -97.155 1.615 -96.225 1.945 ;
        RECT -88.935 1.615 -88.005 1.945 ;
        RECT -97.155 1.090 -96.985 1.615 ;
        RECT -88.175 1.090 -88.005 1.615 ;
        RECT -87.765 1.065 -87.475 2.230 ;
        RECT -87.235 1.945 -87.065 2.230 ;
        RECT -78.255 2.400 -78.085 2.470 ;
        RECT -77.315 2.400 -77.145 2.470 ;
        RECT -78.255 2.230 -77.145 2.400 ;
        RECT -78.255 1.945 -78.085 2.230 ;
        RECT -87.235 1.615 -86.305 1.945 ;
        RECT -79.015 1.615 -78.085 1.945 ;
        RECT -87.235 1.090 -87.065 1.615 ;
        RECT -78.255 1.090 -78.085 1.615 ;
        RECT -77.845 1.065 -77.555 2.230 ;
        RECT -77.315 1.945 -77.145 2.230 ;
        RECT -68.335 2.400 -68.165 2.470 ;
        RECT -67.395 2.400 -67.225 2.470 ;
        RECT -68.335 2.230 -67.225 2.400 ;
        RECT -68.335 1.945 -68.165 2.230 ;
        RECT -77.315 1.615 -76.385 1.945 ;
        RECT -69.095 1.615 -68.165 1.945 ;
        RECT -77.315 1.090 -77.145 1.615 ;
        RECT -68.335 1.090 -68.165 1.615 ;
        RECT -67.925 1.065 -67.635 2.230 ;
        RECT -67.395 1.945 -67.225 2.230 ;
        RECT -58.415 2.400 -58.245 2.470 ;
        RECT -57.475 2.400 -57.305 2.470 ;
        RECT -58.415 2.230 -57.305 2.400 ;
        RECT -58.415 1.945 -58.245 2.230 ;
        RECT -67.395 1.615 -66.465 1.945 ;
        RECT -59.175 1.615 -58.245 1.945 ;
        RECT -67.395 1.090 -67.225 1.615 ;
        RECT -58.415 1.090 -58.245 1.615 ;
        RECT -58.005 1.065 -57.715 2.230 ;
        RECT -57.475 1.945 -57.305 2.230 ;
        RECT -48.495 2.400 -48.325 2.470 ;
        RECT -47.555 2.400 -47.385 2.470 ;
        RECT -48.495 2.230 -47.385 2.400 ;
        RECT -48.495 1.945 -48.325 2.230 ;
        RECT -57.475 1.615 -56.545 1.945 ;
        RECT -49.255 1.615 -48.325 1.945 ;
        RECT -57.475 1.090 -57.305 1.615 ;
        RECT -48.495 1.090 -48.325 1.615 ;
        RECT -48.085 1.065 -47.795 2.230 ;
        RECT -47.555 1.945 -47.385 2.230 ;
        RECT -38.575 2.400 -38.405 2.470 ;
        RECT -37.635 2.400 -37.465 2.470 ;
        RECT -38.575 2.230 -37.465 2.400 ;
        RECT -38.575 1.945 -38.405 2.230 ;
        RECT -47.555 1.615 -46.625 1.945 ;
        RECT -39.335 1.615 -38.405 1.945 ;
        RECT -47.555 1.090 -47.385 1.615 ;
        RECT -38.575 1.090 -38.405 1.615 ;
        RECT -38.165 1.065 -37.875 2.230 ;
        RECT -37.635 1.945 -37.465 2.230 ;
        RECT -28.655 2.400 -28.485 2.470 ;
        RECT -27.715 2.400 -27.545 2.470 ;
        RECT -28.655 2.230 -27.545 2.400 ;
        RECT -28.655 1.945 -28.485 2.230 ;
        RECT -37.635 1.615 -36.705 1.945 ;
        RECT -29.415 1.615 -28.485 1.945 ;
        RECT -37.635 1.090 -37.465 1.615 ;
        RECT -28.655 1.090 -28.485 1.615 ;
        RECT -28.245 1.065 -27.955 2.230 ;
        RECT -27.715 1.945 -27.545 2.230 ;
        RECT -18.735 2.400 -18.565 2.470 ;
        RECT -17.795 2.400 -17.625 2.470 ;
        RECT -18.735 2.230 -17.625 2.400 ;
        RECT -18.735 1.945 -18.565 2.230 ;
        RECT -27.715 1.615 -26.785 1.945 ;
        RECT -19.495 1.615 -18.565 1.945 ;
        RECT -27.715 1.090 -27.545 1.615 ;
        RECT -18.735 1.090 -18.565 1.615 ;
        RECT -18.325 1.065 -18.035 2.230 ;
        RECT -17.795 1.945 -17.625 2.230 ;
        RECT -8.815 2.400 -8.645 2.470 ;
        RECT -7.875 2.400 -7.705 2.470 ;
        RECT -8.815 2.230 -7.705 2.400 ;
        RECT -8.815 1.945 -8.645 2.230 ;
        RECT -17.795 1.615 -16.865 1.945 ;
        RECT -9.575 1.615 -8.645 1.945 ;
        RECT -17.795 1.090 -17.625 1.615 ;
        RECT -8.815 1.090 -8.645 1.615 ;
        RECT -8.405 1.065 -8.115 2.230 ;
        RECT -7.875 1.945 -7.705 2.230 ;
        RECT 1.105 2.400 1.275 2.470 ;
        RECT 2.045 2.400 2.215 2.470 ;
        RECT 1.105 2.230 2.215 2.400 ;
        RECT 1.105 1.945 1.275 2.230 ;
        RECT -7.875 1.615 -6.945 1.945 ;
        RECT 0.345 1.615 1.275 1.945 ;
        RECT -7.875 1.090 -7.705 1.615 ;
        RECT 1.105 1.090 1.275 1.615 ;
        RECT 1.515 1.065 1.805 2.230 ;
        RECT 2.045 1.945 2.215 2.230 ;
        RECT 11.025 2.400 11.195 2.470 ;
        RECT 11.965 2.400 12.135 2.470 ;
        RECT 11.025 2.230 12.135 2.400 ;
        RECT 11.025 1.945 11.195 2.230 ;
        RECT 2.045 1.615 2.975 1.945 ;
        RECT 10.265 1.615 11.195 1.945 ;
        RECT 2.045 1.090 2.215 1.615 ;
        RECT 11.025 1.090 11.195 1.615 ;
        RECT 11.435 1.065 11.725 2.230 ;
        RECT 11.965 1.945 12.135 2.230 ;
        RECT 20.945 2.400 21.115 2.470 ;
        RECT 21.885 2.400 22.055 2.470 ;
        RECT 20.945 2.230 22.055 2.400 ;
        RECT 20.945 1.945 21.115 2.230 ;
        RECT 11.965 1.615 12.895 1.945 ;
        RECT 20.185 1.615 21.115 1.945 ;
        RECT 11.965 1.090 12.135 1.615 ;
        RECT 20.945 1.090 21.115 1.615 ;
        RECT 21.355 1.065 21.645 2.230 ;
        RECT 21.885 1.945 22.055 2.230 ;
        RECT 21.885 1.615 22.815 1.945 ;
        RECT 21.885 1.090 22.055 1.615 ;
        RECT -279.855 -86.070 -279.685 -85.920 ;
        RECT -278.915 -86.070 -278.745 -85.920 ;
        RECT -279.855 -86.240 -278.745 -86.070 ;
        RECT -279.855 -86.445 -279.685 -86.240 ;
        RECT -280.615 -86.775 -279.685 -86.445 ;
        RECT -279.855 -87.300 -279.685 -86.775 ;
        RECT -279.445 -87.405 -279.155 -86.240 ;
        RECT -278.915 -86.445 -278.745 -86.240 ;
        RECT -269.935 -86.070 -269.765 -85.920 ;
        RECT -268.995 -86.070 -268.825 -85.920 ;
        RECT -269.935 -86.240 -268.825 -86.070 ;
        RECT -269.935 -86.445 -269.765 -86.240 ;
        RECT -278.915 -86.775 -277.985 -86.445 ;
        RECT -270.695 -86.775 -269.765 -86.445 ;
        RECT -278.915 -87.300 -278.745 -86.775 ;
        RECT -269.935 -87.300 -269.765 -86.775 ;
        RECT -269.525 -87.405 -269.235 -86.240 ;
        RECT -268.995 -86.445 -268.825 -86.240 ;
        RECT -260.015 -86.070 -259.845 -85.920 ;
        RECT -259.075 -86.070 -258.905 -85.920 ;
        RECT -260.015 -86.240 -258.905 -86.070 ;
        RECT -260.015 -86.445 -259.845 -86.240 ;
        RECT -268.995 -86.775 -268.065 -86.445 ;
        RECT -260.775 -86.775 -259.845 -86.445 ;
        RECT -268.995 -87.300 -268.825 -86.775 ;
        RECT -260.015 -87.300 -259.845 -86.775 ;
        RECT -259.605 -87.405 -259.315 -86.240 ;
        RECT -259.075 -86.445 -258.905 -86.240 ;
        RECT -250.095 -86.070 -249.925 -85.920 ;
        RECT -249.155 -86.070 -248.985 -85.920 ;
        RECT -250.095 -86.240 -248.985 -86.070 ;
        RECT -250.095 -86.445 -249.925 -86.240 ;
        RECT -259.075 -86.775 -258.145 -86.445 ;
        RECT -250.855 -86.775 -249.925 -86.445 ;
        RECT -259.075 -87.300 -258.905 -86.775 ;
        RECT -250.095 -87.300 -249.925 -86.775 ;
        RECT -249.685 -87.405 -249.395 -86.240 ;
        RECT -249.155 -86.445 -248.985 -86.240 ;
        RECT -240.175 -86.070 -240.005 -85.920 ;
        RECT -239.235 -86.070 -239.065 -85.920 ;
        RECT -240.175 -86.240 -239.065 -86.070 ;
        RECT -240.175 -86.445 -240.005 -86.240 ;
        RECT -249.155 -86.775 -248.225 -86.445 ;
        RECT -240.935 -86.775 -240.005 -86.445 ;
        RECT -249.155 -87.300 -248.985 -86.775 ;
        RECT -240.175 -87.300 -240.005 -86.775 ;
        RECT -239.765 -87.405 -239.475 -86.240 ;
        RECT -239.235 -86.445 -239.065 -86.240 ;
        RECT -230.255 -86.070 -230.085 -85.920 ;
        RECT -229.315 -86.070 -229.145 -85.920 ;
        RECT -230.255 -86.240 -229.145 -86.070 ;
        RECT -230.255 -86.445 -230.085 -86.240 ;
        RECT -239.235 -86.775 -238.305 -86.445 ;
        RECT -231.015 -86.775 -230.085 -86.445 ;
        RECT -239.235 -87.300 -239.065 -86.775 ;
        RECT -230.255 -87.300 -230.085 -86.775 ;
        RECT -229.845 -87.405 -229.555 -86.240 ;
        RECT -229.315 -86.445 -229.145 -86.240 ;
        RECT -220.335 -86.070 -220.165 -85.920 ;
        RECT -219.395 -86.070 -219.225 -85.920 ;
        RECT -220.335 -86.240 -219.225 -86.070 ;
        RECT -220.335 -86.445 -220.165 -86.240 ;
        RECT -229.315 -86.775 -228.385 -86.445 ;
        RECT -221.095 -86.775 -220.165 -86.445 ;
        RECT -229.315 -87.300 -229.145 -86.775 ;
        RECT -220.335 -87.300 -220.165 -86.775 ;
        RECT -219.925 -87.405 -219.635 -86.240 ;
        RECT -219.395 -86.445 -219.225 -86.240 ;
        RECT -210.415 -86.070 -210.245 -85.920 ;
        RECT -209.475 -86.070 -209.305 -85.920 ;
        RECT -210.415 -86.240 -209.305 -86.070 ;
        RECT -210.415 -86.445 -210.245 -86.240 ;
        RECT -219.395 -86.775 -218.465 -86.445 ;
        RECT -211.175 -86.775 -210.245 -86.445 ;
        RECT -219.395 -87.300 -219.225 -86.775 ;
        RECT -210.415 -87.300 -210.245 -86.775 ;
        RECT -210.005 -87.405 -209.715 -86.240 ;
        RECT -209.475 -86.445 -209.305 -86.240 ;
        RECT -200.495 -86.070 -200.325 -85.920 ;
        RECT -199.555 -86.070 -199.385 -85.920 ;
        RECT -200.495 -86.240 -199.385 -86.070 ;
        RECT -200.495 -86.445 -200.325 -86.240 ;
        RECT -209.475 -86.775 -208.545 -86.445 ;
        RECT -201.255 -86.775 -200.325 -86.445 ;
        RECT -209.475 -87.300 -209.305 -86.775 ;
        RECT -200.495 -87.300 -200.325 -86.775 ;
        RECT -200.085 -87.405 -199.795 -86.240 ;
        RECT -199.555 -86.445 -199.385 -86.240 ;
        RECT -190.575 -86.070 -190.405 -85.920 ;
        RECT -189.635 -86.070 -189.465 -85.920 ;
        RECT -190.575 -86.240 -189.465 -86.070 ;
        RECT -190.575 -86.445 -190.405 -86.240 ;
        RECT -199.555 -86.775 -198.625 -86.445 ;
        RECT -191.335 -86.775 -190.405 -86.445 ;
        RECT -199.555 -87.300 -199.385 -86.775 ;
        RECT -190.575 -87.300 -190.405 -86.775 ;
        RECT -190.165 -87.405 -189.875 -86.240 ;
        RECT -189.635 -86.445 -189.465 -86.240 ;
        RECT -180.655 -86.070 -180.485 -85.920 ;
        RECT -179.715 -86.070 -179.545 -85.920 ;
        RECT -180.655 -86.240 -179.545 -86.070 ;
        RECT -180.655 -86.445 -180.485 -86.240 ;
        RECT -189.635 -86.775 -188.705 -86.445 ;
        RECT -181.415 -86.775 -180.485 -86.445 ;
        RECT -189.635 -87.300 -189.465 -86.775 ;
        RECT -180.655 -87.300 -180.485 -86.775 ;
        RECT -180.245 -87.405 -179.955 -86.240 ;
        RECT -179.715 -86.445 -179.545 -86.240 ;
        RECT -170.735 -86.070 -170.565 -85.920 ;
        RECT -169.795 -86.070 -169.625 -85.920 ;
        RECT -170.735 -86.240 -169.625 -86.070 ;
        RECT -170.735 -86.445 -170.565 -86.240 ;
        RECT -179.715 -86.775 -178.785 -86.445 ;
        RECT -171.495 -86.775 -170.565 -86.445 ;
        RECT -179.715 -87.300 -179.545 -86.775 ;
        RECT -170.735 -87.300 -170.565 -86.775 ;
        RECT -170.325 -87.405 -170.035 -86.240 ;
        RECT -169.795 -86.445 -169.625 -86.240 ;
        RECT -160.815 -86.070 -160.645 -85.920 ;
        RECT -159.875 -86.070 -159.705 -85.920 ;
        RECT -160.815 -86.240 -159.705 -86.070 ;
        RECT -160.815 -86.445 -160.645 -86.240 ;
        RECT -169.795 -86.775 -168.865 -86.445 ;
        RECT -161.575 -86.775 -160.645 -86.445 ;
        RECT -169.795 -87.300 -169.625 -86.775 ;
        RECT -160.815 -87.300 -160.645 -86.775 ;
        RECT -160.405 -87.405 -160.115 -86.240 ;
        RECT -159.875 -86.445 -159.705 -86.240 ;
        RECT -150.895 -86.070 -150.725 -85.920 ;
        RECT -149.955 -86.070 -149.785 -85.920 ;
        RECT -150.895 -86.240 -149.785 -86.070 ;
        RECT -150.895 -86.445 -150.725 -86.240 ;
        RECT -159.875 -86.775 -158.945 -86.445 ;
        RECT -151.655 -86.775 -150.725 -86.445 ;
        RECT -159.875 -87.300 -159.705 -86.775 ;
        RECT -150.895 -87.300 -150.725 -86.775 ;
        RECT -150.485 -87.405 -150.195 -86.240 ;
        RECT -149.955 -86.445 -149.785 -86.240 ;
        RECT -140.975 -86.070 -140.805 -85.920 ;
        RECT -140.035 -86.070 -139.865 -85.920 ;
        RECT -140.975 -86.240 -139.865 -86.070 ;
        RECT -140.975 -86.445 -140.805 -86.240 ;
        RECT -149.955 -86.775 -149.025 -86.445 ;
        RECT -141.735 -86.775 -140.805 -86.445 ;
        RECT -149.955 -87.300 -149.785 -86.775 ;
        RECT -140.975 -87.300 -140.805 -86.775 ;
        RECT -140.565 -87.405 -140.275 -86.240 ;
        RECT -140.035 -86.445 -139.865 -86.240 ;
        RECT -131.055 -86.070 -130.885 -85.920 ;
        RECT -130.115 -86.070 -129.945 -85.920 ;
        RECT -131.055 -86.240 -129.945 -86.070 ;
        RECT -131.055 -86.445 -130.885 -86.240 ;
        RECT -140.035 -86.775 -139.105 -86.445 ;
        RECT -131.815 -86.775 -130.885 -86.445 ;
        RECT -140.035 -87.300 -139.865 -86.775 ;
        RECT -131.055 -87.300 -130.885 -86.775 ;
        RECT -130.645 -87.405 -130.355 -86.240 ;
        RECT -130.115 -86.445 -129.945 -86.240 ;
        RECT -121.135 -86.070 -120.965 -85.920 ;
        RECT -120.195 -86.070 -120.025 -85.920 ;
        RECT -121.135 -86.240 -120.025 -86.070 ;
        RECT -121.135 -86.445 -120.965 -86.240 ;
        RECT -130.115 -86.775 -129.185 -86.445 ;
        RECT -121.895 -86.775 -120.965 -86.445 ;
        RECT -130.115 -87.300 -129.945 -86.775 ;
        RECT -121.135 -87.300 -120.965 -86.775 ;
        RECT -120.725 -87.405 -120.435 -86.240 ;
        RECT -120.195 -86.445 -120.025 -86.240 ;
        RECT -111.215 -86.070 -111.045 -85.920 ;
        RECT -110.275 -86.070 -110.105 -85.920 ;
        RECT -111.215 -86.240 -110.105 -86.070 ;
        RECT -111.215 -86.445 -111.045 -86.240 ;
        RECT -120.195 -86.775 -119.265 -86.445 ;
        RECT -111.975 -86.775 -111.045 -86.445 ;
        RECT -120.195 -87.300 -120.025 -86.775 ;
        RECT -111.215 -87.300 -111.045 -86.775 ;
        RECT -110.805 -87.405 -110.515 -86.240 ;
        RECT -110.275 -86.445 -110.105 -86.240 ;
        RECT -101.295 -86.070 -101.125 -85.920 ;
        RECT -100.355 -86.070 -100.185 -85.920 ;
        RECT -101.295 -86.240 -100.185 -86.070 ;
        RECT -101.295 -86.445 -101.125 -86.240 ;
        RECT -110.275 -86.775 -109.345 -86.445 ;
        RECT -102.055 -86.775 -101.125 -86.445 ;
        RECT -110.275 -87.300 -110.105 -86.775 ;
        RECT -101.295 -87.300 -101.125 -86.775 ;
        RECT -100.885 -87.405 -100.595 -86.240 ;
        RECT -100.355 -86.445 -100.185 -86.240 ;
        RECT -91.375 -86.070 -91.205 -85.920 ;
        RECT -90.435 -86.070 -90.265 -85.920 ;
        RECT -91.375 -86.240 -90.265 -86.070 ;
        RECT -91.375 -86.445 -91.205 -86.240 ;
        RECT -100.355 -86.775 -99.425 -86.445 ;
        RECT -92.135 -86.775 -91.205 -86.445 ;
        RECT -100.355 -87.300 -100.185 -86.775 ;
        RECT -91.375 -87.300 -91.205 -86.775 ;
        RECT -90.965 -87.405 -90.675 -86.240 ;
        RECT -90.435 -86.445 -90.265 -86.240 ;
        RECT -81.455 -86.070 -81.285 -85.920 ;
        RECT -80.515 -86.070 -80.345 -85.920 ;
        RECT -81.455 -86.240 -80.345 -86.070 ;
        RECT -81.455 -86.445 -81.285 -86.240 ;
        RECT -90.435 -86.775 -89.505 -86.445 ;
        RECT -82.215 -86.775 -81.285 -86.445 ;
        RECT -90.435 -87.300 -90.265 -86.775 ;
        RECT -81.455 -87.300 -81.285 -86.775 ;
        RECT -81.045 -87.405 -80.755 -86.240 ;
        RECT -80.515 -86.445 -80.345 -86.240 ;
        RECT -71.535 -86.070 -71.365 -85.920 ;
        RECT -70.595 -86.070 -70.425 -85.920 ;
        RECT -71.535 -86.240 -70.425 -86.070 ;
        RECT -71.535 -86.445 -71.365 -86.240 ;
        RECT -80.515 -86.775 -79.585 -86.445 ;
        RECT -72.295 -86.775 -71.365 -86.445 ;
        RECT -80.515 -87.300 -80.345 -86.775 ;
        RECT -71.535 -87.300 -71.365 -86.775 ;
        RECT -71.125 -87.405 -70.835 -86.240 ;
        RECT -70.595 -86.445 -70.425 -86.240 ;
        RECT -61.615 -86.070 -61.445 -85.920 ;
        RECT -60.675 -86.070 -60.505 -85.920 ;
        RECT -61.615 -86.240 -60.505 -86.070 ;
        RECT -61.615 -86.445 -61.445 -86.240 ;
        RECT -70.595 -86.775 -69.665 -86.445 ;
        RECT -62.375 -86.775 -61.445 -86.445 ;
        RECT -70.595 -87.300 -70.425 -86.775 ;
        RECT -61.615 -87.300 -61.445 -86.775 ;
        RECT -61.205 -87.405 -60.915 -86.240 ;
        RECT -60.675 -86.445 -60.505 -86.240 ;
        RECT -51.695 -86.070 -51.525 -85.920 ;
        RECT -50.755 -86.070 -50.585 -85.920 ;
        RECT -51.695 -86.240 -50.585 -86.070 ;
        RECT -51.695 -86.445 -51.525 -86.240 ;
        RECT -60.675 -86.775 -59.745 -86.445 ;
        RECT -52.455 -86.775 -51.525 -86.445 ;
        RECT -60.675 -87.300 -60.505 -86.775 ;
        RECT -51.695 -87.300 -51.525 -86.775 ;
        RECT -51.285 -87.405 -50.995 -86.240 ;
        RECT -50.755 -86.445 -50.585 -86.240 ;
        RECT -41.775 -86.070 -41.605 -85.920 ;
        RECT -40.835 -86.070 -40.665 -85.920 ;
        RECT -41.775 -86.240 -40.665 -86.070 ;
        RECT -41.775 -86.445 -41.605 -86.240 ;
        RECT -50.755 -86.775 -49.825 -86.445 ;
        RECT -42.535 -86.775 -41.605 -86.445 ;
        RECT -50.755 -87.300 -50.585 -86.775 ;
        RECT -41.775 -87.300 -41.605 -86.775 ;
        RECT -41.365 -87.405 -41.075 -86.240 ;
        RECT -40.835 -86.445 -40.665 -86.240 ;
        RECT -31.855 -86.070 -31.685 -85.920 ;
        RECT -30.915 -86.070 -30.745 -85.920 ;
        RECT -31.855 -86.240 -30.745 -86.070 ;
        RECT -31.855 -86.445 -31.685 -86.240 ;
        RECT -40.835 -86.775 -39.905 -86.445 ;
        RECT -32.615 -86.775 -31.685 -86.445 ;
        RECT -40.835 -87.300 -40.665 -86.775 ;
        RECT -31.855 -87.300 -31.685 -86.775 ;
        RECT -31.445 -87.405 -31.155 -86.240 ;
        RECT -30.915 -86.445 -30.745 -86.240 ;
        RECT -21.935 -86.070 -21.765 -85.920 ;
        RECT -20.995 -86.070 -20.825 -85.920 ;
        RECT -21.935 -86.240 -20.825 -86.070 ;
        RECT -21.935 -86.445 -21.765 -86.240 ;
        RECT -30.915 -86.775 -29.985 -86.445 ;
        RECT -22.695 -86.775 -21.765 -86.445 ;
        RECT -30.915 -87.300 -30.745 -86.775 ;
        RECT -21.935 -87.300 -21.765 -86.775 ;
        RECT -21.525 -87.405 -21.235 -86.240 ;
        RECT -20.995 -86.445 -20.825 -86.240 ;
        RECT -12.015 -86.070 -11.845 -85.920 ;
        RECT -11.075 -86.070 -10.905 -85.920 ;
        RECT -12.015 -86.240 -10.905 -86.070 ;
        RECT -12.015 -86.445 -11.845 -86.240 ;
        RECT -20.995 -86.775 -20.065 -86.445 ;
        RECT -12.775 -86.775 -11.845 -86.445 ;
        RECT -20.995 -87.300 -20.825 -86.775 ;
        RECT -12.015 -87.300 -11.845 -86.775 ;
        RECT -11.605 -87.405 -11.315 -86.240 ;
        RECT -11.075 -86.445 -10.905 -86.240 ;
        RECT -2.095 -86.070 -1.925 -85.920 ;
        RECT -1.155 -86.070 -0.985 -85.920 ;
        RECT -2.095 -86.240 -0.985 -86.070 ;
        RECT -2.095 -86.445 -1.925 -86.240 ;
        RECT -11.075 -86.775 -10.145 -86.445 ;
        RECT -2.855 -86.775 -1.925 -86.445 ;
        RECT -11.075 -87.300 -10.905 -86.775 ;
        RECT -2.095 -87.300 -1.925 -86.775 ;
        RECT -1.685 -87.405 -1.395 -86.240 ;
        RECT -1.155 -86.445 -0.985 -86.240 ;
        RECT 7.825 -86.070 7.995 -85.920 ;
        RECT 8.765 -86.070 8.935 -85.920 ;
        RECT 7.825 -86.240 8.935 -86.070 ;
        RECT 7.825 -86.445 7.995 -86.240 ;
        RECT -1.155 -86.775 -0.225 -86.445 ;
        RECT 7.065 -86.775 7.995 -86.445 ;
        RECT -1.155 -87.300 -0.985 -86.775 ;
        RECT 7.825 -87.300 7.995 -86.775 ;
        RECT 8.235 -87.405 8.525 -86.240 ;
        RECT 8.765 -86.445 8.935 -86.240 ;
        RECT 17.745 -86.070 17.915 -85.920 ;
        RECT 18.685 -86.070 18.855 -85.920 ;
        RECT 17.745 -86.240 18.855 -86.070 ;
        RECT 17.745 -86.445 17.915 -86.240 ;
        RECT 8.765 -86.775 9.695 -86.445 ;
        RECT 16.985 -86.775 17.915 -86.445 ;
        RECT 8.765 -87.300 8.935 -86.775 ;
        RECT 17.745 -87.300 17.915 -86.775 ;
        RECT 18.155 -87.405 18.445 -86.240 ;
        RECT 18.685 -86.445 18.855 -86.240 ;
        RECT 27.665 -86.070 27.835 -85.920 ;
        RECT 27.665 -86.240 28.450 -86.070 ;
        RECT 27.665 -86.445 27.835 -86.240 ;
        RECT 18.685 -86.775 19.615 -86.445 ;
        RECT 26.905 -86.775 27.835 -86.445 ;
        RECT 18.685 -87.300 18.855 -86.775 ;
        RECT 27.665 -87.300 27.835 -86.775 ;
        RECT 28.075 -87.405 28.365 -86.240 ;
        RECT -285.870 -87.815 -282.650 -87.645 ;
        RECT -275.950 -87.815 -272.730 -87.645 ;
        RECT -266.030 -87.815 -262.810 -87.645 ;
        RECT -256.110 -87.815 -252.890 -87.645 ;
        RECT -246.190 -87.815 -242.970 -87.645 ;
        RECT -236.270 -87.815 -233.050 -87.645 ;
        RECT -226.350 -87.815 -223.130 -87.645 ;
        RECT -216.430 -87.815 -213.210 -87.645 ;
        RECT -206.510 -87.815 -203.290 -87.645 ;
        RECT -196.590 -87.815 -193.370 -87.645 ;
        RECT -186.670 -87.815 -183.450 -87.645 ;
        RECT -176.750 -87.815 -173.530 -87.645 ;
        RECT -166.830 -87.815 -163.610 -87.645 ;
        RECT -156.910 -87.815 -153.690 -87.645 ;
        RECT -146.990 -87.815 -143.770 -87.645 ;
        RECT -137.070 -87.815 -133.850 -87.645 ;
        RECT -127.150 -87.815 -123.930 -87.645 ;
        RECT -117.230 -87.815 -114.010 -87.645 ;
        RECT -107.310 -87.815 -104.090 -87.645 ;
        RECT -97.390 -87.815 -94.170 -87.645 ;
        RECT -87.470 -87.815 -84.250 -87.645 ;
        RECT -77.550 -87.815 -74.330 -87.645 ;
        RECT -67.630 -87.815 -64.410 -87.645 ;
        RECT -57.710 -87.815 -54.490 -87.645 ;
        RECT -47.790 -87.815 -44.570 -87.645 ;
        RECT -37.870 -87.815 -34.650 -87.645 ;
        RECT -27.950 -87.815 -24.730 -87.645 ;
        RECT -18.030 -87.815 -14.810 -87.645 ;
        RECT -8.110 -87.815 -4.890 -87.645 ;
        RECT 1.810 -87.815 5.030 -87.645 ;
        RECT 11.730 -87.815 14.950 -87.645 ;
        RECT 21.650 -87.815 24.870 -87.645 ;
        RECT -285.785 -88.955 -285.525 -87.815 ;
        RECT -284.855 -88.955 -284.575 -87.815 ;
        RECT -284.405 -88.980 -284.115 -87.815 ;
        RECT -283.945 -88.955 -283.665 -87.815 ;
        RECT -282.995 -88.955 -282.735 -87.815 ;
        RECT -275.865 -88.955 -275.605 -87.815 ;
        RECT -274.935 -88.955 -274.655 -87.815 ;
        RECT -274.485 -88.980 -274.195 -87.815 ;
        RECT -274.025 -88.955 -273.745 -87.815 ;
        RECT -273.075 -88.955 -272.815 -87.815 ;
        RECT -265.945 -88.955 -265.685 -87.815 ;
        RECT -265.015 -88.955 -264.735 -87.815 ;
        RECT -264.565 -88.980 -264.275 -87.815 ;
        RECT -264.105 -88.955 -263.825 -87.815 ;
        RECT -263.155 -88.955 -262.895 -87.815 ;
        RECT -256.025 -88.955 -255.765 -87.815 ;
        RECT -255.095 -88.955 -254.815 -87.815 ;
        RECT -254.645 -88.980 -254.355 -87.815 ;
        RECT -254.185 -88.955 -253.905 -87.815 ;
        RECT -253.235 -88.955 -252.975 -87.815 ;
        RECT -246.105 -88.955 -245.845 -87.815 ;
        RECT -245.175 -88.955 -244.895 -87.815 ;
        RECT -244.725 -88.980 -244.435 -87.815 ;
        RECT -244.265 -88.955 -243.985 -87.815 ;
        RECT -243.315 -88.955 -243.055 -87.815 ;
        RECT -236.185 -88.955 -235.925 -87.815 ;
        RECT -235.255 -88.955 -234.975 -87.815 ;
        RECT -234.805 -88.980 -234.515 -87.815 ;
        RECT -234.345 -88.955 -234.065 -87.815 ;
        RECT -233.395 -88.955 -233.135 -87.815 ;
        RECT -226.265 -88.955 -226.005 -87.815 ;
        RECT -225.335 -88.955 -225.055 -87.815 ;
        RECT -224.885 -88.980 -224.595 -87.815 ;
        RECT -224.425 -88.955 -224.145 -87.815 ;
        RECT -223.475 -88.955 -223.215 -87.815 ;
        RECT -216.345 -88.955 -216.085 -87.815 ;
        RECT -215.415 -88.955 -215.135 -87.815 ;
        RECT -214.965 -88.980 -214.675 -87.815 ;
        RECT -214.505 -88.955 -214.225 -87.815 ;
        RECT -213.555 -88.955 -213.295 -87.815 ;
        RECT -206.425 -88.955 -206.165 -87.815 ;
        RECT -205.495 -88.955 -205.215 -87.815 ;
        RECT -205.045 -88.980 -204.755 -87.815 ;
        RECT -204.585 -88.955 -204.305 -87.815 ;
        RECT -203.635 -88.955 -203.375 -87.815 ;
        RECT -196.505 -88.955 -196.245 -87.815 ;
        RECT -195.575 -88.955 -195.295 -87.815 ;
        RECT -195.125 -88.980 -194.835 -87.815 ;
        RECT -194.665 -88.955 -194.385 -87.815 ;
        RECT -193.715 -88.955 -193.455 -87.815 ;
        RECT -186.585 -88.955 -186.325 -87.815 ;
        RECT -185.655 -88.955 -185.375 -87.815 ;
        RECT -185.205 -88.980 -184.915 -87.815 ;
        RECT -184.745 -88.955 -184.465 -87.815 ;
        RECT -183.795 -88.955 -183.535 -87.815 ;
        RECT -176.665 -88.955 -176.405 -87.815 ;
        RECT -175.735 -88.955 -175.455 -87.815 ;
        RECT -175.285 -88.980 -174.995 -87.815 ;
        RECT -174.825 -88.955 -174.545 -87.815 ;
        RECT -173.875 -88.955 -173.615 -87.815 ;
        RECT -166.745 -88.955 -166.485 -87.815 ;
        RECT -165.815 -88.955 -165.535 -87.815 ;
        RECT -165.365 -88.980 -165.075 -87.815 ;
        RECT -164.905 -88.955 -164.625 -87.815 ;
        RECT -163.955 -88.955 -163.695 -87.815 ;
        RECT -156.825 -88.955 -156.565 -87.815 ;
        RECT -155.895 -88.955 -155.615 -87.815 ;
        RECT -155.445 -88.980 -155.155 -87.815 ;
        RECT -154.985 -88.955 -154.705 -87.815 ;
        RECT -154.035 -88.955 -153.775 -87.815 ;
        RECT -146.905 -88.955 -146.645 -87.815 ;
        RECT -145.975 -88.955 -145.695 -87.815 ;
        RECT -145.525 -88.980 -145.235 -87.815 ;
        RECT -145.065 -88.955 -144.785 -87.815 ;
        RECT -144.115 -88.955 -143.855 -87.815 ;
        RECT -136.985 -88.955 -136.725 -87.815 ;
        RECT -136.055 -88.955 -135.775 -87.815 ;
        RECT -135.605 -88.980 -135.315 -87.815 ;
        RECT -135.145 -88.955 -134.865 -87.815 ;
        RECT -134.195 -88.955 -133.935 -87.815 ;
        RECT -127.065 -88.955 -126.805 -87.815 ;
        RECT -126.135 -88.955 -125.855 -87.815 ;
        RECT -125.685 -88.980 -125.395 -87.815 ;
        RECT -125.225 -88.955 -124.945 -87.815 ;
        RECT -124.275 -88.955 -124.015 -87.815 ;
        RECT -117.145 -88.955 -116.885 -87.815 ;
        RECT -116.215 -88.955 -115.935 -87.815 ;
        RECT -115.765 -88.980 -115.475 -87.815 ;
        RECT -115.305 -88.955 -115.025 -87.815 ;
        RECT -114.355 -88.955 -114.095 -87.815 ;
        RECT -107.225 -88.955 -106.965 -87.815 ;
        RECT -106.295 -88.955 -106.015 -87.815 ;
        RECT -105.845 -88.980 -105.555 -87.815 ;
        RECT -105.385 -88.955 -105.105 -87.815 ;
        RECT -104.435 -88.955 -104.175 -87.815 ;
        RECT -97.305 -88.955 -97.045 -87.815 ;
        RECT -96.375 -88.955 -96.095 -87.815 ;
        RECT -95.925 -88.980 -95.635 -87.815 ;
        RECT -95.465 -88.955 -95.185 -87.815 ;
        RECT -94.515 -88.955 -94.255 -87.815 ;
        RECT -87.385 -88.955 -87.125 -87.815 ;
        RECT -86.455 -88.955 -86.175 -87.815 ;
        RECT -86.005 -88.980 -85.715 -87.815 ;
        RECT -85.545 -88.955 -85.265 -87.815 ;
        RECT -84.595 -88.955 -84.335 -87.815 ;
        RECT -77.465 -88.955 -77.205 -87.815 ;
        RECT -76.535 -88.955 -76.255 -87.815 ;
        RECT -76.085 -88.980 -75.795 -87.815 ;
        RECT -75.625 -88.955 -75.345 -87.815 ;
        RECT -74.675 -88.955 -74.415 -87.815 ;
        RECT -67.545 -88.955 -67.285 -87.815 ;
        RECT -66.615 -88.955 -66.335 -87.815 ;
        RECT -66.165 -88.980 -65.875 -87.815 ;
        RECT -65.705 -88.955 -65.425 -87.815 ;
        RECT -64.755 -88.955 -64.495 -87.815 ;
        RECT -57.625 -88.955 -57.365 -87.815 ;
        RECT -56.695 -88.955 -56.415 -87.815 ;
        RECT -56.245 -88.980 -55.955 -87.815 ;
        RECT -55.785 -88.955 -55.505 -87.815 ;
        RECT -54.835 -88.955 -54.575 -87.815 ;
        RECT -47.705 -88.955 -47.445 -87.815 ;
        RECT -46.775 -88.955 -46.495 -87.815 ;
        RECT -46.325 -88.980 -46.035 -87.815 ;
        RECT -45.865 -88.955 -45.585 -87.815 ;
        RECT -44.915 -88.955 -44.655 -87.815 ;
        RECT -37.785 -88.955 -37.525 -87.815 ;
        RECT -36.855 -88.955 -36.575 -87.815 ;
        RECT -36.405 -88.980 -36.115 -87.815 ;
        RECT -35.945 -88.955 -35.665 -87.815 ;
        RECT -34.995 -88.955 -34.735 -87.815 ;
        RECT -27.865 -88.955 -27.605 -87.815 ;
        RECT -26.935 -88.955 -26.655 -87.815 ;
        RECT -26.485 -88.980 -26.195 -87.815 ;
        RECT -26.025 -88.955 -25.745 -87.815 ;
        RECT -25.075 -88.955 -24.815 -87.815 ;
        RECT -17.945 -88.955 -17.685 -87.815 ;
        RECT -17.015 -88.955 -16.735 -87.815 ;
        RECT -16.565 -88.980 -16.275 -87.815 ;
        RECT -16.105 -88.955 -15.825 -87.815 ;
        RECT -15.155 -88.955 -14.895 -87.815 ;
        RECT -8.025 -88.955 -7.765 -87.815 ;
        RECT -7.095 -88.955 -6.815 -87.815 ;
        RECT -6.645 -88.980 -6.355 -87.815 ;
        RECT -6.185 -88.955 -5.905 -87.815 ;
        RECT -5.235 -88.955 -4.975 -87.815 ;
        RECT 1.895 -88.955 2.155 -87.815 ;
        RECT 2.825 -88.955 3.105 -87.815 ;
        RECT 3.275 -88.980 3.565 -87.815 ;
        RECT 3.735 -88.955 4.015 -87.815 ;
        RECT 4.685 -88.955 4.945 -87.815 ;
        RECT 11.815 -88.955 12.075 -87.815 ;
        RECT 12.745 -88.955 13.025 -87.815 ;
        RECT 13.195 -88.980 13.485 -87.815 ;
        RECT 13.655 -88.955 13.935 -87.815 ;
        RECT 14.605 -88.955 14.865 -87.815 ;
        RECT 21.735 -88.955 21.995 -87.815 ;
        RECT 22.665 -88.955 22.945 -87.815 ;
        RECT 23.115 -88.980 23.405 -87.815 ;
        RECT 23.575 -88.955 23.855 -87.815 ;
        RECT 24.525 -88.955 24.785 -87.815 ;
        RECT -280.825 -90.365 -280.565 -89.225 ;
        RECT -279.895 -90.365 -279.615 -89.225 ;
        RECT -279.445 -90.365 -279.155 -89.200 ;
        RECT -278.985 -90.365 -278.705 -89.225 ;
        RECT -278.035 -90.365 -277.775 -89.225 ;
        RECT -270.905 -90.365 -270.645 -89.225 ;
        RECT -269.975 -90.365 -269.695 -89.225 ;
        RECT -269.525 -90.365 -269.235 -89.200 ;
        RECT -269.065 -90.365 -268.785 -89.225 ;
        RECT -268.115 -90.365 -267.855 -89.225 ;
        RECT -260.985 -90.365 -260.725 -89.225 ;
        RECT -260.055 -90.365 -259.775 -89.225 ;
        RECT -259.605 -90.365 -259.315 -89.200 ;
        RECT -259.145 -90.365 -258.865 -89.225 ;
        RECT -258.195 -90.365 -257.935 -89.225 ;
        RECT -251.065 -90.365 -250.805 -89.225 ;
        RECT -250.135 -90.365 -249.855 -89.225 ;
        RECT -249.685 -90.365 -249.395 -89.200 ;
        RECT -249.225 -90.365 -248.945 -89.225 ;
        RECT -248.275 -90.365 -248.015 -89.225 ;
        RECT -241.145 -90.365 -240.885 -89.225 ;
        RECT -240.215 -90.365 -239.935 -89.225 ;
        RECT -239.765 -90.365 -239.475 -89.200 ;
        RECT -239.305 -90.365 -239.025 -89.225 ;
        RECT -238.355 -90.365 -238.095 -89.225 ;
        RECT -231.225 -90.365 -230.965 -89.225 ;
        RECT -230.295 -90.365 -230.015 -89.225 ;
        RECT -229.845 -90.365 -229.555 -89.200 ;
        RECT -229.385 -90.365 -229.105 -89.225 ;
        RECT -228.435 -90.365 -228.175 -89.225 ;
        RECT -221.305 -90.365 -221.045 -89.225 ;
        RECT -220.375 -90.365 -220.095 -89.225 ;
        RECT -219.925 -90.365 -219.635 -89.200 ;
        RECT -219.465 -90.365 -219.185 -89.225 ;
        RECT -218.515 -90.365 -218.255 -89.225 ;
        RECT -211.385 -90.365 -211.125 -89.225 ;
        RECT -210.455 -90.365 -210.175 -89.225 ;
        RECT -210.005 -90.365 -209.715 -89.200 ;
        RECT -209.545 -90.365 -209.265 -89.225 ;
        RECT -208.595 -90.365 -208.335 -89.225 ;
        RECT -201.465 -90.365 -201.205 -89.225 ;
        RECT -200.535 -90.365 -200.255 -89.225 ;
        RECT -200.085 -90.365 -199.795 -89.200 ;
        RECT -199.625 -90.365 -199.345 -89.225 ;
        RECT -198.675 -90.365 -198.415 -89.225 ;
        RECT -191.545 -90.365 -191.285 -89.225 ;
        RECT -190.615 -90.365 -190.335 -89.225 ;
        RECT -190.165 -90.365 -189.875 -89.200 ;
        RECT -189.705 -90.365 -189.425 -89.225 ;
        RECT -188.755 -90.365 -188.495 -89.225 ;
        RECT -181.625 -90.365 -181.365 -89.225 ;
        RECT -180.695 -90.365 -180.415 -89.225 ;
        RECT -180.245 -90.365 -179.955 -89.200 ;
        RECT -179.785 -90.365 -179.505 -89.225 ;
        RECT -178.835 -90.365 -178.575 -89.225 ;
        RECT -171.705 -90.365 -171.445 -89.225 ;
        RECT -170.775 -90.365 -170.495 -89.225 ;
        RECT -170.325 -90.365 -170.035 -89.200 ;
        RECT -169.865 -90.365 -169.585 -89.225 ;
        RECT -168.915 -90.365 -168.655 -89.225 ;
        RECT -161.785 -90.365 -161.525 -89.225 ;
        RECT -160.855 -90.365 -160.575 -89.225 ;
        RECT -160.405 -90.365 -160.115 -89.200 ;
        RECT -159.945 -90.365 -159.665 -89.225 ;
        RECT -158.995 -90.365 -158.735 -89.225 ;
        RECT -151.865 -90.365 -151.605 -89.225 ;
        RECT -150.935 -90.365 -150.655 -89.225 ;
        RECT -150.485 -90.365 -150.195 -89.200 ;
        RECT -150.025 -90.365 -149.745 -89.225 ;
        RECT -149.075 -90.365 -148.815 -89.225 ;
        RECT -141.945 -90.365 -141.685 -89.225 ;
        RECT -141.015 -90.365 -140.735 -89.225 ;
        RECT -140.565 -90.365 -140.275 -89.200 ;
        RECT -140.105 -90.365 -139.825 -89.225 ;
        RECT -139.155 -90.365 -138.895 -89.225 ;
        RECT -132.025 -90.365 -131.765 -89.225 ;
        RECT -131.095 -90.365 -130.815 -89.225 ;
        RECT -130.645 -90.365 -130.355 -89.200 ;
        RECT -130.185 -90.365 -129.905 -89.225 ;
        RECT -129.235 -90.365 -128.975 -89.225 ;
        RECT -122.105 -90.365 -121.845 -89.225 ;
        RECT -121.175 -90.365 -120.895 -89.225 ;
        RECT -120.725 -90.365 -120.435 -89.200 ;
        RECT -120.265 -90.365 -119.985 -89.225 ;
        RECT -119.315 -90.365 -119.055 -89.225 ;
        RECT -112.185 -90.365 -111.925 -89.225 ;
        RECT -111.255 -90.365 -110.975 -89.225 ;
        RECT -110.805 -90.365 -110.515 -89.200 ;
        RECT -110.345 -90.365 -110.065 -89.225 ;
        RECT -109.395 -90.365 -109.135 -89.225 ;
        RECT -102.265 -90.365 -102.005 -89.225 ;
        RECT -101.335 -90.365 -101.055 -89.225 ;
        RECT -100.885 -90.365 -100.595 -89.200 ;
        RECT -100.425 -90.365 -100.145 -89.225 ;
        RECT -99.475 -90.365 -99.215 -89.225 ;
        RECT -92.345 -90.365 -92.085 -89.225 ;
        RECT -91.415 -90.365 -91.135 -89.225 ;
        RECT -90.965 -90.365 -90.675 -89.200 ;
        RECT -90.505 -90.365 -90.225 -89.225 ;
        RECT -89.555 -90.365 -89.295 -89.225 ;
        RECT -82.425 -90.365 -82.165 -89.225 ;
        RECT -81.495 -90.365 -81.215 -89.225 ;
        RECT -81.045 -90.365 -80.755 -89.200 ;
        RECT -80.585 -90.365 -80.305 -89.225 ;
        RECT -79.635 -90.365 -79.375 -89.225 ;
        RECT -72.505 -90.365 -72.245 -89.225 ;
        RECT -71.575 -90.365 -71.295 -89.225 ;
        RECT -71.125 -90.365 -70.835 -89.200 ;
        RECT -70.665 -90.365 -70.385 -89.225 ;
        RECT -69.715 -90.365 -69.455 -89.225 ;
        RECT -62.585 -90.365 -62.325 -89.225 ;
        RECT -61.655 -90.365 -61.375 -89.225 ;
        RECT -61.205 -90.365 -60.915 -89.200 ;
        RECT -60.745 -90.365 -60.465 -89.225 ;
        RECT -59.795 -90.365 -59.535 -89.225 ;
        RECT -52.665 -90.365 -52.405 -89.225 ;
        RECT -51.735 -90.365 -51.455 -89.225 ;
        RECT -51.285 -90.365 -50.995 -89.200 ;
        RECT -50.825 -90.365 -50.545 -89.225 ;
        RECT -49.875 -90.365 -49.615 -89.225 ;
        RECT -42.745 -90.365 -42.485 -89.225 ;
        RECT -41.815 -90.365 -41.535 -89.225 ;
        RECT -41.365 -90.365 -41.075 -89.200 ;
        RECT -40.905 -90.365 -40.625 -89.225 ;
        RECT -39.955 -90.365 -39.695 -89.225 ;
        RECT -32.825 -90.365 -32.565 -89.225 ;
        RECT -31.895 -90.365 -31.615 -89.225 ;
        RECT -31.445 -90.365 -31.155 -89.200 ;
        RECT -30.985 -90.365 -30.705 -89.225 ;
        RECT -30.035 -90.365 -29.775 -89.225 ;
        RECT -22.905 -90.365 -22.645 -89.225 ;
        RECT -21.975 -90.365 -21.695 -89.225 ;
        RECT -21.525 -90.365 -21.235 -89.200 ;
        RECT -21.065 -90.365 -20.785 -89.225 ;
        RECT -20.115 -90.365 -19.855 -89.225 ;
        RECT -12.985 -90.365 -12.725 -89.225 ;
        RECT -12.055 -90.365 -11.775 -89.225 ;
        RECT -11.605 -90.365 -11.315 -89.200 ;
        RECT -11.145 -90.365 -10.865 -89.225 ;
        RECT -10.195 -90.365 -9.935 -89.225 ;
        RECT -3.065 -90.365 -2.805 -89.225 ;
        RECT -2.135 -90.365 -1.855 -89.225 ;
        RECT -1.685 -90.365 -1.395 -89.200 ;
        RECT -1.225 -90.365 -0.945 -89.225 ;
        RECT -0.275 -90.365 -0.015 -89.225 ;
        RECT 6.855 -90.365 7.115 -89.225 ;
        RECT 7.785 -90.365 8.065 -89.225 ;
        RECT 8.235 -90.365 8.525 -89.200 ;
        RECT 8.695 -90.365 8.975 -89.225 ;
        RECT 9.645 -90.365 9.905 -89.225 ;
        RECT 16.775 -90.365 17.035 -89.225 ;
        RECT 17.705 -90.365 17.985 -89.225 ;
        RECT 18.155 -90.365 18.445 -89.200 ;
        RECT 18.615 -90.365 18.895 -89.225 ;
        RECT 19.565 -90.365 19.825 -89.225 ;
        RECT 26.695 -90.365 26.955 -89.225 ;
        RECT 27.625 -90.365 27.905 -89.225 ;
        RECT 28.075 -90.365 28.365 -89.200 ;
        RECT -280.910 -90.535 -277.690 -90.365 ;
        RECT -270.990 -90.535 -267.770 -90.365 ;
        RECT -261.070 -90.535 -257.850 -90.365 ;
        RECT -251.150 -90.535 -247.930 -90.365 ;
        RECT -241.230 -90.535 -238.010 -90.365 ;
        RECT -231.310 -90.535 -228.090 -90.365 ;
        RECT -221.390 -90.535 -218.170 -90.365 ;
        RECT -211.470 -90.535 -208.250 -90.365 ;
        RECT -201.550 -90.535 -198.330 -90.365 ;
        RECT -191.630 -90.535 -188.410 -90.365 ;
        RECT -181.710 -90.535 -178.490 -90.365 ;
        RECT -171.790 -90.535 -168.570 -90.365 ;
        RECT -161.870 -90.535 -158.650 -90.365 ;
        RECT -151.950 -90.535 -148.730 -90.365 ;
        RECT -142.030 -90.535 -138.810 -90.365 ;
        RECT -132.110 -90.535 -128.890 -90.365 ;
        RECT -122.190 -90.535 -118.970 -90.365 ;
        RECT -112.270 -90.535 -109.050 -90.365 ;
        RECT -102.350 -90.535 -99.130 -90.365 ;
        RECT -92.430 -90.535 -89.210 -90.365 ;
        RECT -82.510 -90.535 -79.290 -90.365 ;
        RECT -72.590 -90.535 -69.370 -90.365 ;
        RECT -62.670 -90.535 -59.450 -90.365 ;
        RECT -52.750 -90.535 -49.530 -90.365 ;
        RECT -42.830 -90.535 -39.610 -90.365 ;
        RECT -32.910 -90.535 -29.690 -90.365 ;
        RECT -22.990 -90.535 -19.770 -90.365 ;
        RECT -13.070 -90.535 -9.850 -90.365 ;
        RECT -3.150 -90.535 0.070 -90.365 ;
        RECT 6.770 -90.535 9.990 -90.365 ;
        RECT 16.690 -90.535 19.910 -90.365 ;
        RECT 26.610 -90.535 28.450 -90.365 ;
        RECT -284.815 -90.950 -284.645 -90.880 ;
        RECT -283.875 -90.950 -283.705 -90.880 ;
        RECT -284.815 -91.120 -283.705 -90.950 ;
        RECT -284.815 -91.405 -284.645 -91.120 ;
        RECT -285.575 -91.735 -284.645 -91.405 ;
        RECT -284.815 -92.260 -284.645 -91.735 ;
        RECT -284.405 -92.285 -284.115 -91.120 ;
        RECT -283.875 -91.405 -283.705 -91.120 ;
        RECT -274.895 -90.950 -274.725 -90.880 ;
        RECT -273.955 -90.950 -273.785 -90.880 ;
        RECT -274.895 -91.120 -273.785 -90.950 ;
        RECT -274.895 -91.405 -274.725 -91.120 ;
        RECT -283.875 -91.735 -282.945 -91.405 ;
        RECT -275.655 -91.735 -274.725 -91.405 ;
        RECT -283.875 -92.260 -283.705 -91.735 ;
        RECT -274.895 -92.260 -274.725 -91.735 ;
        RECT -274.485 -92.285 -274.195 -91.120 ;
        RECT -273.955 -91.405 -273.785 -91.120 ;
        RECT -264.975 -90.950 -264.805 -90.880 ;
        RECT -264.035 -90.950 -263.865 -90.880 ;
        RECT -264.975 -91.120 -263.865 -90.950 ;
        RECT -264.975 -91.405 -264.805 -91.120 ;
        RECT -273.955 -91.735 -273.025 -91.405 ;
        RECT -265.735 -91.735 -264.805 -91.405 ;
        RECT -273.955 -92.260 -273.785 -91.735 ;
        RECT -264.975 -92.260 -264.805 -91.735 ;
        RECT -264.565 -92.285 -264.275 -91.120 ;
        RECT -264.035 -91.405 -263.865 -91.120 ;
        RECT -255.055 -90.950 -254.885 -90.880 ;
        RECT -254.115 -90.950 -253.945 -90.880 ;
        RECT -255.055 -91.120 -253.945 -90.950 ;
        RECT -255.055 -91.405 -254.885 -91.120 ;
        RECT -264.035 -91.735 -263.105 -91.405 ;
        RECT -255.815 -91.735 -254.885 -91.405 ;
        RECT -264.035 -92.260 -263.865 -91.735 ;
        RECT -255.055 -92.260 -254.885 -91.735 ;
        RECT -254.645 -92.285 -254.355 -91.120 ;
        RECT -254.115 -91.405 -253.945 -91.120 ;
        RECT -245.135 -90.950 -244.965 -90.880 ;
        RECT -244.195 -90.950 -244.025 -90.880 ;
        RECT -245.135 -91.120 -244.025 -90.950 ;
        RECT -245.135 -91.405 -244.965 -91.120 ;
        RECT -254.115 -91.735 -253.185 -91.405 ;
        RECT -245.895 -91.735 -244.965 -91.405 ;
        RECT -254.115 -92.260 -253.945 -91.735 ;
        RECT -245.135 -92.260 -244.965 -91.735 ;
        RECT -244.725 -92.285 -244.435 -91.120 ;
        RECT -244.195 -91.405 -244.025 -91.120 ;
        RECT -235.215 -90.950 -235.045 -90.880 ;
        RECT -234.275 -90.950 -234.105 -90.880 ;
        RECT -235.215 -91.120 -234.105 -90.950 ;
        RECT -235.215 -91.405 -235.045 -91.120 ;
        RECT -244.195 -91.735 -243.265 -91.405 ;
        RECT -235.975 -91.735 -235.045 -91.405 ;
        RECT -244.195 -92.260 -244.025 -91.735 ;
        RECT -235.215 -92.260 -235.045 -91.735 ;
        RECT -234.805 -92.285 -234.515 -91.120 ;
        RECT -234.275 -91.405 -234.105 -91.120 ;
        RECT -225.295 -90.950 -225.125 -90.880 ;
        RECT -224.355 -90.950 -224.185 -90.880 ;
        RECT -225.295 -91.120 -224.185 -90.950 ;
        RECT -225.295 -91.405 -225.125 -91.120 ;
        RECT -234.275 -91.735 -233.345 -91.405 ;
        RECT -226.055 -91.735 -225.125 -91.405 ;
        RECT -234.275 -92.260 -234.105 -91.735 ;
        RECT -225.295 -92.260 -225.125 -91.735 ;
        RECT -224.885 -92.285 -224.595 -91.120 ;
        RECT -224.355 -91.405 -224.185 -91.120 ;
        RECT -215.375 -90.950 -215.205 -90.880 ;
        RECT -214.435 -90.950 -214.265 -90.880 ;
        RECT -215.375 -91.120 -214.265 -90.950 ;
        RECT -215.375 -91.405 -215.205 -91.120 ;
        RECT -224.355 -91.735 -223.425 -91.405 ;
        RECT -216.135 -91.735 -215.205 -91.405 ;
        RECT -224.355 -92.260 -224.185 -91.735 ;
        RECT -215.375 -92.260 -215.205 -91.735 ;
        RECT -214.965 -92.285 -214.675 -91.120 ;
        RECT -214.435 -91.405 -214.265 -91.120 ;
        RECT -205.455 -90.950 -205.285 -90.880 ;
        RECT -204.515 -90.950 -204.345 -90.880 ;
        RECT -205.455 -91.120 -204.345 -90.950 ;
        RECT -205.455 -91.405 -205.285 -91.120 ;
        RECT -214.435 -91.735 -213.505 -91.405 ;
        RECT -206.215 -91.735 -205.285 -91.405 ;
        RECT -214.435 -92.260 -214.265 -91.735 ;
        RECT -205.455 -92.260 -205.285 -91.735 ;
        RECT -205.045 -92.285 -204.755 -91.120 ;
        RECT -204.515 -91.405 -204.345 -91.120 ;
        RECT -195.535 -90.950 -195.365 -90.880 ;
        RECT -194.595 -90.950 -194.425 -90.880 ;
        RECT -195.535 -91.120 -194.425 -90.950 ;
        RECT -195.535 -91.405 -195.365 -91.120 ;
        RECT -204.515 -91.735 -203.585 -91.405 ;
        RECT -196.295 -91.735 -195.365 -91.405 ;
        RECT -204.515 -92.260 -204.345 -91.735 ;
        RECT -195.535 -92.260 -195.365 -91.735 ;
        RECT -195.125 -92.285 -194.835 -91.120 ;
        RECT -194.595 -91.405 -194.425 -91.120 ;
        RECT -185.615 -90.950 -185.445 -90.880 ;
        RECT -184.675 -90.950 -184.505 -90.880 ;
        RECT -185.615 -91.120 -184.505 -90.950 ;
        RECT -185.615 -91.405 -185.445 -91.120 ;
        RECT -194.595 -91.735 -193.665 -91.405 ;
        RECT -186.375 -91.735 -185.445 -91.405 ;
        RECT -194.595 -92.260 -194.425 -91.735 ;
        RECT -185.615 -92.260 -185.445 -91.735 ;
        RECT -185.205 -92.285 -184.915 -91.120 ;
        RECT -184.675 -91.405 -184.505 -91.120 ;
        RECT -175.695 -90.950 -175.525 -90.880 ;
        RECT -174.755 -90.950 -174.585 -90.880 ;
        RECT -175.695 -91.120 -174.585 -90.950 ;
        RECT -175.695 -91.405 -175.525 -91.120 ;
        RECT -184.675 -91.735 -183.745 -91.405 ;
        RECT -176.455 -91.735 -175.525 -91.405 ;
        RECT -184.675 -92.260 -184.505 -91.735 ;
        RECT -175.695 -92.260 -175.525 -91.735 ;
        RECT -175.285 -92.285 -174.995 -91.120 ;
        RECT -174.755 -91.405 -174.585 -91.120 ;
        RECT -165.775 -90.950 -165.605 -90.880 ;
        RECT -164.835 -90.950 -164.665 -90.880 ;
        RECT -165.775 -91.120 -164.665 -90.950 ;
        RECT -165.775 -91.405 -165.605 -91.120 ;
        RECT -174.755 -91.735 -173.825 -91.405 ;
        RECT -166.535 -91.735 -165.605 -91.405 ;
        RECT -174.755 -92.260 -174.585 -91.735 ;
        RECT -165.775 -92.260 -165.605 -91.735 ;
        RECT -165.365 -92.285 -165.075 -91.120 ;
        RECT -164.835 -91.405 -164.665 -91.120 ;
        RECT -155.855 -90.950 -155.685 -90.880 ;
        RECT -154.915 -90.950 -154.745 -90.880 ;
        RECT -155.855 -91.120 -154.745 -90.950 ;
        RECT -155.855 -91.405 -155.685 -91.120 ;
        RECT -164.835 -91.735 -163.905 -91.405 ;
        RECT -156.615 -91.735 -155.685 -91.405 ;
        RECT -164.835 -92.260 -164.665 -91.735 ;
        RECT -155.855 -92.260 -155.685 -91.735 ;
        RECT -155.445 -92.285 -155.155 -91.120 ;
        RECT -154.915 -91.405 -154.745 -91.120 ;
        RECT -145.935 -90.950 -145.765 -90.880 ;
        RECT -144.995 -90.950 -144.825 -90.880 ;
        RECT -145.935 -91.120 -144.825 -90.950 ;
        RECT -145.935 -91.405 -145.765 -91.120 ;
        RECT -154.915 -91.735 -153.985 -91.405 ;
        RECT -146.695 -91.735 -145.765 -91.405 ;
        RECT -154.915 -92.260 -154.745 -91.735 ;
        RECT -145.935 -92.260 -145.765 -91.735 ;
        RECT -145.525 -92.285 -145.235 -91.120 ;
        RECT -144.995 -91.405 -144.825 -91.120 ;
        RECT -136.015 -90.950 -135.845 -90.880 ;
        RECT -135.075 -90.950 -134.905 -90.880 ;
        RECT -136.015 -91.120 -134.905 -90.950 ;
        RECT -136.015 -91.405 -135.845 -91.120 ;
        RECT -144.995 -91.735 -144.065 -91.405 ;
        RECT -136.775 -91.735 -135.845 -91.405 ;
        RECT -144.995 -92.260 -144.825 -91.735 ;
        RECT -136.015 -92.260 -135.845 -91.735 ;
        RECT -135.605 -92.285 -135.315 -91.120 ;
        RECT -135.075 -91.405 -134.905 -91.120 ;
        RECT -126.095 -90.950 -125.925 -90.880 ;
        RECT -125.155 -90.950 -124.985 -90.880 ;
        RECT -126.095 -91.120 -124.985 -90.950 ;
        RECT -126.095 -91.405 -125.925 -91.120 ;
        RECT -135.075 -91.735 -134.145 -91.405 ;
        RECT -126.855 -91.735 -125.925 -91.405 ;
        RECT -135.075 -92.260 -134.905 -91.735 ;
        RECT -126.095 -92.260 -125.925 -91.735 ;
        RECT -125.685 -92.285 -125.395 -91.120 ;
        RECT -125.155 -91.405 -124.985 -91.120 ;
        RECT -116.175 -90.950 -116.005 -90.880 ;
        RECT -115.235 -90.950 -115.065 -90.880 ;
        RECT -116.175 -91.120 -115.065 -90.950 ;
        RECT -116.175 -91.405 -116.005 -91.120 ;
        RECT -125.155 -91.735 -124.225 -91.405 ;
        RECT -116.935 -91.735 -116.005 -91.405 ;
        RECT -125.155 -92.260 -124.985 -91.735 ;
        RECT -116.175 -92.260 -116.005 -91.735 ;
        RECT -115.765 -92.285 -115.475 -91.120 ;
        RECT -115.235 -91.405 -115.065 -91.120 ;
        RECT -106.255 -90.950 -106.085 -90.880 ;
        RECT -105.315 -90.950 -105.145 -90.880 ;
        RECT -106.255 -91.120 -105.145 -90.950 ;
        RECT -106.255 -91.405 -106.085 -91.120 ;
        RECT -115.235 -91.735 -114.305 -91.405 ;
        RECT -107.015 -91.735 -106.085 -91.405 ;
        RECT -115.235 -92.260 -115.065 -91.735 ;
        RECT -106.255 -92.260 -106.085 -91.735 ;
        RECT -105.845 -92.285 -105.555 -91.120 ;
        RECT -105.315 -91.405 -105.145 -91.120 ;
        RECT -96.335 -90.950 -96.165 -90.880 ;
        RECT -95.395 -90.950 -95.225 -90.880 ;
        RECT -96.335 -91.120 -95.225 -90.950 ;
        RECT -96.335 -91.405 -96.165 -91.120 ;
        RECT -105.315 -91.735 -104.385 -91.405 ;
        RECT -97.095 -91.735 -96.165 -91.405 ;
        RECT -105.315 -92.260 -105.145 -91.735 ;
        RECT -96.335 -92.260 -96.165 -91.735 ;
        RECT -95.925 -92.285 -95.635 -91.120 ;
        RECT -95.395 -91.405 -95.225 -91.120 ;
        RECT -86.415 -90.950 -86.245 -90.880 ;
        RECT -85.475 -90.950 -85.305 -90.880 ;
        RECT -86.415 -91.120 -85.305 -90.950 ;
        RECT -86.415 -91.405 -86.245 -91.120 ;
        RECT -95.395 -91.735 -94.465 -91.405 ;
        RECT -87.175 -91.735 -86.245 -91.405 ;
        RECT -95.395 -92.260 -95.225 -91.735 ;
        RECT -86.415 -92.260 -86.245 -91.735 ;
        RECT -86.005 -92.285 -85.715 -91.120 ;
        RECT -85.475 -91.405 -85.305 -91.120 ;
        RECT -76.495 -90.950 -76.325 -90.880 ;
        RECT -75.555 -90.950 -75.385 -90.880 ;
        RECT -76.495 -91.120 -75.385 -90.950 ;
        RECT -76.495 -91.405 -76.325 -91.120 ;
        RECT -85.475 -91.735 -84.545 -91.405 ;
        RECT -77.255 -91.735 -76.325 -91.405 ;
        RECT -85.475 -92.260 -85.305 -91.735 ;
        RECT -76.495 -92.260 -76.325 -91.735 ;
        RECT -76.085 -92.285 -75.795 -91.120 ;
        RECT -75.555 -91.405 -75.385 -91.120 ;
        RECT -66.575 -90.950 -66.405 -90.880 ;
        RECT -65.635 -90.950 -65.465 -90.880 ;
        RECT -66.575 -91.120 -65.465 -90.950 ;
        RECT -66.575 -91.405 -66.405 -91.120 ;
        RECT -75.555 -91.735 -74.625 -91.405 ;
        RECT -67.335 -91.735 -66.405 -91.405 ;
        RECT -75.555 -92.260 -75.385 -91.735 ;
        RECT -66.575 -92.260 -66.405 -91.735 ;
        RECT -66.165 -92.285 -65.875 -91.120 ;
        RECT -65.635 -91.405 -65.465 -91.120 ;
        RECT -56.655 -90.950 -56.485 -90.880 ;
        RECT -55.715 -90.950 -55.545 -90.880 ;
        RECT -56.655 -91.120 -55.545 -90.950 ;
        RECT -56.655 -91.405 -56.485 -91.120 ;
        RECT -65.635 -91.735 -64.705 -91.405 ;
        RECT -57.415 -91.735 -56.485 -91.405 ;
        RECT -65.635 -92.260 -65.465 -91.735 ;
        RECT -56.655 -92.260 -56.485 -91.735 ;
        RECT -56.245 -92.285 -55.955 -91.120 ;
        RECT -55.715 -91.405 -55.545 -91.120 ;
        RECT -46.735 -90.950 -46.565 -90.880 ;
        RECT -45.795 -90.950 -45.625 -90.880 ;
        RECT -46.735 -91.120 -45.625 -90.950 ;
        RECT -46.735 -91.405 -46.565 -91.120 ;
        RECT -55.715 -91.735 -54.785 -91.405 ;
        RECT -47.495 -91.735 -46.565 -91.405 ;
        RECT -55.715 -92.260 -55.545 -91.735 ;
        RECT -46.735 -92.260 -46.565 -91.735 ;
        RECT -46.325 -92.285 -46.035 -91.120 ;
        RECT -45.795 -91.405 -45.625 -91.120 ;
        RECT -36.815 -90.950 -36.645 -90.880 ;
        RECT -35.875 -90.950 -35.705 -90.880 ;
        RECT -36.815 -91.120 -35.705 -90.950 ;
        RECT -36.815 -91.405 -36.645 -91.120 ;
        RECT -45.795 -91.735 -44.865 -91.405 ;
        RECT -37.575 -91.735 -36.645 -91.405 ;
        RECT -45.795 -92.260 -45.625 -91.735 ;
        RECT -36.815 -92.260 -36.645 -91.735 ;
        RECT -36.405 -92.285 -36.115 -91.120 ;
        RECT -35.875 -91.405 -35.705 -91.120 ;
        RECT -26.895 -90.950 -26.725 -90.880 ;
        RECT -25.955 -90.950 -25.785 -90.880 ;
        RECT -26.895 -91.120 -25.785 -90.950 ;
        RECT -26.895 -91.405 -26.725 -91.120 ;
        RECT -35.875 -91.735 -34.945 -91.405 ;
        RECT -27.655 -91.735 -26.725 -91.405 ;
        RECT -35.875 -92.260 -35.705 -91.735 ;
        RECT -26.895 -92.260 -26.725 -91.735 ;
        RECT -26.485 -92.285 -26.195 -91.120 ;
        RECT -25.955 -91.405 -25.785 -91.120 ;
        RECT -16.975 -90.950 -16.805 -90.880 ;
        RECT -16.035 -90.950 -15.865 -90.880 ;
        RECT -16.975 -91.120 -15.865 -90.950 ;
        RECT -16.975 -91.405 -16.805 -91.120 ;
        RECT -25.955 -91.735 -25.025 -91.405 ;
        RECT -17.735 -91.735 -16.805 -91.405 ;
        RECT -25.955 -92.260 -25.785 -91.735 ;
        RECT -16.975 -92.260 -16.805 -91.735 ;
        RECT -16.565 -92.285 -16.275 -91.120 ;
        RECT -16.035 -91.405 -15.865 -91.120 ;
        RECT -7.055 -90.950 -6.885 -90.880 ;
        RECT -6.115 -90.950 -5.945 -90.880 ;
        RECT -7.055 -91.120 -5.945 -90.950 ;
        RECT -7.055 -91.405 -6.885 -91.120 ;
        RECT -16.035 -91.735 -15.105 -91.405 ;
        RECT -7.815 -91.735 -6.885 -91.405 ;
        RECT -16.035 -92.260 -15.865 -91.735 ;
        RECT -7.055 -92.260 -6.885 -91.735 ;
        RECT -6.645 -92.285 -6.355 -91.120 ;
        RECT -6.115 -91.405 -5.945 -91.120 ;
        RECT 2.865 -90.950 3.035 -90.880 ;
        RECT 3.805 -90.950 3.975 -90.880 ;
        RECT 2.865 -91.120 3.975 -90.950 ;
        RECT 2.865 -91.405 3.035 -91.120 ;
        RECT -6.115 -91.735 -5.185 -91.405 ;
        RECT 2.105 -91.735 3.035 -91.405 ;
        RECT -6.115 -92.260 -5.945 -91.735 ;
        RECT 2.865 -92.260 3.035 -91.735 ;
        RECT 3.275 -92.285 3.565 -91.120 ;
        RECT 3.805 -91.405 3.975 -91.120 ;
        RECT 12.785 -90.950 12.955 -90.880 ;
        RECT 13.725 -90.950 13.895 -90.880 ;
        RECT 12.785 -91.120 13.895 -90.950 ;
        RECT 12.785 -91.405 12.955 -91.120 ;
        RECT 3.805 -91.735 4.735 -91.405 ;
        RECT 12.025 -91.735 12.955 -91.405 ;
        RECT 3.805 -92.260 3.975 -91.735 ;
        RECT 12.785 -92.260 12.955 -91.735 ;
        RECT 13.195 -92.285 13.485 -91.120 ;
        RECT 13.725 -91.405 13.895 -91.120 ;
        RECT 22.705 -90.950 22.875 -90.880 ;
        RECT 23.645 -90.950 23.815 -90.880 ;
        RECT 22.705 -91.120 23.815 -90.950 ;
        RECT 22.705 -91.405 22.875 -91.120 ;
        RECT 13.725 -91.735 14.655 -91.405 ;
        RECT 21.945 -91.735 22.875 -91.405 ;
        RECT 13.725 -92.260 13.895 -91.735 ;
        RECT 22.705 -92.260 22.875 -91.735 ;
        RECT 23.115 -92.285 23.405 -91.120 ;
        RECT 23.645 -91.405 23.815 -91.120 ;
        RECT 23.645 -91.735 24.575 -91.405 ;
        RECT 23.645 -92.260 23.815 -91.735 ;
        RECT -279.605 -173.780 -279.435 -173.630 ;
        RECT -278.665 -173.780 -278.495 -173.630 ;
        RECT -279.605 -173.950 -278.495 -173.780 ;
        RECT -279.605 -174.155 -279.435 -173.950 ;
        RECT -280.365 -174.485 -279.435 -174.155 ;
        RECT -279.605 -175.010 -279.435 -174.485 ;
        RECT -279.195 -175.115 -278.905 -173.950 ;
        RECT -278.665 -174.155 -278.495 -173.950 ;
        RECT -269.685 -173.780 -269.515 -173.630 ;
        RECT -268.745 -173.780 -268.575 -173.630 ;
        RECT -269.685 -173.950 -268.575 -173.780 ;
        RECT -269.685 -174.155 -269.515 -173.950 ;
        RECT -278.665 -174.485 -277.735 -174.155 ;
        RECT -270.445 -174.485 -269.515 -174.155 ;
        RECT -278.665 -175.010 -278.495 -174.485 ;
        RECT -269.685 -175.010 -269.515 -174.485 ;
        RECT -269.275 -175.115 -268.985 -173.950 ;
        RECT -268.745 -174.155 -268.575 -173.950 ;
        RECT -259.765 -173.780 -259.595 -173.630 ;
        RECT -258.825 -173.780 -258.655 -173.630 ;
        RECT -259.765 -173.950 -258.655 -173.780 ;
        RECT -259.765 -174.155 -259.595 -173.950 ;
        RECT -268.745 -174.485 -267.815 -174.155 ;
        RECT -260.525 -174.485 -259.595 -174.155 ;
        RECT -268.745 -175.010 -268.575 -174.485 ;
        RECT -259.765 -175.010 -259.595 -174.485 ;
        RECT -259.355 -175.115 -259.065 -173.950 ;
        RECT -258.825 -174.155 -258.655 -173.950 ;
        RECT -249.845 -173.780 -249.675 -173.630 ;
        RECT -248.905 -173.780 -248.735 -173.630 ;
        RECT -249.845 -173.950 -248.735 -173.780 ;
        RECT -249.845 -174.155 -249.675 -173.950 ;
        RECT -258.825 -174.485 -257.895 -174.155 ;
        RECT -250.605 -174.485 -249.675 -174.155 ;
        RECT -258.825 -175.010 -258.655 -174.485 ;
        RECT -249.845 -175.010 -249.675 -174.485 ;
        RECT -249.435 -175.115 -249.145 -173.950 ;
        RECT -248.905 -174.155 -248.735 -173.950 ;
        RECT -239.925 -173.780 -239.755 -173.630 ;
        RECT -238.985 -173.780 -238.815 -173.630 ;
        RECT -239.925 -173.950 -238.815 -173.780 ;
        RECT -239.925 -174.155 -239.755 -173.950 ;
        RECT -248.905 -174.485 -247.975 -174.155 ;
        RECT -240.685 -174.485 -239.755 -174.155 ;
        RECT -248.905 -175.010 -248.735 -174.485 ;
        RECT -239.925 -175.010 -239.755 -174.485 ;
        RECT -239.515 -175.115 -239.225 -173.950 ;
        RECT -238.985 -174.155 -238.815 -173.950 ;
        RECT -230.005 -173.780 -229.835 -173.630 ;
        RECT -229.065 -173.780 -228.895 -173.630 ;
        RECT -230.005 -173.950 -228.895 -173.780 ;
        RECT -230.005 -174.155 -229.835 -173.950 ;
        RECT -238.985 -174.485 -238.055 -174.155 ;
        RECT -230.765 -174.485 -229.835 -174.155 ;
        RECT -238.985 -175.010 -238.815 -174.485 ;
        RECT -230.005 -175.010 -229.835 -174.485 ;
        RECT -229.595 -175.115 -229.305 -173.950 ;
        RECT -229.065 -174.155 -228.895 -173.950 ;
        RECT -220.085 -173.780 -219.915 -173.630 ;
        RECT -219.145 -173.780 -218.975 -173.630 ;
        RECT -220.085 -173.950 -218.975 -173.780 ;
        RECT -220.085 -174.155 -219.915 -173.950 ;
        RECT -229.065 -174.485 -228.135 -174.155 ;
        RECT -220.845 -174.485 -219.915 -174.155 ;
        RECT -229.065 -175.010 -228.895 -174.485 ;
        RECT -220.085 -175.010 -219.915 -174.485 ;
        RECT -219.675 -175.115 -219.385 -173.950 ;
        RECT -219.145 -174.155 -218.975 -173.950 ;
        RECT -210.165 -173.780 -209.995 -173.630 ;
        RECT -209.225 -173.780 -209.055 -173.630 ;
        RECT -210.165 -173.950 -209.055 -173.780 ;
        RECT -210.165 -174.155 -209.995 -173.950 ;
        RECT -219.145 -174.485 -218.215 -174.155 ;
        RECT -210.925 -174.485 -209.995 -174.155 ;
        RECT -219.145 -175.010 -218.975 -174.485 ;
        RECT -210.165 -175.010 -209.995 -174.485 ;
        RECT -209.755 -175.115 -209.465 -173.950 ;
        RECT -209.225 -174.155 -209.055 -173.950 ;
        RECT -200.245 -173.780 -200.075 -173.630 ;
        RECT -199.305 -173.780 -199.135 -173.630 ;
        RECT -200.245 -173.950 -199.135 -173.780 ;
        RECT -200.245 -174.155 -200.075 -173.950 ;
        RECT -209.225 -174.485 -208.295 -174.155 ;
        RECT -201.005 -174.485 -200.075 -174.155 ;
        RECT -209.225 -175.010 -209.055 -174.485 ;
        RECT -200.245 -175.010 -200.075 -174.485 ;
        RECT -199.835 -175.115 -199.545 -173.950 ;
        RECT -199.305 -174.155 -199.135 -173.950 ;
        RECT -190.325 -173.780 -190.155 -173.630 ;
        RECT -189.385 -173.780 -189.215 -173.630 ;
        RECT -190.325 -173.950 -189.215 -173.780 ;
        RECT -190.325 -174.155 -190.155 -173.950 ;
        RECT -199.305 -174.485 -198.375 -174.155 ;
        RECT -191.085 -174.485 -190.155 -174.155 ;
        RECT -199.305 -175.010 -199.135 -174.485 ;
        RECT -190.325 -175.010 -190.155 -174.485 ;
        RECT -189.915 -175.115 -189.625 -173.950 ;
        RECT -189.385 -174.155 -189.215 -173.950 ;
        RECT -180.405 -173.780 -180.235 -173.630 ;
        RECT -179.465 -173.780 -179.295 -173.630 ;
        RECT -180.405 -173.950 -179.295 -173.780 ;
        RECT -180.405 -174.155 -180.235 -173.950 ;
        RECT -189.385 -174.485 -188.455 -174.155 ;
        RECT -181.165 -174.485 -180.235 -174.155 ;
        RECT -189.385 -175.010 -189.215 -174.485 ;
        RECT -180.405 -175.010 -180.235 -174.485 ;
        RECT -179.995 -175.115 -179.705 -173.950 ;
        RECT -179.465 -174.155 -179.295 -173.950 ;
        RECT -170.485 -173.780 -170.315 -173.630 ;
        RECT -169.545 -173.780 -169.375 -173.630 ;
        RECT -170.485 -173.950 -169.375 -173.780 ;
        RECT -170.485 -174.155 -170.315 -173.950 ;
        RECT -179.465 -174.485 -178.535 -174.155 ;
        RECT -171.245 -174.485 -170.315 -174.155 ;
        RECT -179.465 -175.010 -179.295 -174.485 ;
        RECT -170.485 -175.010 -170.315 -174.485 ;
        RECT -170.075 -175.115 -169.785 -173.950 ;
        RECT -169.545 -174.155 -169.375 -173.950 ;
        RECT -160.565 -173.780 -160.395 -173.630 ;
        RECT -159.625 -173.780 -159.455 -173.630 ;
        RECT -160.565 -173.950 -159.455 -173.780 ;
        RECT -160.565 -174.155 -160.395 -173.950 ;
        RECT -169.545 -174.485 -168.615 -174.155 ;
        RECT -161.325 -174.485 -160.395 -174.155 ;
        RECT -169.545 -175.010 -169.375 -174.485 ;
        RECT -160.565 -175.010 -160.395 -174.485 ;
        RECT -160.155 -175.115 -159.865 -173.950 ;
        RECT -159.625 -174.155 -159.455 -173.950 ;
        RECT -150.645 -173.780 -150.475 -173.630 ;
        RECT -149.705 -173.780 -149.535 -173.630 ;
        RECT -150.645 -173.950 -149.535 -173.780 ;
        RECT -150.645 -174.155 -150.475 -173.950 ;
        RECT -159.625 -174.485 -158.695 -174.155 ;
        RECT -151.405 -174.485 -150.475 -174.155 ;
        RECT -159.625 -175.010 -159.455 -174.485 ;
        RECT -150.645 -175.010 -150.475 -174.485 ;
        RECT -150.235 -175.115 -149.945 -173.950 ;
        RECT -149.705 -174.155 -149.535 -173.950 ;
        RECT -140.725 -173.780 -140.555 -173.630 ;
        RECT -139.785 -173.780 -139.615 -173.630 ;
        RECT -140.725 -173.950 -139.615 -173.780 ;
        RECT -140.725 -174.155 -140.555 -173.950 ;
        RECT -149.705 -174.485 -148.775 -174.155 ;
        RECT -141.485 -174.485 -140.555 -174.155 ;
        RECT -149.705 -175.010 -149.535 -174.485 ;
        RECT -140.725 -175.010 -140.555 -174.485 ;
        RECT -140.315 -175.115 -140.025 -173.950 ;
        RECT -139.785 -174.155 -139.615 -173.950 ;
        RECT -130.805 -173.780 -130.635 -173.630 ;
        RECT -129.865 -173.780 -129.695 -173.630 ;
        RECT -130.805 -173.950 -129.695 -173.780 ;
        RECT -130.805 -174.155 -130.635 -173.950 ;
        RECT -139.785 -174.485 -138.855 -174.155 ;
        RECT -131.565 -174.485 -130.635 -174.155 ;
        RECT -139.785 -175.010 -139.615 -174.485 ;
        RECT -130.805 -175.010 -130.635 -174.485 ;
        RECT -130.395 -175.115 -130.105 -173.950 ;
        RECT -129.865 -174.155 -129.695 -173.950 ;
        RECT -120.885 -173.780 -120.715 -173.630 ;
        RECT -119.945 -173.780 -119.775 -173.630 ;
        RECT -120.885 -173.950 -119.775 -173.780 ;
        RECT -120.885 -174.155 -120.715 -173.950 ;
        RECT -129.865 -174.485 -128.935 -174.155 ;
        RECT -121.645 -174.485 -120.715 -174.155 ;
        RECT -129.865 -175.010 -129.695 -174.485 ;
        RECT -120.885 -175.010 -120.715 -174.485 ;
        RECT -120.475 -175.115 -120.185 -173.950 ;
        RECT -119.945 -174.155 -119.775 -173.950 ;
        RECT -110.965 -173.780 -110.795 -173.630 ;
        RECT -110.025 -173.780 -109.855 -173.630 ;
        RECT -110.965 -173.950 -109.855 -173.780 ;
        RECT -110.965 -174.155 -110.795 -173.950 ;
        RECT -119.945 -174.485 -119.015 -174.155 ;
        RECT -111.725 -174.485 -110.795 -174.155 ;
        RECT -119.945 -175.010 -119.775 -174.485 ;
        RECT -110.965 -175.010 -110.795 -174.485 ;
        RECT -110.555 -175.115 -110.265 -173.950 ;
        RECT -110.025 -174.155 -109.855 -173.950 ;
        RECT -101.045 -173.780 -100.875 -173.630 ;
        RECT -100.105 -173.780 -99.935 -173.630 ;
        RECT -101.045 -173.950 -99.935 -173.780 ;
        RECT -101.045 -174.155 -100.875 -173.950 ;
        RECT -110.025 -174.485 -109.095 -174.155 ;
        RECT -101.805 -174.485 -100.875 -174.155 ;
        RECT -110.025 -175.010 -109.855 -174.485 ;
        RECT -101.045 -175.010 -100.875 -174.485 ;
        RECT -100.635 -175.115 -100.345 -173.950 ;
        RECT -100.105 -174.155 -99.935 -173.950 ;
        RECT -91.125 -173.780 -90.955 -173.630 ;
        RECT -90.185 -173.780 -90.015 -173.630 ;
        RECT -91.125 -173.950 -90.015 -173.780 ;
        RECT -91.125 -174.155 -90.955 -173.950 ;
        RECT -100.105 -174.485 -99.175 -174.155 ;
        RECT -91.885 -174.485 -90.955 -174.155 ;
        RECT -100.105 -175.010 -99.935 -174.485 ;
        RECT -91.125 -175.010 -90.955 -174.485 ;
        RECT -90.715 -175.115 -90.425 -173.950 ;
        RECT -90.185 -174.155 -90.015 -173.950 ;
        RECT -81.205 -173.780 -81.035 -173.630 ;
        RECT -80.265 -173.780 -80.095 -173.630 ;
        RECT -81.205 -173.950 -80.095 -173.780 ;
        RECT -81.205 -174.155 -81.035 -173.950 ;
        RECT -90.185 -174.485 -89.255 -174.155 ;
        RECT -81.965 -174.485 -81.035 -174.155 ;
        RECT -90.185 -175.010 -90.015 -174.485 ;
        RECT -81.205 -175.010 -81.035 -174.485 ;
        RECT -80.795 -175.115 -80.505 -173.950 ;
        RECT -80.265 -174.155 -80.095 -173.950 ;
        RECT -71.285 -173.780 -71.115 -173.630 ;
        RECT -70.345 -173.780 -70.175 -173.630 ;
        RECT -71.285 -173.950 -70.175 -173.780 ;
        RECT -71.285 -174.155 -71.115 -173.950 ;
        RECT -80.265 -174.485 -79.335 -174.155 ;
        RECT -72.045 -174.485 -71.115 -174.155 ;
        RECT -80.265 -175.010 -80.095 -174.485 ;
        RECT -71.285 -175.010 -71.115 -174.485 ;
        RECT -70.875 -175.115 -70.585 -173.950 ;
        RECT -70.345 -174.155 -70.175 -173.950 ;
        RECT -61.365 -173.780 -61.195 -173.630 ;
        RECT -60.425 -173.780 -60.255 -173.630 ;
        RECT -61.365 -173.950 -60.255 -173.780 ;
        RECT -61.365 -174.155 -61.195 -173.950 ;
        RECT -70.345 -174.485 -69.415 -174.155 ;
        RECT -62.125 -174.485 -61.195 -174.155 ;
        RECT -70.345 -175.010 -70.175 -174.485 ;
        RECT -61.365 -175.010 -61.195 -174.485 ;
        RECT -60.955 -175.115 -60.665 -173.950 ;
        RECT -60.425 -174.155 -60.255 -173.950 ;
        RECT -51.445 -173.780 -51.275 -173.630 ;
        RECT -50.505 -173.780 -50.335 -173.630 ;
        RECT -51.445 -173.950 -50.335 -173.780 ;
        RECT -51.445 -174.155 -51.275 -173.950 ;
        RECT -60.425 -174.485 -59.495 -174.155 ;
        RECT -52.205 -174.485 -51.275 -174.155 ;
        RECT -60.425 -175.010 -60.255 -174.485 ;
        RECT -51.445 -175.010 -51.275 -174.485 ;
        RECT -51.035 -175.115 -50.745 -173.950 ;
        RECT -50.505 -174.155 -50.335 -173.950 ;
        RECT -41.525 -173.780 -41.355 -173.630 ;
        RECT -40.585 -173.780 -40.415 -173.630 ;
        RECT -41.525 -173.950 -40.415 -173.780 ;
        RECT -41.525 -174.155 -41.355 -173.950 ;
        RECT -50.505 -174.485 -49.575 -174.155 ;
        RECT -42.285 -174.485 -41.355 -174.155 ;
        RECT -50.505 -175.010 -50.335 -174.485 ;
        RECT -41.525 -175.010 -41.355 -174.485 ;
        RECT -41.115 -175.115 -40.825 -173.950 ;
        RECT -40.585 -174.155 -40.415 -173.950 ;
        RECT -31.605 -173.780 -31.435 -173.630 ;
        RECT -30.665 -173.780 -30.495 -173.630 ;
        RECT -31.605 -173.950 -30.495 -173.780 ;
        RECT -31.605 -174.155 -31.435 -173.950 ;
        RECT -40.585 -174.485 -39.655 -174.155 ;
        RECT -32.365 -174.485 -31.435 -174.155 ;
        RECT -40.585 -175.010 -40.415 -174.485 ;
        RECT -31.605 -175.010 -31.435 -174.485 ;
        RECT -31.195 -175.115 -30.905 -173.950 ;
        RECT -30.665 -174.155 -30.495 -173.950 ;
        RECT -21.685 -173.780 -21.515 -173.630 ;
        RECT -20.745 -173.780 -20.575 -173.630 ;
        RECT -21.685 -173.950 -20.575 -173.780 ;
        RECT -21.685 -174.155 -21.515 -173.950 ;
        RECT -30.665 -174.485 -29.735 -174.155 ;
        RECT -22.445 -174.485 -21.515 -174.155 ;
        RECT -30.665 -175.010 -30.495 -174.485 ;
        RECT -21.685 -175.010 -21.515 -174.485 ;
        RECT -21.275 -175.115 -20.985 -173.950 ;
        RECT -20.745 -174.155 -20.575 -173.950 ;
        RECT -11.765 -173.780 -11.595 -173.630 ;
        RECT -10.825 -173.780 -10.655 -173.630 ;
        RECT -11.765 -173.950 -10.655 -173.780 ;
        RECT -11.765 -174.155 -11.595 -173.950 ;
        RECT -20.745 -174.485 -19.815 -174.155 ;
        RECT -12.525 -174.485 -11.595 -174.155 ;
        RECT -20.745 -175.010 -20.575 -174.485 ;
        RECT -11.765 -175.010 -11.595 -174.485 ;
        RECT -11.355 -175.115 -11.065 -173.950 ;
        RECT -10.825 -174.155 -10.655 -173.950 ;
        RECT -1.845 -173.780 -1.675 -173.630 ;
        RECT -0.905 -173.780 -0.735 -173.630 ;
        RECT -1.845 -173.950 -0.735 -173.780 ;
        RECT -1.845 -174.155 -1.675 -173.950 ;
        RECT -10.825 -174.485 -9.895 -174.155 ;
        RECT -2.605 -174.485 -1.675 -174.155 ;
        RECT -10.825 -175.010 -10.655 -174.485 ;
        RECT -1.845 -175.010 -1.675 -174.485 ;
        RECT -1.435 -175.115 -1.145 -173.950 ;
        RECT -0.905 -174.155 -0.735 -173.950 ;
        RECT 8.075 -173.780 8.245 -173.630 ;
        RECT 9.015 -173.780 9.185 -173.630 ;
        RECT 8.075 -173.950 9.185 -173.780 ;
        RECT 8.075 -174.155 8.245 -173.950 ;
        RECT -0.905 -174.485 0.025 -174.155 ;
        RECT 7.315 -174.485 8.245 -174.155 ;
        RECT -0.905 -175.010 -0.735 -174.485 ;
        RECT 8.075 -175.010 8.245 -174.485 ;
        RECT 8.485 -175.115 8.775 -173.950 ;
        RECT 9.015 -174.155 9.185 -173.950 ;
        RECT 17.995 -173.780 18.165 -173.630 ;
        RECT 18.935 -173.780 19.105 -173.630 ;
        RECT 17.995 -173.950 19.105 -173.780 ;
        RECT 17.995 -174.155 18.165 -173.950 ;
        RECT 9.015 -174.485 9.945 -174.155 ;
        RECT 17.235 -174.485 18.165 -174.155 ;
        RECT 9.015 -175.010 9.185 -174.485 ;
        RECT 17.995 -175.010 18.165 -174.485 ;
        RECT 18.405 -175.115 18.695 -173.950 ;
        RECT 18.935 -174.155 19.105 -173.950 ;
        RECT 27.915 -173.780 28.085 -173.630 ;
        RECT 27.915 -173.950 28.700 -173.780 ;
        RECT 27.915 -174.155 28.085 -173.950 ;
        RECT 18.935 -174.485 19.865 -174.155 ;
        RECT 27.155 -174.485 28.085 -174.155 ;
        RECT 18.935 -175.010 19.105 -174.485 ;
        RECT 27.915 -175.010 28.085 -174.485 ;
        RECT 28.325 -175.115 28.615 -173.950 ;
        RECT -285.620 -175.525 -282.400 -175.355 ;
        RECT -275.700 -175.525 -272.480 -175.355 ;
        RECT -265.780 -175.525 -262.560 -175.355 ;
        RECT -255.860 -175.525 -252.640 -175.355 ;
        RECT -245.940 -175.525 -242.720 -175.355 ;
        RECT -236.020 -175.525 -232.800 -175.355 ;
        RECT -226.100 -175.525 -222.880 -175.355 ;
        RECT -216.180 -175.525 -212.960 -175.355 ;
        RECT -206.260 -175.525 -203.040 -175.355 ;
        RECT -196.340 -175.525 -193.120 -175.355 ;
        RECT -186.420 -175.525 -183.200 -175.355 ;
        RECT -176.500 -175.525 -173.280 -175.355 ;
        RECT -166.580 -175.525 -163.360 -175.355 ;
        RECT -156.660 -175.525 -153.440 -175.355 ;
        RECT -146.740 -175.525 -143.520 -175.355 ;
        RECT -136.820 -175.525 -133.600 -175.355 ;
        RECT -126.900 -175.525 -123.680 -175.355 ;
        RECT -116.980 -175.525 -113.760 -175.355 ;
        RECT -107.060 -175.525 -103.840 -175.355 ;
        RECT -97.140 -175.525 -93.920 -175.355 ;
        RECT -87.220 -175.525 -84.000 -175.355 ;
        RECT -77.300 -175.525 -74.080 -175.355 ;
        RECT -67.380 -175.525 -64.160 -175.355 ;
        RECT -57.460 -175.525 -54.240 -175.355 ;
        RECT -47.540 -175.525 -44.320 -175.355 ;
        RECT -37.620 -175.525 -34.400 -175.355 ;
        RECT -27.700 -175.525 -24.480 -175.355 ;
        RECT -17.780 -175.525 -14.560 -175.355 ;
        RECT -7.860 -175.525 -4.640 -175.355 ;
        RECT 2.060 -175.525 5.280 -175.355 ;
        RECT 11.980 -175.525 15.200 -175.355 ;
        RECT 21.900 -175.525 25.120 -175.355 ;
        RECT -285.535 -176.665 -285.275 -175.525 ;
        RECT -284.605 -176.665 -284.325 -175.525 ;
        RECT -284.155 -176.690 -283.865 -175.525 ;
        RECT -283.695 -176.665 -283.415 -175.525 ;
        RECT -282.745 -176.665 -282.485 -175.525 ;
        RECT -275.615 -176.665 -275.355 -175.525 ;
        RECT -274.685 -176.665 -274.405 -175.525 ;
        RECT -274.235 -176.690 -273.945 -175.525 ;
        RECT -273.775 -176.665 -273.495 -175.525 ;
        RECT -272.825 -176.665 -272.565 -175.525 ;
        RECT -265.695 -176.665 -265.435 -175.525 ;
        RECT -264.765 -176.665 -264.485 -175.525 ;
        RECT -264.315 -176.690 -264.025 -175.525 ;
        RECT -263.855 -176.665 -263.575 -175.525 ;
        RECT -262.905 -176.665 -262.645 -175.525 ;
        RECT -255.775 -176.665 -255.515 -175.525 ;
        RECT -254.845 -176.665 -254.565 -175.525 ;
        RECT -254.395 -176.690 -254.105 -175.525 ;
        RECT -253.935 -176.665 -253.655 -175.525 ;
        RECT -252.985 -176.665 -252.725 -175.525 ;
        RECT -245.855 -176.665 -245.595 -175.525 ;
        RECT -244.925 -176.665 -244.645 -175.525 ;
        RECT -244.475 -176.690 -244.185 -175.525 ;
        RECT -244.015 -176.665 -243.735 -175.525 ;
        RECT -243.065 -176.665 -242.805 -175.525 ;
        RECT -235.935 -176.665 -235.675 -175.525 ;
        RECT -235.005 -176.665 -234.725 -175.525 ;
        RECT -234.555 -176.690 -234.265 -175.525 ;
        RECT -234.095 -176.665 -233.815 -175.525 ;
        RECT -233.145 -176.665 -232.885 -175.525 ;
        RECT -226.015 -176.665 -225.755 -175.525 ;
        RECT -225.085 -176.665 -224.805 -175.525 ;
        RECT -224.635 -176.690 -224.345 -175.525 ;
        RECT -224.175 -176.665 -223.895 -175.525 ;
        RECT -223.225 -176.665 -222.965 -175.525 ;
        RECT -216.095 -176.665 -215.835 -175.525 ;
        RECT -215.165 -176.665 -214.885 -175.525 ;
        RECT -214.715 -176.690 -214.425 -175.525 ;
        RECT -214.255 -176.665 -213.975 -175.525 ;
        RECT -213.305 -176.665 -213.045 -175.525 ;
        RECT -206.175 -176.665 -205.915 -175.525 ;
        RECT -205.245 -176.665 -204.965 -175.525 ;
        RECT -204.795 -176.690 -204.505 -175.525 ;
        RECT -204.335 -176.665 -204.055 -175.525 ;
        RECT -203.385 -176.665 -203.125 -175.525 ;
        RECT -196.255 -176.665 -195.995 -175.525 ;
        RECT -195.325 -176.665 -195.045 -175.525 ;
        RECT -194.875 -176.690 -194.585 -175.525 ;
        RECT -194.415 -176.665 -194.135 -175.525 ;
        RECT -193.465 -176.665 -193.205 -175.525 ;
        RECT -186.335 -176.665 -186.075 -175.525 ;
        RECT -185.405 -176.665 -185.125 -175.525 ;
        RECT -184.955 -176.690 -184.665 -175.525 ;
        RECT -184.495 -176.665 -184.215 -175.525 ;
        RECT -183.545 -176.665 -183.285 -175.525 ;
        RECT -176.415 -176.665 -176.155 -175.525 ;
        RECT -175.485 -176.665 -175.205 -175.525 ;
        RECT -175.035 -176.690 -174.745 -175.525 ;
        RECT -174.575 -176.665 -174.295 -175.525 ;
        RECT -173.625 -176.665 -173.365 -175.525 ;
        RECT -166.495 -176.665 -166.235 -175.525 ;
        RECT -165.565 -176.665 -165.285 -175.525 ;
        RECT -165.115 -176.690 -164.825 -175.525 ;
        RECT -164.655 -176.665 -164.375 -175.525 ;
        RECT -163.705 -176.665 -163.445 -175.525 ;
        RECT -156.575 -176.665 -156.315 -175.525 ;
        RECT -155.645 -176.665 -155.365 -175.525 ;
        RECT -155.195 -176.690 -154.905 -175.525 ;
        RECT -154.735 -176.665 -154.455 -175.525 ;
        RECT -153.785 -176.665 -153.525 -175.525 ;
        RECT -146.655 -176.665 -146.395 -175.525 ;
        RECT -145.725 -176.665 -145.445 -175.525 ;
        RECT -145.275 -176.690 -144.985 -175.525 ;
        RECT -144.815 -176.665 -144.535 -175.525 ;
        RECT -143.865 -176.665 -143.605 -175.525 ;
        RECT -136.735 -176.665 -136.475 -175.525 ;
        RECT -135.805 -176.665 -135.525 -175.525 ;
        RECT -135.355 -176.690 -135.065 -175.525 ;
        RECT -134.895 -176.665 -134.615 -175.525 ;
        RECT -133.945 -176.665 -133.685 -175.525 ;
        RECT -126.815 -176.665 -126.555 -175.525 ;
        RECT -125.885 -176.665 -125.605 -175.525 ;
        RECT -125.435 -176.690 -125.145 -175.525 ;
        RECT -124.975 -176.665 -124.695 -175.525 ;
        RECT -124.025 -176.665 -123.765 -175.525 ;
        RECT -116.895 -176.665 -116.635 -175.525 ;
        RECT -115.965 -176.665 -115.685 -175.525 ;
        RECT -115.515 -176.690 -115.225 -175.525 ;
        RECT -115.055 -176.665 -114.775 -175.525 ;
        RECT -114.105 -176.665 -113.845 -175.525 ;
        RECT -106.975 -176.665 -106.715 -175.525 ;
        RECT -106.045 -176.665 -105.765 -175.525 ;
        RECT -105.595 -176.690 -105.305 -175.525 ;
        RECT -105.135 -176.665 -104.855 -175.525 ;
        RECT -104.185 -176.665 -103.925 -175.525 ;
        RECT -97.055 -176.665 -96.795 -175.525 ;
        RECT -96.125 -176.665 -95.845 -175.525 ;
        RECT -95.675 -176.690 -95.385 -175.525 ;
        RECT -95.215 -176.665 -94.935 -175.525 ;
        RECT -94.265 -176.665 -94.005 -175.525 ;
        RECT -87.135 -176.665 -86.875 -175.525 ;
        RECT -86.205 -176.665 -85.925 -175.525 ;
        RECT -85.755 -176.690 -85.465 -175.525 ;
        RECT -85.295 -176.665 -85.015 -175.525 ;
        RECT -84.345 -176.665 -84.085 -175.525 ;
        RECT -77.215 -176.665 -76.955 -175.525 ;
        RECT -76.285 -176.665 -76.005 -175.525 ;
        RECT -75.835 -176.690 -75.545 -175.525 ;
        RECT -75.375 -176.665 -75.095 -175.525 ;
        RECT -74.425 -176.665 -74.165 -175.525 ;
        RECT -67.295 -176.665 -67.035 -175.525 ;
        RECT -66.365 -176.665 -66.085 -175.525 ;
        RECT -65.915 -176.690 -65.625 -175.525 ;
        RECT -65.455 -176.665 -65.175 -175.525 ;
        RECT -64.505 -176.665 -64.245 -175.525 ;
        RECT -57.375 -176.665 -57.115 -175.525 ;
        RECT -56.445 -176.665 -56.165 -175.525 ;
        RECT -55.995 -176.690 -55.705 -175.525 ;
        RECT -55.535 -176.665 -55.255 -175.525 ;
        RECT -54.585 -176.665 -54.325 -175.525 ;
        RECT -47.455 -176.665 -47.195 -175.525 ;
        RECT -46.525 -176.665 -46.245 -175.525 ;
        RECT -46.075 -176.690 -45.785 -175.525 ;
        RECT -45.615 -176.665 -45.335 -175.525 ;
        RECT -44.665 -176.665 -44.405 -175.525 ;
        RECT -37.535 -176.665 -37.275 -175.525 ;
        RECT -36.605 -176.665 -36.325 -175.525 ;
        RECT -36.155 -176.690 -35.865 -175.525 ;
        RECT -35.695 -176.665 -35.415 -175.525 ;
        RECT -34.745 -176.665 -34.485 -175.525 ;
        RECT -27.615 -176.665 -27.355 -175.525 ;
        RECT -26.685 -176.665 -26.405 -175.525 ;
        RECT -26.235 -176.690 -25.945 -175.525 ;
        RECT -25.775 -176.665 -25.495 -175.525 ;
        RECT -24.825 -176.665 -24.565 -175.525 ;
        RECT -17.695 -176.665 -17.435 -175.525 ;
        RECT -16.765 -176.665 -16.485 -175.525 ;
        RECT -16.315 -176.690 -16.025 -175.525 ;
        RECT -15.855 -176.665 -15.575 -175.525 ;
        RECT -14.905 -176.665 -14.645 -175.525 ;
        RECT -7.775 -176.665 -7.515 -175.525 ;
        RECT -6.845 -176.665 -6.565 -175.525 ;
        RECT -6.395 -176.690 -6.105 -175.525 ;
        RECT -5.935 -176.665 -5.655 -175.525 ;
        RECT -4.985 -176.665 -4.725 -175.525 ;
        RECT 2.145 -176.665 2.405 -175.525 ;
        RECT 3.075 -176.665 3.355 -175.525 ;
        RECT 3.525 -176.690 3.815 -175.525 ;
        RECT 3.985 -176.665 4.265 -175.525 ;
        RECT 4.935 -176.665 5.195 -175.525 ;
        RECT 12.065 -176.665 12.325 -175.525 ;
        RECT 12.995 -176.665 13.275 -175.525 ;
        RECT 13.445 -176.690 13.735 -175.525 ;
        RECT 13.905 -176.665 14.185 -175.525 ;
        RECT 14.855 -176.665 15.115 -175.525 ;
        RECT 21.985 -176.665 22.245 -175.525 ;
        RECT 22.915 -176.665 23.195 -175.525 ;
        RECT 23.365 -176.690 23.655 -175.525 ;
        RECT 23.825 -176.665 24.105 -175.525 ;
        RECT 24.775 -176.665 25.035 -175.525 ;
        RECT -280.575 -178.075 -280.315 -176.935 ;
        RECT -279.645 -178.075 -279.365 -176.935 ;
        RECT -279.195 -178.075 -278.905 -176.910 ;
        RECT -278.735 -178.075 -278.455 -176.935 ;
        RECT -277.785 -178.075 -277.525 -176.935 ;
        RECT -270.655 -178.075 -270.395 -176.935 ;
        RECT -269.725 -178.075 -269.445 -176.935 ;
        RECT -269.275 -178.075 -268.985 -176.910 ;
        RECT -268.815 -178.075 -268.535 -176.935 ;
        RECT -267.865 -178.075 -267.605 -176.935 ;
        RECT -260.735 -178.075 -260.475 -176.935 ;
        RECT -259.805 -178.075 -259.525 -176.935 ;
        RECT -259.355 -178.075 -259.065 -176.910 ;
        RECT -258.895 -178.075 -258.615 -176.935 ;
        RECT -257.945 -178.075 -257.685 -176.935 ;
        RECT -250.815 -178.075 -250.555 -176.935 ;
        RECT -249.885 -178.075 -249.605 -176.935 ;
        RECT -249.435 -178.075 -249.145 -176.910 ;
        RECT -248.975 -178.075 -248.695 -176.935 ;
        RECT -248.025 -178.075 -247.765 -176.935 ;
        RECT -240.895 -178.075 -240.635 -176.935 ;
        RECT -239.965 -178.075 -239.685 -176.935 ;
        RECT -239.515 -178.075 -239.225 -176.910 ;
        RECT -239.055 -178.075 -238.775 -176.935 ;
        RECT -238.105 -178.075 -237.845 -176.935 ;
        RECT -230.975 -178.075 -230.715 -176.935 ;
        RECT -230.045 -178.075 -229.765 -176.935 ;
        RECT -229.595 -178.075 -229.305 -176.910 ;
        RECT -229.135 -178.075 -228.855 -176.935 ;
        RECT -228.185 -178.075 -227.925 -176.935 ;
        RECT -221.055 -178.075 -220.795 -176.935 ;
        RECT -220.125 -178.075 -219.845 -176.935 ;
        RECT -219.675 -178.075 -219.385 -176.910 ;
        RECT -219.215 -178.075 -218.935 -176.935 ;
        RECT -218.265 -178.075 -218.005 -176.935 ;
        RECT -211.135 -178.075 -210.875 -176.935 ;
        RECT -210.205 -178.075 -209.925 -176.935 ;
        RECT -209.755 -178.075 -209.465 -176.910 ;
        RECT -209.295 -178.075 -209.015 -176.935 ;
        RECT -208.345 -178.075 -208.085 -176.935 ;
        RECT -201.215 -178.075 -200.955 -176.935 ;
        RECT -200.285 -178.075 -200.005 -176.935 ;
        RECT -199.835 -178.075 -199.545 -176.910 ;
        RECT -199.375 -178.075 -199.095 -176.935 ;
        RECT -198.425 -178.075 -198.165 -176.935 ;
        RECT -191.295 -178.075 -191.035 -176.935 ;
        RECT -190.365 -178.075 -190.085 -176.935 ;
        RECT -189.915 -178.075 -189.625 -176.910 ;
        RECT -189.455 -178.075 -189.175 -176.935 ;
        RECT -188.505 -178.075 -188.245 -176.935 ;
        RECT -181.375 -178.075 -181.115 -176.935 ;
        RECT -180.445 -178.075 -180.165 -176.935 ;
        RECT -179.995 -178.075 -179.705 -176.910 ;
        RECT -179.535 -178.075 -179.255 -176.935 ;
        RECT -178.585 -178.075 -178.325 -176.935 ;
        RECT -171.455 -178.075 -171.195 -176.935 ;
        RECT -170.525 -178.075 -170.245 -176.935 ;
        RECT -170.075 -178.075 -169.785 -176.910 ;
        RECT -169.615 -178.075 -169.335 -176.935 ;
        RECT -168.665 -178.075 -168.405 -176.935 ;
        RECT -161.535 -178.075 -161.275 -176.935 ;
        RECT -160.605 -178.075 -160.325 -176.935 ;
        RECT -160.155 -178.075 -159.865 -176.910 ;
        RECT -159.695 -178.075 -159.415 -176.935 ;
        RECT -158.745 -178.075 -158.485 -176.935 ;
        RECT -151.615 -178.075 -151.355 -176.935 ;
        RECT -150.685 -178.075 -150.405 -176.935 ;
        RECT -150.235 -178.075 -149.945 -176.910 ;
        RECT -149.775 -178.075 -149.495 -176.935 ;
        RECT -148.825 -178.075 -148.565 -176.935 ;
        RECT -141.695 -178.075 -141.435 -176.935 ;
        RECT -140.765 -178.075 -140.485 -176.935 ;
        RECT -140.315 -178.075 -140.025 -176.910 ;
        RECT -139.855 -178.075 -139.575 -176.935 ;
        RECT -138.905 -178.075 -138.645 -176.935 ;
        RECT -131.775 -178.075 -131.515 -176.935 ;
        RECT -130.845 -178.075 -130.565 -176.935 ;
        RECT -130.395 -178.075 -130.105 -176.910 ;
        RECT -129.935 -178.075 -129.655 -176.935 ;
        RECT -128.985 -178.075 -128.725 -176.935 ;
        RECT -121.855 -178.075 -121.595 -176.935 ;
        RECT -120.925 -178.075 -120.645 -176.935 ;
        RECT -120.475 -178.075 -120.185 -176.910 ;
        RECT -120.015 -178.075 -119.735 -176.935 ;
        RECT -119.065 -178.075 -118.805 -176.935 ;
        RECT -111.935 -178.075 -111.675 -176.935 ;
        RECT -111.005 -178.075 -110.725 -176.935 ;
        RECT -110.555 -178.075 -110.265 -176.910 ;
        RECT -110.095 -178.075 -109.815 -176.935 ;
        RECT -109.145 -178.075 -108.885 -176.935 ;
        RECT -102.015 -178.075 -101.755 -176.935 ;
        RECT -101.085 -178.075 -100.805 -176.935 ;
        RECT -100.635 -178.075 -100.345 -176.910 ;
        RECT -100.175 -178.075 -99.895 -176.935 ;
        RECT -99.225 -178.075 -98.965 -176.935 ;
        RECT -92.095 -178.075 -91.835 -176.935 ;
        RECT -91.165 -178.075 -90.885 -176.935 ;
        RECT -90.715 -178.075 -90.425 -176.910 ;
        RECT -90.255 -178.075 -89.975 -176.935 ;
        RECT -89.305 -178.075 -89.045 -176.935 ;
        RECT -82.175 -178.075 -81.915 -176.935 ;
        RECT -81.245 -178.075 -80.965 -176.935 ;
        RECT -80.795 -178.075 -80.505 -176.910 ;
        RECT -80.335 -178.075 -80.055 -176.935 ;
        RECT -79.385 -178.075 -79.125 -176.935 ;
        RECT -72.255 -178.075 -71.995 -176.935 ;
        RECT -71.325 -178.075 -71.045 -176.935 ;
        RECT -70.875 -178.075 -70.585 -176.910 ;
        RECT -70.415 -178.075 -70.135 -176.935 ;
        RECT -69.465 -178.075 -69.205 -176.935 ;
        RECT -62.335 -178.075 -62.075 -176.935 ;
        RECT -61.405 -178.075 -61.125 -176.935 ;
        RECT -60.955 -178.075 -60.665 -176.910 ;
        RECT -60.495 -178.075 -60.215 -176.935 ;
        RECT -59.545 -178.075 -59.285 -176.935 ;
        RECT -52.415 -178.075 -52.155 -176.935 ;
        RECT -51.485 -178.075 -51.205 -176.935 ;
        RECT -51.035 -178.075 -50.745 -176.910 ;
        RECT -50.575 -178.075 -50.295 -176.935 ;
        RECT -49.625 -178.075 -49.365 -176.935 ;
        RECT -42.495 -178.075 -42.235 -176.935 ;
        RECT -41.565 -178.075 -41.285 -176.935 ;
        RECT -41.115 -178.075 -40.825 -176.910 ;
        RECT -40.655 -178.075 -40.375 -176.935 ;
        RECT -39.705 -178.075 -39.445 -176.935 ;
        RECT -32.575 -178.075 -32.315 -176.935 ;
        RECT -31.645 -178.075 -31.365 -176.935 ;
        RECT -31.195 -178.075 -30.905 -176.910 ;
        RECT -30.735 -178.075 -30.455 -176.935 ;
        RECT -29.785 -178.075 -29.525 -176.935 ;
        RECT -22.655 -178.075 -22.395 -176.935 ;
        RECT -21.725 -178.075 -21.445 -176.935 ;
        RECT -21.275 -178.075 -20.985 -176.910 ;
        RECT -20.815 -178.075 -20.535 -176.935 ;
        RECT -19.865 -178.075 -19.605 -176.935 ;
        RECT -12.735 -178.075 -12.475 -176.935 ;
        RECT -11.805 -178.075 -11.525 -176.935 ;
        RECT -11.355 -178.075 -11.065 -176.910 ;
        RECT -10.895 -178.075 -10.615 -176.935 ;
        RECT -9.945 -178.075 -9.685 -176.935 ;
        RECT -2.815 -178.075 -2.555 -176.935 ;
        RECT -1.885 -178.075 -1.605 -176.935 ;
        RECT -1.435 -178.075 -1.145 -176.910 ;
        RECT -0.975 -178.075 -0.695 -176.935 ;
        RECT -0.025 -178.075 0.235 -176.935 ;
        RECT 7.105 -178.075 7.365 -176.935 ;
        RECT 8.035 -178.075 8.315 -176.935 ;
        RECT 8.485 -178.075 8.775 -176.910 ;
        RECT 8.945 -178.075 9.225 -176.935 ;
        RECT 9.895 -178.075 10.155 -176.935 ;
        RECT 17.025 -178.075 17.285 -176.935 ;
        RECT 17.955 -178.075 18.235 -176.935 ;
        RECT 18.405 -178.075 18.695 -176.910 ;
        RECT 18.865 -178.075 19.145 -176.935 ;
        RECT 19.815 -178.075 20.075 -176.935 ;
        RECT 26.945 -178.075 27.205 -176.935 ;
        RECT 27.875 -178.075 28.155 -176.935 ;
        RECT 28.325 -178.075 28.615 -176.910 ;
        RECT -280.660 -178.245 -277.440 -178.075 ;
        RECT -270.740 -178.245 -267.520 -178.075 ;
        RECT -260.820 -178.245 -257.600 -178.075 ;
        RECT -250.900 -178.245 -247.680 -178.075 ;
        RECT -240.980 -178.245 -237.760 -178.075 ;
        RECT -231.060 -178.245 -227.840 -178.075 ;
        RECT -221.140 -178.245 -217.920 -178.075 ;
        RECT -211.220 -178.245 -208.000 -178.075 ;
        RECT -201.300 -178.245 -198.080 -178.075 ;
        RECT -191.380 -178.245 -188.160 -178.075 ;
        RECT -181.460 -178.245 -178.240 -178.075 ;
        RECT -171.540 -178.245 -168.320 -178.075 ;
        RECT -161.620 -178.245 -158.400 -178.075 ;
        RECT -151.700 -178.245 -148.480 -178.075 ;
        RECT -141.780 -178.245 -138.560 -178.075 ;
        RECT -131.860 -178.245 -128.640 -178.075 ;
        RECT -121.940 -178.245 -118.720 -178.075 ;
        RECT -112.020 -178.245 -108.800 -178.075 ;
        RECT -102.100 -178.245 -98.880 -178.075 ;
        RECT -92.180 -178.245 -88.960 -178.075 ;
        RECT -82.260 -178.245 -79.040 -178.075 ;
        RECT -72.340 -178.245 -69.120 -178.075 ;
        RECT -62.420 -178.245 -59.200 -178.075 ;
        RECT -52.500 -178.245 -49.280 -178.075 ;
        RECT -42.580 -178.245 -39.360 -178.075 ;
        RECT -32.660 -178.245 -29.440 -178.075 ;
        RECT -22.740 -178.245 -19.520 -178.075 ;
        RECT -12.820 -178.245 -9.600 -178.075 ;
        RECT -2.900 -178.245 0.320 -178.075 ;
        RECT 7.020 -178.245 10.240 -178.075 ;
        RECT 16.940 -178.245 20.160 -178.075 ;
        RECT 26.860 -178.245 28.700 -178.075 ;
        RECT -284.565 -178.660 -284.395 -178.590 ;
        RECT -283.625 -178.660 -283.455 -178.590 ;
        RECT -284.565 -178.830 -283.455 -178.660 ;
        RECT -284.565 -179.115 -284.395 -178.830 ;
        RECT -285.325 -179.445 -284.395 -179.115 ;
        RECT -284.565 -179.970 -284.395 -179.445 ;
        RECT -284.155 -179.995 -283.865 -178.830 ;
        RECT -283.625 -179.115 -283.455 -178.830 ;
        RECT -274.645 -178.660 -274.475 -178.590 ;
        RECT -273.705 -178.660 -273.535 -178.590 ;
        RECT -274.645 -178.830 -273.535 -178.660 ;
        RECT -274.645 -179.115 -274.475 -178.830 ;
        RECT -283.625 -179.445 -282.695 -179.115 ;
        RECT -275.405 -179.445 -274.475 -179.115 ;
        RECT -283.625 -179.970 -283.455 -179.445 ;
        RECT -274.645 -179.970 -274.475 -179.445 ;
        RECT -274.235 -179.995 -273.945 -178.830 ;
        RECT -273.705 -179.115 -273.535 -178.830 ;
        RECT -264.725 -178.660 -264.555 -178.590 ;
        RECT -263.785 -178.660 -263.615 -178.590 ;
        RECT -264.725 -178.830 -263.615 -178.660 ;
        RECT -264.725 -179.115 -264.555 -178.830 ;
        RECT -273.705 -179.445 -272.775 -179.115 ;
        RECT -265.485 -179.445 -264.555 -179.115 ;
        RECT -273.705 -179.970 -273.535 -179.445 ;
        RECT -264.725 -179.970 -264.555 -179.445 ;
        RECT -264.315 -179.995 -264.025 -178.830 ;
        RECT -263.785 -179.115 -263.615 -178.830 ;
        RECT -254.805 -178.660 -254.635 -178.590 ;
        RECT -253.865 -178.660 -253.695 -178.590 ;
        RECT -254.805 -178.830 -253.695 -178.660 ;
        RECT -254.805 -179.115 -254.635 -178.830 ;
        RECT -263.785 -179.445 -262.855 -179.115 ;
        RECT -255.565 -179.445 -254.635 -179.115 ;
        RECT -263.785 -179.970 -263.615 -179.445 ;
        RECT -254.805 -179.970 -254.635 -179.445 ;
        RECT -254.395 -179.995 -254.105 -178.830 ;
        RECT -253.865 -179.115 -253.695 -178.830 ;
        RECT -244.885 -178.660 -244.715 -178.590 ;
        RECT -243.945 -178.660 -243.775 -178.590 ;
        RECT -244.885 -178.830 -243.775 -178.660 ;
        RECT -244.885 -179.115 -244.715 -178.830 ;
        RECT -253.865 -179.445 -252.935 -179.115 ;
        RECT -245.645 -179.445 -244.715 -179.115 ;
        RECT -253.865 -179.970 -253.695 -179.445 ;
        RECT -244.885 -179.970 -244.715 -179.445 ;
        RECT -244.475 -179.995 -244.185 -178.830 ;
        RECT -243.945 -179.115 -243.775 -178.830 ;
        RECT -234.965 -178.660 -234.795 -178.590 ;
        RECT -234.025 -178.660 -233.855 -178.590 ;
        RECT -234.965 -178.830 -233.855 -178.660 ;
        RECT -234.965 -179.115 -234.795 -178.830 ;
        RECT -243.945 -179.445 -243.015 -179.115 ;
        RECT -235.725 -179.445 -234.795 -179.115 ;
        RECT -243.945 -179.970 -243.775 -179.445 ;
        RECT -234.965 -179.970 -234.795 -179.445 ;
        RECT -234.555 -179.995 -234.265 -178.830 ;
        RECT -234.025 -179.115 -233.855 -178.830 ;
        RECT -225.045 -178.660 -224.875 -178.590 ;
        RECT -224.105 -178.660 -223.935 -178.590 ;
        RECT -225.045 -178.830 -223.935 -178.660 ;
        RECT -225.045 -179.115 -224.875 -178.830 ;
        RECT -234.025 -179.445 -233.095 -179.115 ;
        RECT -225.805 -179.445 -224.875 -179.115 ;
        RECT -234.025 -179.970 -233.855 -179.445 ;
        RECT -225.045 -179.970 -224.875 -179.445 ;
        RECT -224.635 -179.995 -224.345 -178.830 ;
        RECT -224.105 -179.115 -223.935 -178.830 ;
        RECT -215.125 -178.660 -214.955 -178.590 ;
        RECT -214.185 -178.660 -214.015 -178.590 ;
        RECT -215.125 -178.830 -214.015 -178.660 ;
        RECT -215.125 -179.115 -214.955 -178.830 ;
        RECT -224.105 -179.445 -223.175 -179.115 ;
        RECT -215.885 -179.445 -214.955 -179.115 ;
        RECT -224.105 -179.970 -223.935 -179.445 ;
        RECT -215.125 -179.970 -214.955 -179.445 ;
        RECT -214.715 -179.995 -214.425 -178.830 ;
        RECT -214.185 -179.115 -214.015 -178.830 ;
        RECT -205.205 -178.660 -205.035 -178.590 ;
        RECT -204.265 -178.660 -204.095 -178.590 ;
        RECT -205.205 -178.830 -204.095 -178.660 ;
        RECT -205.205 -179.115 -205.035 -178.830 ;
        RECT -214.185 -179.445 -213.255 -179.115 ;
        RECT -205.965 -179.445 -205.035 -179.115 ;
        RECT -214.185 -179.970 -214.015 -179.445 ;
        RECT -205.205 -179.970 -205.035 -179.445 ;
        RECT -204.795 -179.995 -204.505 -178.830 ;
        RECT -204.265 -179.115 -204.095 -178.830 ;
        RECT -195.285 -178.660 -195.115 -178.590 ;
        RECT -194.345 -178.660 -194.175 -178.590 ;
        RECT -195.285 -178.830 -194.175 -178.660 ;
        RECT -195.285 -179.115 -195.115 -178.830 ;
        RECT -204.265 -179.445 -203.335 -179.115 ;
        RECT -196.045 -179.445 -195.115 -179.115 ;
        RECT -204.265 -179.970 -204.095 -179.445 ;
        RECT -195.285 -179.970 -195.115 -179.445 ;
        RECT -194.875 -179.995 -194.585 -178.830 ;
        RECT -194.345 -179.115 -194.175 -178.830 ;
        RECT -185.365 -178.660 -185.195 -178.590 ;
        RECT -184.425 -178.660 -184.255 -178.590 ;
        RECT -185.365 -178.830 -184.255 -178.660 ;
        RECT -185.365 -179.115 -185.195 -178.830 ;
        RECT -194.345 -179.445 -193.415 -179.115 ;
        RECT -186.125 -179.445 -185.195 -179.115 ;
        RECT -194.345 -179.970 -194.175 -179.445 ;
        RECT -185.365 -179.970 -185.195 -179.445 ;
        RECT -184.955 -179.995 -184.665 -178.830 ;
        RECT -184.425 -179.115 -184.255 -178.830 ;
        RECT -175.445 -178.660 -175.275 -178.590 ;
        RECT -174.505 -178.660 -174.335 -178.590 ;
        RECT -175.445 -178.830 -174.335 -178.660 ;
        RECT -175.445 -179.115 -175.275 -178.830 ;
        RECT -184.425 -179.445 -183.495 -179.115 ;
        RECT -176.205 -179.445 -175.275 -179.115 ;
        RECT -184.425 -179.970 -184.255 -179.445 ;
        RECT -175.445 -179.970 -175.275 -179.445 ;
        RECT -175.035 -179.995 -174.745 -178.830 ;
        RECT -174.505 -179.115 -174.335 -178.830 ;
        RECT -165.525 -178.660 -165.355 -178.590 ;
        RECT -164.585 -178.660 -164.415 -178.590 ;
        RECT -165.525 -178.830 -164.415 -178.660 ;
        RECT -165.525 -179.115 -165.355 -178.830 ;
        RECT -174.505 -179.445 -173.575 -179.115 ;
        RECT -166.285 -179.445 -165.355 -179.115 ;
        RECT -174.505 -179.970 -174.335 -179.445 ;
        RECT -165.525 -179.970 -165.355 -179.445 ;
        RECT -165.115 -179.995 -164.825 -178.830 ;
        RECT -164.585 -179.115 -164.415 -178.830 ;
        RECT -155.605 -178.660 -155.435 -178.590 ;
        RECT -154.665 -178.660 -154.495 -178.590 ;
        RECT -155.605 -178.830 -154.495 -178.660 ;
        RECT -155.605 -179.115 -155.435 -178.830 ;
        RECT -164.585 -179.445 -163.655 -179.115 ;
        RECT -156.365 -179.445 -155.435 -179.115 ;
        RECT -164.585 -179.970 -164.415 -179.445 ;
        RECT -155.605 -179.970 -155.435 -179.445 ;
        RECT -155.195 -179.995 -154.905 -178.830 ;
        RECT -154.665 -179.115 -154.495 -178.830 ;
        RECT -145.685 -178.660 -145.515 -178.590 ;
        RECT -144.745 -178.660 -144.575 -178.590 ;
        RECT -145.685 -178.830 -144.575 -178.660 ;
        RECT -145.685 -179.115 -145.515 -178.830 ;
        RECT -154.665 -179.445 -153.735 -179.115 ;
        RECT -146.445 -179.445 -145.515 -179.115 ;
        RECT -154.665 -179.970 -154.495 -179.445 ;
        RECT -145.685 -179.970 -145.515 -179.445 ;
        RECT -145.275 -179.995 -144.985 -178.830 ;
        RECT -144.745 -179.115 -144.575 -178.830 ;
        RECT -135.765 -178.660 -135.595 -178.590 ;
        RECT -134.825 -178.660 -134.655 -178.590 ;
        RECT -135.765 -178.830 -134.655 -178.660 ;
        RECT -135.765 -179.115 -135.595 -178.830 ;
        RECT -144.745 -179.445 -143.815 -179.115 ;
        RECT -136.525 -179.445 -135.595 -179.115 ;
        RECT -144.745 -179.970 -144.575 -179.445 ;
        RECT -135.765 -179.970 -135.595 -179.445 ;
        RECT -135.355 -179.995 -135.065 -178.830 ;
        RECT -134.825 -179.115 -134.655 -178.830 ;
        RECT -125.845 -178.660 -125.675 -178.590 ;
        RECT -124.905 -178.660 -124.735 -178.590 ;
        RECT -125.845 -178.830 -124.735 -178.660 ;
        RECT -125.845 -179.115 -125.675 -178.830 ;
        RECT -134.825 -179.445 -133.895 -179.115 ;
        RECT -126.605 -179.445 -125.675 -179.115 ;
        RECT -134.825 -179.970 -134.655 -179.445 ;
        RECT -125.845 -179.970 -125.675 -179.445 ;
        RECT -125.435 -179.995 -125.145 -178.830 ;
        RECT -124.905 -179.115 -124.735 -178.830 ;
        RECT -115.925 -178.660 -115.755 -178.590 ;
        RECT -114.985 -178.660 -114.815 -178.590 ;
        RECT -115.925 -178.830 -114.815 -178.660 ;
        RECT -115.925 -179.115 -115.755 -178.830 ;
        RECT -124.905 -179.445 -123.975 -179.115 ;
        RECT -116.685 -179.445 -115.755 -179.115 ;
        RECT -124.905 -179.970 -124.735 -179.445 ;
        RECT -115.925 -179.970 -115.755 -179.445 ;
        RECT -115.515 -179.995 -115.225 -178.830 ;
        RECT -114.985 -179.115 -114.815 -178.830 ;
        RECT -106.005 -178.660 -105.835 -178.590 ;
        RECT -105.065 -178.660 -104.895 -178.590 ;
        RECT -106.005 -178.830 -104.895 -178.660 ;
        RECT -106.005 -179.115 -105.835 -178.830 ;
        RECT -114.985 -179.445 -114.055 -179.115 ;
        RECT -106.765 -179.445 -105.835 -179.115 ;
        RECT -114.985 -179.970 -114.815 -179.445 ;
        RECT -106.005 -179.970 -105.835 -179.445 ;
        RECT -105.595 -179.995 -105.305 -178.830 ;
        RECT -105.065 -179.115 -104.895 -178.830 ;
        RECT -96.085 -178.660 -95.915 -178.590 ;
        RECT -95.145 -178.660 -94.975 -178.590 ;
        RECT -96.085 -178.830 -94.975 -178.660 ;
        RECT -96.085 -179.115 -95.915 -178.830 ;
        RECT -105.065 -179.445 -104.135 -179.115 ;
        RECT -96.845 -179.445 -95.915 -179.115 ;
        RECT -105.065 -179.970 -104.895 -179.445 ;
        RECT -96.085 -179.970 -95.915 -179.445 ;
        RECT -95.675 -179.995 -95.385 -178.830 ;
        RECT -95.145 -179.115 -94.975 -178.830 ;
        RECT -86.165 -178.660 -85.995 -178.590 ;
        RECT -85.225 -178.660 -85.055 -178.590 ;
        RECT -86.165 -178.830 -85.055 -178.660 ;
        RECT -86.165 -179.115 -85.995 -178.830 ;
        RECT -95.145 -179.445 -94.215 -179.115 ;
        RECT -86.925 -179.445 -85.995 -179.115 ;
        RECT -95.145 -179.970 -94.975 -179.445 ;
        RECT -86.165 -179.970 -85.995 -179.445 ;
        RECT -85.755 -179.995 -85.465 -178.830 ;
        RECT -85.225 -179.115 -85.055 -178.830 ;
        RECT -76.245 -178.660 -76.075 -178.590 ;
        RECT -75.305 -178.660 -75.135 -178.590 ;
        RECT -76.245 -178.830 -75.135 -178.660 ;
        RECT -76.245 -179.115 -76.075 -178.830 ;
        RECT -85.225 -179.445 -84.295 -179.115 ;
        RECT -77.005 -179.445 -76.075 -179.115 ;
        RECT -85.225 -179.970 -85.055 -179.445 ;
        RECT -76.245 -179.970 -76.075 -179.445 ;
        RECT -75.835 -179.995 -75.545 -178.830 ;
        RECT -75.305 -179.115 -75.135 -178.830 ;
        RECT -66.325 -178.660 -66.155 -178.590 ;
        RECT -65.385 -178.660 -65.215 -178.590 ;
        RECT -66.325 -178.830 -65.215 -178.660 ;
        RECT -66.325 -179.115 -66.155 -178.830 ;
        RECT -75.305 -179.445 -74.375 -179.115 ;
        RECT -67.085 -179.445 -66.155 -179.115 ;
        RECT -75.305 -179.970 -75.135 -179.445 ;
        RECT -66.325 -179.970 -66.155 -179.445 ;
        RECT -65.915 -179.995 -65.625 -178.830 ;
        RECT -65.385 -179.115 -65.215 -178.830 ;
        RECT -56.405 -178.660 -56.235 -178.590 ;
        RECT -55.465 -178.660 -55.295 -178.590 ;
        RECT -56.405 -178.830 -55.295 -178.660 ;
        RECT -56.405 -179.115 -56.235 -178.830 ;
        RECT -65.385 -179.445 -64.455 -179.115 ;
        RECT -57.165 -179.445 -56.235 -179.115 ;
        RECT -65.385 -179.970 -65.215 -179.445 ;
        RECT -56.405 -179.970 -56.235 -179.445 ;
        RECT -55.995 -179.995 -55.705 -178.830 ;
        RECT -55.465 -179.115 -55.295 -178.830 ;
        RECT -46.485 -178.660 -46.315 -178.590 ;
        RECT -45.545 -178.660 -45.375 -178.590 ;
        RECT -46.485 -178.830 -45.375 -178.660 ;
        RECT -46.485 -179.115 -46.315 -178.830 ;
        RECT -55.465 -179.445 -54.535 -179.115 ;
        RECT -47.245 -179.445 -46.315 -179.115 ;
        RECT -55.465 -179.970 -55.295 -179.445 ;
        RECT -46.485 -179.970 -46.315 -179.445 ;
        RECT -46.075 -179.995 -45.785 -178.830 ;
        RECT -45.545 -179.115 -45.375 -178.830 ;
        RECT -36.565 -178.660 -36.395 -178.590 ;
        RECT -35.625 -178.660 -35.455 -178.590 ;
        RECT -36.565 -178.830 -35.455 -178.660 ;
        RECT -36.565 -179.115 -36.395 -178.830 ;
        RECT -45.545 -179.445 -44.615 -179.115 ;
        RECT -37.325 -179.445 -36.395 -179.115 ;
        RECT -45.545 -179.970 -45.375 -179.445 ;
        RECT -36.565 -179.970 -36.395 -179.445 ;
        RECT -36.155 -179.995 -35.865 -178.830 ;
        RECT -35.625 -179.115 -35.455 -178.830 ;
        RECT -26.645 -178.660 -26.475 -178.590 ;
        RECT -25.705 -178.660 -25.535 -178.590 ;
        RECT -26.645 -178.830 -25.535 -178.660 ;
        RECT -26.645 -179.115 -26.475 -178.830 ;
        RECT -35.625 -179.445 -34.695 -179.115 ;
        RECT -27.405 -179.445 -26.475 -179.115 ;
        RECT -35.625 -179.970 -35.455 -179.445 ;
        RECT -26.645 -179.970 -26.475 -179.445 ;
        RECT -26.235 -179.995 -25.945 -178.830 ;
        RECT -25.705 -179.115 -25.535 -178.830 ;
        RECT -16.725 -178.660 -16.555 -178.590 ;
        RECT -15.785 -178.660 -15.615 -178.590 ;
        RECT -16.725 -178.830 -15.615 -178.660 ;
        RECT -16.725 -179.115 -16.555 -178.830 ;
        RECT -25.705 -179.445 -24.775 -179.115 ;
        RECT -17.485 -179.445 -16.555 -179.115 ;
        RECT -25.705 -179.970 -25.535 -179.445 ;
        RECT -16.725 -179.970 -16.555 -179.445 ;
        RECT -16.315 -179.995 -16.025 -178.830 ;
        RECT -15.785 -179.115 -15.615 -178.830 ;
        RECT -6.805 -178.660 -6.635 -178.590 ;
        RECT -5.865 -178.660 -5.695 -178.590 ;
        RECT -6.805 -178.830 -5.695 -178.660 ;
        RECT -6.805 -179.115 -6.635 -178.830 ;
        RECT -15.785 -179.445 -14.855 -179.115 ;
        RECT -7.565 -179.445 -6.635 -179.115 ;
        RECT -15.785 -179.970 -15.615 -179.445 ;
        RECT -6.805 -179.970 -6.635 -179.445 ;
        RECT -6.395 -179.995 -6.105 -178.830 ;
        RECT -5.865 -179.115 -5.695 -178.830 ;
        RECT 3.115 -178.660 3.285 -178.590 ;
        RECT 4.055 -178.660 4.225 -178.590 ;
        RECT 3.115 -178.830 4.225 -178.660 ;
        RECT 3.115 -179.115 3.285 -178.830 ;
        RECT -5.865 -179.445 -4.935 -179.115 ;
        RECT 2.355 -179.445 3.285 -179.115 ;
        RECT -5.865 -179.970 -5.695 -179.445 ;
        RECT 3.115 -179.970 3.285 -179.445 ;
        RECT 3.525 -179.995 3.815 -178.830 ;
        RECT 4.055 -179.115 4.225 -178.830 ;
        RECT 13.035 -178.660 13.205 -178.590 ;
        RECT 13.975 -178.660 14.145 -178.590 ;
        RECT 13.035 -178.830 14.145 -178.660 ;
        RECT 13.035 -179.115 13.205 -178.830 ;
        RECT 4.055 -179.445 4.985 -179.115 ;
        RECT 12.275 -179.445 13.205 -179.115 ;
        RECT 4.055 -179.970 4.225 -179.445 ;
        RECT 13.035 -179.970 13.205 -179.445 ;
        RECT 13.445 -179.995 13.735 -178.830 ;
        RECT 13.975 -179.115 14.145 -178.830 ;
        RECT 22.955 -178.660 23.125 -178.590 ;
        RECT 23.895 -178.660 24.065 -178.590 ;
        RECT 22.955 -178.830 24.065 -178.660 ;
        RECT 22.955 -179.115 23.125 -178.830 ;
        RECT 13.975 -179.445 14.905 -179.115 ;
        RECT 22.195 -179.445 23.125 -179.115 ;
        RECT 13.975 -179.970 14.145 -179.445 ;
        RECT 22.955 -179.970 23.125 -179.445 ;
        RECT 23.365 -179.995 23.655 -178.830 ;
        RECT 23.895 -179.115 24.065 -178.830 ;
        RECT 23.895 -179.445 24.825 -179.115 ;
        RECT 23.895 -179.970 24.065 -179.445 ;
      LAYER mcon ;
        RECT -281.865 94.825 -281.695 94.995 ;
        RECT -281.395 94.820 -281.225 94.990 ;
        RECT -280.925 94.825 -280.755 94.995 ;
        RECT -281.865 94.365 -281.695 94.535 ;
        RECT -281.865 93.905 -281.695 94.075 ;
        RECT -271.945 94.825 -271.775 94.995 ;
        RECT -271.475 94.820 -271.305 94.990 ;
        RECT -271.005 94.825 -270.835 94.995 ;
        RECT -280.925 94.365 -280.755 94.535 ;
        RECT -271.945 94.365 -271.775 94.535 ;
        RECT -280.925 93.905 -280.755 94.075 ;
        RECT -271.945 93.905 -271.775 94.075 ;
        RECT -262.025 94.825 -261.855 94.995 ;
        RECT -261.555 94.820 -261.385 94.990 ;
        RECT -261.085 94.825 -260.915 94.995 ;
        RECT -271.005 94.365 -270.835 94.535 ;
        RECT -262.025 94.365 -261.855 94.535 ;
        RECT -271.005 93.905 -270.835 94.075 ;
        RECT -262.025 93.905 -261.855 94.075 ;
        RECT -252.105 94.825 -251.935 94.995 ;
        RECT -251.635 94.820 -251.465 94.990 ;
        RECT -251.165 94.825 -250.995 94.995 ;
        RECT -261.085 94.365 -260.915 94.535 ;
        RECT -252.105 94.365 -251.935 94.535 ;
        RECT -261.085 93.905 -260.915 94.075 ;
        RECT -252.105 93.905 -251.935 94.075 ;
        RECT -242.185 94.825 -242.015 94.995 ;
        RECT -241.715 94.820 -241.545 94.990 ;
        RECT -241.245 94.825 -241.075 94.995 ;
        RECT -251.165 94.365 -250.995 94.535 ;
        RECT -242.185 94.365 -242.015 94.535 ;
        RECT -251.165 93.905 -250.995 94.075 ;
        RECT -242.185 93.905 -242.015 94.075 ;
        RECT -232.265 94.825 -232.095 94.995 ;
        RECT -231.795 94.820 -231.625 94.990 ;
        RECT -231.325 94.825 -231.155 94.995 ;
        RECT -241.245 94.365 -241.075 94.535 ;
        RECT -232.265 94.365 -232.095 94.535 ;
        RECT -241.245 93.905 -241.075 94.075 ;
        RECT -232.265 93.905 -232.095 94.075 ;
        RECT -222.345 94.825 -222.175 94.995 ;
        RECT -221.875 94.820 -221.705 94.990 ;
        RECT -221.405 94.825 -221.235 94.995 ;
        RECT -231.325 94.365 -231.155 94.535 ;
        RECT -222.345 94.365 -222.175 94.535 ;
        RECT -231.325 93.905 -231.155 94.075 ;
        RECT -222.345 93.905 -222.175 94.075 ;
        RECT -212.425 94.825 -212.255 94.995 ;
        RECT -211.955 94.820 -211.785 94.990 ;
        RECT -211.485 94.825 -211.315 94.995 ;
        RECT -221.405 94.365 -221.235 94.535 ;
        RECT -212.425 94.365 -212.255 94.535 ;
        RECT -221.405 93.905 -221.235 94.075 ;
        RECT -212.425 93.905 -212.255 94.075 ;
        RECT -202.505 94.825 -202.335 94.995 ;
        RECT -202.035 94.820 -201.865 94.990 ;
        RECT -201.565 94.825 -201.395 94.995 ;
        RECT -211.485 94.365 -211.315 94.535 ;
        RECT -202.505 94.365 -202.335 94.535 ;
        RECT -211.485 93.905 -211.315 94.075 ;
        RECT -202.505 93.905 -202.335 94.075 ;
        RECT -192.585 94.825 -192.415 94.995 ;
        RECT -192.115 94.820 -191.945 94.990 ;
        RECT -191.645 94.825 -191.475 94.995 ;
        RECT -201.565 94.365 -201.395 94.535 ;
        RECT -192.585 94.365 -192.415 94.535 ;
        RECT -201.565 93.905 -201.395 94.075 ;
        RECT -192.585 93.905 -192.415 94.075 ;
        RECT -182.665 94.825 -182.495 94.995 ;
        RECT -182.195 94.820 -182.025 94.990 ;
        RECT -181.725 94.825 -181.555 94.995 ;
        RECT -191.645 94.365 -191.475 94.535 ;
        RECT -182.665 94.365 -182.495 94.535 ;
        RECT -191.645 93.905 -191.475 94.075 ;
        RECT -182.665 93.905 -182.495 94.075 ;
        RECT -172.745 94.825 -172.575 94.995 ;
        RECT -172.275 94.820 -172.105 94.990 ;
        RECT -171.805 94.825 -171.635 94.995 ;
        RECT -181.725 94.365 -181.555 94.535 ;
        RECT -172.745 94.365 -172.575 94.535 ;
        RECT -181.725 93.905 -181.555 94.075 ;
        RECT -172.745 93.905 -172.575 94.075 ;
        RECT -162.825 94.825 -162.655 94.995 ;
        RECT -162.355 94.820 -162.185 94.990 ;
        RECT -161.885 94.825 -161.715 94.995 ;
        RECT -171.805 94.365 -171.635 94.535 ;
        RECT -162.825 94.365 -162.655 94.535 ;
        RECT -171.805 93.905 -171.635 94.075 ;
        RECT -162.825 93.905 -162.655 94.075 ;
        RECT -152.905 94.825 -152.735 94.995 ;
        RECT -152.435 94.820 -152.265 94.990 ;
        RECT -151.965 94.825 -151.795 94.995 ;
        RECT -161.885 94.365 -161.715 94.535 ;
        RECT -152.905 94.365 -152.735 94.535 ;
        RECT -161.885 93.905 -161.715 94.075 ;
        RECT -152.905 93.905 -152.735 94.075 ;
        RECT -142.985 94.825 -142.815 94.995 ;
        RECT -142.515 94.820 -142.345 94.990 ;
        RECT -142.045 94.825 -141.875 94.995 ;
        RECT -151.965 94.365 -151.795 94.535 ;
        RECT -142.985 94.365 -142.815 94.535 ;
        RECT -151.965 93.905 -151.795 94.075 ;
        RECT -142.985 93.905 -142.815 94.075 ;
        RECT -133.065 94.825 -132.895 94.995 ;
        RECT -132.595 94.820 -132.425 94.990 ;
        RECT -132.125 94.825 -131.955 94.995 ;
        RECT -142.045 94.365 -141.875 94.535 ;
        RECT -133.065 94.365 -132.895 94.535 ;
        RECT -142.045 93.905 -141.875 94.075 ;
        RECT -133.065 93.905 -132.895 94.075 ;
        RECT -123.145 94.825 -122.975 94.995 ;
        RECT -122.675 94.820 -122.505 94.990 ;
        RECT -122.205 94.825 -122.035 94.995 ;
        RECT -132.125 94.365 -131.955 94.535 ;
        RECT -123.145 94.365 -122.975 94.535 ;
        RECT -132.125 93.905 -131.955 94.075 ;
        RECT -123.145 93.905 -122.975 94.075 ;
        RECT -113.225 94.825 -113.055 94.995 ;
        RECT -112.755 94.820 -112.585 94.990 ;
        RECT -112.285 94.825 -112.115 94.995 ;
        RECT -122.205 94.365 -122.035 94.535 ;
        RECT -113.225 94.365 -113.055 94.535 ;
        RECT -122.205 93.905 -122.035 94.075 ;
        RECT -113.225 93.905 -113.055 94.075 ;
        RECT -103.305 94.825 -103.135 94.995 ;
        RECT -102.835 94.820 -102.665 94.990 ;
        RECT -102.365 94.825 -102.195 94.995 ;
        RECT -112.285 94.365 -112.115 94.535 ;
        RECT -103.305 94.365 -103.135 94.535 ;
        RECT -112.285 93.905 -112.115 94.075 ;
        RECT -103.305 93.905 -103.135 94.075 ;
        RECT -93.385 94.825 -93.215 94.995 ;
        RECT -92.915 94.820 -92.745 94.990 ;
        RECT -92.445 94.825 -92.275 94.995 ;
        RECT -102.365 94.365 -102.195 94.535 ;
        RECT -93.385 94.365 -93.215 94.535 ;
        RECT -102.365 93.905 -102.195 94.075 ;
        RECT -93.385 93.905 -93.215 94.075 ;
        RECT -83.465 94.825 -83.295 94.995 ;
        RECT -82.995 94.820 -82.825 94.990 ;
        RECT -82.525 94.825 -82.355 94.995 ;
        RECT -92.445 94.365 -92.275 94.535 ;
        RECT -83.465 94.365 -83.295 94.535 ;
        RECT -92.445 93.905 -92.275 94.075 ;
        RECT -83.465 93.905 -83.295 94.075 ;
        RECT -73.545 94.825 -73.375 94.995 ;
        RECT -73.075 94.820 -72.905 94.990 ;
        RECT -72.605 94.825 -72.435 94.995 ;
        RECT -82.525 94.365 -82.355 94.535 ;
        RECT -73.545 94.365 -73.375 94.535 ;
        RECT -82.525 93.905 -82.355 94.075 ;
        RECT -73.545 93.905 -73.375 94.075 ;
        RECT -63.625 94.825 -63.455 94.995 ;
        RECT -63.155 94.820 -62.985 94.990 ;
        RECT -62.685 94.825 -62.515 94.995 ;
        RECT -72.605 94.365 -72.435 94.535 ;
        RECT -63.625 94.365 -63.455 94.535 ;
        RECT -72.605 93.905 -72.435 94.075 ;
        RECT -63.625 93.905 -63.455 94.075 ;
        RECT -53.705 94.825 -53.535 94.995 ;
        RECT -53.235 94.820 -53.065 94.990 ;
        RECT -52.765 94.825 -52.595 94.995 ;
        RECT -62.685 94.365 -62.515 94.535 ;
        RECT -53.705 94.365 -53.535 94.535 ;
        RECT -62.685 93.905 -62.515 94.075 ;
        RECT -53.705 93.905 -53.535 94.075 ;
        RECT -43.785 94.825 -43.615 94.995 ;
        RECT -43.315 94.820 -43.145 94.990 ;
        RECT -42.845 94.825 -42.675 94.995 ;
        RECT -52.765 94.365 -52.595 94.535 ;
        RECT -43.785 94.365 -43.615 94.535 ;
        RECT -52.765 93.905 -52.595 94.075 ;
        RECT -43.785 93.905 -43.615 94.075 ;
        RECT -33.865 94.825 -33.695 94.995 ;
        RECT -33.395 94.820 -33.225 94.990 ;
        RECT -32.925 94.825 -32.755 94.995 ;
        RECT -42.845 94.365 -42.675 94.535 ;
        RECT -33.865 94.365 -33.695 94.535 ;
        RECT -42.845 93.905 -42.675 94.075 ;
        RECT -33.865 93.905 -33.695 94.075 ;
        RECT -23.945 94.825 -23.775 94.995 ;
        RECT -23.475 94.820 -23.305 94.990 ;
        RECT -23.005 94.825 -22.835 94.995 ;
        RECT -32.925 94.365 -32.755 94.535 ;
        RECT -23.945 94.365 -23.775 94.535 ;
        RECT -32.925 93.905 -32.755 94.075 ;
        RECT -23.945 93.905 -23.775 94.075 ;
        RECT -14.025 94.825 -13.855 94.995 ;
        RECT -13.555 94.820 -13.385 94.990 ;
        RECT -13.085 94.825 -12.915 94.995 ;
        RECT -23.005 94.365 -22.835 94.535 ;
        RECT -14.025 94.365 -13.855 94.535 ;
        RECT -23.005 93.905 -22.835 94.075 ;
        RECT -14.025 93.905 -13.855 94.075 ;
        RECT -4.105 94.825 -3.935 94.995 ;
        RECT -3.635 94.820 -3.465 94.990 ;
        RECT -3.165 94.825 -2.995 94.995 ;
        RECT -13.085 94.365 -12.915 94.535 ;
        RECT -4.105 94.365 -3.935 94.535 ;
        RECT -13.085 93.905 -12.915 94.075 ;
        RECT -4.105 93.905 -3.935 94.075 ;
        RECT 5.815 94.825 5.985 94.995 ;
        RECT 6.285 94.820 6.455 94.990 ;
        RECT 6.755 94.825 6.925 94.995 ;
        RECT -3.165 94.365 -2.995 94.535 ;
        RECT 5.815 94.365 5.985 94.535 ;
        RECT -3.165 93.905 -2.995 94.075 ;
        RECT 5.815 93.905 5.985 94.075 ;
        RECT 15.735 94.825 15.905 94.995 ;
        RECT 16.205 94.820 16.375 94.990 ;
        RECT 16.675 94.825 16.845 94.995 ;
        RECT 6.755 94.365 6.925 94.535 ;
        RECT 15.735 94.365 15.905 94.535 ;
        RECT 6.755 93.905 6.925 94.075 ;
        RECT 15.735 93.905 15.905 94.075 ;
        RECT 25.655 94.825 25.825 94.995 ;
        RECT 26.125 94.820 26.295 94.990 ;
        RECT 16.675 94.365 16.845 94.535 ;
        RECT 25.655 94.365 25.825 94.535 ;
        RECT 16.675 93.905 16.845 94.075 ;
        RECT 25.655 93.905 25.825 94.075 ;
        RECT -287.735 93.245 -287.565 93.415 ;
        RECT -287.275 93.245 -287.105 93.415 ;
        RECT -286.815 93.245 -286.645 93.415 ;
        RECT -286.355 93.245 -286.185 93.415 ;
        RECT -285.895 93.245 -285.725 93.415 ;
        RECT -285.435 93.245 -285.265 93.415 ;
        RECT -284.975 93.245 -284.805 93.415 ;
        RECT -277.815 93.245 -277.645 93.415 ;
        RECT -277.355 93.245 -277.185 93.415 ;
        RECT -276.895 93.245 -276.725 93.415 ;
        RECT -276.435 93.245 -276.265 93.415 ;
        RECT -275.975 93.245 -275.805 93.415 ;
        RECT -275.515 93.245 -275.345 93.415 ;
        RECT -275.055 93.245 -274.885 93.415 ;
        RECT -267.895 93.245 -267.725 93.415 ;
        RECT -267.435 93.245 -267.265 93.415 ;
        RECT -266.975 93.245 -266.805 93.415 ;
        RECT -266.515 93.245 -266.345 93.415 ;
        RECT -266.055 93.245 -265.885 93.415 ;
        RECT -265.595 93.245 -265.425 93.415 ;
        RECT -265.135 93.245 -264.965 93.415 ;
        RECT -257.975 93.245 -257.805 93.415 ;
        RECT -257.515 93.245 -257.345 93.415 ;
        RECT -257.055 93.245 -256.885 93.415 ;
        RECT -256.595 93.245 -256.425 93.415 ;
        RECT -256.135 93.245 -255.965 93.415 ;
        RECT -255.675 93.245 -255.505 93.415 ;
        RECT -255.215 93.245 -255.045 93.415 ;
        RECT -248.055 93.245 -247.885 93.415 ;
        RECT -247.595 93.245 -247.425 93.415 ;
        RECT -247.135 93.245 -246.965 93.415 ;
        RECT -246.675 93.245 -246.505 93.415 ;
        RECT -246.215 93.245 -246.045 93.415 ;
        RECT -245.755 93.245 -245.585 93.415 ;
        RECT -245.295 93.245 -245.125 93.415 ;
        RECT -238.135 93.245 -237.965 93.415 ;
        RECT -237.675 93.245 -237.505 93.415 ;
        RECT -237.215 93.245 -237.045 93.415 ;
        RECT -236.755 93.245 -236.585 93.415 ;
        RECT -236.295 93.245 -236.125 93.415 ;
        RECT -235.835 93.245 -235.665 93.415 ;
        RECT -235.375 93.245 -235.205 93.415 ;
        RECT -228.215 93.245 -228.045 93.415 ;
        RECT -227.755 93.245 -227.585 93.415 ;
        RECT -227.295 93.245 -227.125 93.415 ;
        RECT -226.835 93.245 -226.665 93.415 ;
        RECT -226.375 93.245 -226.205 93.415 ;
        RECT -225.915 93.245 -225.745 93.415 ;
        RECT -225.455 93.245 -225.285 93.415 ;
        RECT -218.295 93.245 -218.125 93.415 ;
        RECT -217.835 93.245 -217.665 93.415 ;
        RECT -217.375 93.245 -217.205 93.415 ;
        RECT -216.915 93.245 -216.745 93.415 ;
        RECT -216.455 93.245 -216.285 93.415 ;
        RECT -215.995 93.245 -215.825 93.415 ;
        RECT -215.535 93.245 -215.365 93.415 ;
        RECT -208.375 93.245 -208.205 93.415 ;
        RECT -207.915 93.245 -207.745 93.415 ;
        RECT -207.455 93.245 -207.285 93.415 ;
        RECT -206.995 93.245 -206.825 93.415 ;
        RECT -206.535 93.245 -206.365 93.415 ;
        RECT -206.075 93.245 -205.905 93.415 ;
        RECT -205.615 93.245 -205.445 93.415 ;
        RECT -198.455 93.245 -198.285 93.415 ;
        RECT -197.995 93.245 -197.825 93.415 ;
        RECT -197.535 93.245 -197.365 93.415 ;
        RECT -197.075 93.245 -196.905 93.415 ;
        RECT -196.615 93.245 -196.445 93.415 ;
        RECT -196.155 93.245 -195.985 93.415 ;
        RECT -195.695 93.245 -195.525 93.415 ;
        RECT -188.535 93.245 -188.365 93.415 ;
        RECT -188.075 93.245 -187.905 93.415 ;
        RECT -187.615 93.245 -187.445 93.415 ;
        RECT -187.155 93.245 -186.985 93.415 ;
        RECT -186.695 93.245 -186.525 93.415 ;
        RECT -186.235 93.245 -186.065 93.415 ;
        RECT -185.775 93.245 -185.605 93.415 ;
        RECT -178.615 93.245 -178.445 93.415 ;
        RECT -178.155 93.245 -177.985 93.415 ;
        RECT -177.695 93.245 -177.525 93.415 ;
        RECT -177.235 93.245 -177.065 93.415 ;
        RECT -176.775 93.245 -176.605 93.415 ;
        RECT -176.315 93.245 -176.145 93.415 ;
        RECT -175.855 93.245 -175.685 93.415 ;
        RECT -168.695 93.245 -168.525 93.415 ;
        RECT -168.235 93.245 -168.065 93.415 ;
        RECT -167.775 93.245 -167.605 93.415 ;
        RECT -167.315 93.245 -167.145 93.415 ;
        RECT -166.855 93.245 -166.685 93.415 ;
        RECT -166.395 93.245 -166.225 93.415 ;
        RECT -165.935 93.245 -165.765 93.415 ;
        RECT -158.775 93.245 -158.605 93.415 ;
        RECT -158.315 93.245 -158.145 93.415 ;
        RECT -157.855 93.245 -157.685 93.415 ;
        RECT -157.395 93.245 -157.225 93.415 ;
        RECT -156.935 93.245 -156.765 93.415 ;
        RECT -156.475 93.245 -156.305 93.415 ;
        RECT -156.015 93.245 -155.845 93.415 ;
        RECT -148.855 93.245 -148.685 93.415 ;
        RECT -148.395 93.245 -148.225 93.415 ;
        RECT -147.935 93.245 -147.765 93.415 ;
        RECT -147.475 93.245 -147.305 93.415 ;
        RECT -147.015 93.245 -146.845 93.415 ;
        RECT -146.555 93.245 -146.385 93.415 ;
        RECT -146.095 93.245 -145.925 93.415 ;
        RECT -138.935 93.245 -138.765 93.415 ;
        RECT -138.475 93.245 -138.305 93.415 ;
        RECT -138.015 93.245 -137.845 93.415 ;
        RECT -137.555 93.245 -137.385 93.415 ;
        RECT -137.095 93.245 -136.925 93.415 ;
        RECT -136.635 93.245 -136.465 93.415 ;
        RECT -136.175 93.245 -136.005 93.415 ;
        RECT -129.015 93.245 -128.845 93.415 ;
        RECT -128.555 93.245 -128.385 93.415 ;
        RECT -128.095 93.245 -127.925 93.415 ;
        RECT -127.635 93.245 -127.465 93.415 ;
        RECT -127.175 93.245 -127.005 93.415 ;
        RECT -126.715 93.245 -126.545 93.415 ;
        RECT -126.255 93.245 -126.085 93.415 ;
        RECT -119.095 93.245 -118.925 93.415 ;
        RECT -118.635 93.245 -118.465 93.415 ;
        RECT -118.175 93.245 -118.005 93.415 ;
        RECT -117.715 93.245 -117.545 93.415 ;
        RECT -117.255 93.245 -117.085 93.415 ;
        RECT -116.795 93.245 -116.625 93.415 ;
        RECT -116.335 93.245 -116.165 93.415 ;
        RECT -109.175 93.245 -109.005 93.415 ;
        RECT -108.715 93.245 -108.545 93.415 ;
        RECT -108.255 93.245 -108.085 93.415 ;
        RECT -107.795 93.245 -107.625 93.415 ;
        RECT -107.335 93.245 -107.165 93.415 ;
        RECT -106.875 93.245 -106.705 93.415 ;
        RECT -106.415 93.245 -106.245 93.415 ;
        RECT -99.255 93.245 -99.085 93.415 ;
        RECT -98.795 93.245 -98.625 93.415 ;
        RECT -98.335 93.245 -98.165 93.415 ;
        RECT -97.875 93.245 -97.705 93.415 ;
        RECT -97.415 93.245 -97.245 93.415 ;
        RECT -96.955 93.245 -96.785 93.415 ;
        RECT -96.495 93.245 -96.325 93.415 ;
        RECT -89.335 93.245 -89.165 93.415 ;
        RECT -88.875 93.245 -88.705 93.415 ;
        RECT -88.415 93.245 -88.245 93.415 ;
        RECT -87.955 93.245 -87.785 93.415 ;
        RECT -87.495 93.245 -87.325 93.415 ;
        RECT -87.035 93.245 -86.865 93.415 ;
        RECT -86.575 93.245 -86.405 93.415 ;
        RECT -79.415 93.245 -79.245 93.415 ;
        RECT -78.955 93.245 -78.785 93.415 ;
        RECT -78.495 93.245 -78.325 93.415 ;
        RECT -78.035 93.245 -77.865 93.415 ;
        RECT -77.575 93.245 -77.405 93.415 ;
        RECT -77.115 93.245 -76.945 93.415 ;
        RECT -76.655 93.245 -76.485 93.415 ;
        RECT -69.495 93.245 -69.325 93.415 ;
        RECT -69.035 93.245 -68.865 93.415 ;
        RECT -68.575 93.245 -68.405 93.415 ;
        RECT -68.115 93.245 -67.945 93.415 ;
        RECT -67.655 93.245 -67.485 93.415 ;
        RECT -67.195 93.245 -67.025 93.415 ;
        RECT -66.735 93.245 -66.565 93.415 ;
        RECT -59.575 93.245 -59.405 93.415 ;
        RECT -59.115 93.245 -58.945 93.415 ;
        RECT -58.655 93.245 -58.485 93.415 ;
        RECT -58.195 93.245 -58.025 93.415 ;
        RECT -57.735 93.245 -57.565 93.415 ;
        RECT -57.275 93.245 -57.105 93.415 ;
        RECT -56.815 93.245 -56.645 93.415 ;
        RECT -49.655 93.245 -49.485 93.415 ;
        RECT -49.195 93.245 -49.025 93.415 ;
        RECT -48.735 93.245 -48.565 93.415 ;
        RECT -48.275 93.245 -48.105 93.415 ;
        RECT -47.815 93.245 -47.645 93.415 ;
        RECT -47.355 93.245 -47.185 93.415 ;
        RECT -46.895 93.245 -46.725 93.415 ;
        RECT -39.735 93.245 -39.565 93.415 ;
        RECT -39.275 93.245 -39.105 93.415 ;
        RECT -38.815 93.245 -38.645 93.415 ;
        RECT -38.355 93.245 -38.185 93.415 ;
        RECT -37.895 93.245 -37.725 93.415 ;
        RECT -37.435 93.245 -37.265 93.415 ;
        RECT -36.975 93.245 -36.805 93.415 ;
        RECT -29.815 93.245 -29.645 93.415 ;
        RECT -29.355 93.245 -29.185 93.415 ;
        RECT -28.895 93.245 -28.725 93.415 ;
        RECT -28.435 93.245 -28.265 93.415 ;
        RECT -27.975 93.245 -27.805 93.415 ;
        RECT -27.515 93.245 -27.345 93.415 ;
        RECT -27.055 93.245 -26.885 93.415 ;
        RECT -19.895 93.245 -19.725 93.415 ;
        RECT -19.435 93.245 -19.265 93.415 ;
        RECT -18.975 93.245 -18.805 93.415 ;
        RECT -18.515 93.245 -18.345 93.415 ;
        RECT -18.055 93.245 -17.885 93.415 ;
        RECT -17.595 93.245 -17.425 93.415 ;
        RECT -17.135 93.245 -16.965 93.415 ;
        RECT -9.975 93.245 -9.805 93.415 ;
        RECT -9.515 93.245 -9.345 93.415 ;
        RECT -9.055 93.245 -8.885 93.415 ;
        RECT -8.595 93.245 -8.425 93.415 ;
        RECT -8.135 93.245 -7.965 93.415 ;
        RECT -7.675 93.245 -7.505 93.415 ;
        RECT -7.215 93.245 -7.045 93.415 ;
        RECT -0.055 93.245 0.115 93.415 ;
        RECT 0.405 93.245 0.575 93.415 ;
        RECT 0.865 93.245 1.035 93.415 ;
        RECT 1.325 93.245 1.495 93.415 ;
        RECT 1.785 93.245 1.955 93.415 ;
        RECT 2.245 93.245 2.415 93.415 ;
        RECT 2.705 93.245 2.875 93.415 ;
        RECT 9.865 93.245 10.035 93.415 ;
        RECT 10.325 93.245 10.495 93.415 ;
        RECT 10.785 93.245 10.955 93.415 ;
        RECT 11.245 93.245 11.415 93.415 ;
        RECT 11.705 93.245 11.875 93.415 ;
        RECT 12.165 93.245 12.335 93.415 ;
        RECT 12.625 93.245 12.795 93.415 ;
        RECT 19.785 93.245 19.955 93.415 ;
        RECT 20.245 93.245 20.415 93.415 ;
        RECT 20.705 93.245 20.875 93.415 ;
        RECT 21.165 93.245 21.335 93.415 ;
        RECT 21.625 93.245 21.795 93.415 ;
        RECT 22.085 93.245 22.255 93.415 ;
        RECT 22.545 93.245 22.715 93.415 ;
        RECT -282.775 90.525 -282.605 90.695 ;
        RECT -282.315 90.525 -282.145 90.695 ;
        RECT -281.855 90.525 -281.685 90.695 ;
        RECT -281.395 90.525 -281.225 90.695 ;
        RECT -280.935 90.525 -280.765 90.695 ;
        RECT -280.475 90.525 -280.305 90.695 ;
        RECT -280.015 90.525 -279.845 90.695 ;
        RECT -272.855 90.525 -272.685 90.695 ;
        RECT -272.395 90.525 -272.225 90.695 ;
        RECT -271.935 90.525 -271.765 90.695 ;
        RECT -271.475 90.525 -271.305 90.695 ;
        RECT -271.015 90.525 -270.845 90.695 ;
        RECT -270.555 90.525 -270.385 90.695 ;
        RECT -270.095 90.525 -269.925 90.695 ;
        RECT -262.935 90.525 -262.765 90.695 ;
        RECT -262.475 90.525 -262.305 90.695 ;
        RECT -262.015 90.525 -261.845 90.695 ;
        RECT -261.555 90.525 -261.385 90.695 ;
        RECT -261.095 90.525 -260.925 90.695 ;
        RECT -260.635 90.525 -260.465 90.695 ;
        RECT -260.175 90.525 -260.005 90.695 ;
        RECT -253.015 90.525 -252.845 90.695 ;
        RECT -252.555 90.525 -252.385 90.695 ;
        RECT -252.095 90.525 -251.925 90.695 ;
        RECT -251.635 90.525 -251.465 90.695 ;
        RECT -251.175 90.525 -251.005 90.695 ;
        RECT -250.715 90.525 -250.545 90.695 ;
        RECT -250.255 90.525 -250.085 90.695 ;
        RECT -243.095 90.525 -242.925 90.695 ;
        RECT -242.635 90.525 -242.465 90.695 ;
        RECT -242.175 90.525 -242.005 90.695 ;
        RECT -241.715 90.525 -241.545 90.695 ;
        RECT -241.255 90.525 -241.085 90.695 ;
        RECT -240.795 90.525 -240.625 90.695 ;
        RECT -240.335 90.525 -240.165 90.695 ;
        RECT -233.175 90.525 -233.005 90.695 ;
        RECT -232.715 90.525 -232.545 90.695 ;
        RECT -232.255 90.525 -232.085 90.695 ;
        RECT -231.795 90.525 -231.625 90.695 ;
        RECT -231.335 90.525 -231.165 90.695 ;
        RECT -230.875 90.525 -230.705 90.695 ;
        RECT -230.415 90.525 -230.245 90.695 ;
        RECT -223.255 90.525 -223.085 90.695 ;
        RECT -222.795 90.525 -222.625 90.695 ;
        RECT -222.335 90.525 -222.165 90.695 ;
        RECT -221.875 90.525 -221.705 90.695 ;
        RECT -221.415 90.525 -221.245 90.695 ;
        RECT -220.955 90.525 -220.785 90.695 ;
        RECT -220.495 90.525 -220.325 90.695 ;
        RECT -213.335 90.525 -213.165 90.695 ;
        RECT -212.875 90.525 -212.705 90.695 ;
        RECT -212.415 90.525 -212.245 90.695 ;
        RECT -211.955 90.525 -211.785 90.695 ;
        RECT -211.495 90.525 -211.325 90.695 ;
        RECT -211.035 90.525 -210.865 90.695 ;
        RECT -210.575 90.525 -210.405 90.695 ;
        RECT -203.415 90.525 -203.245 90.695 ;
        RECT -202.955 90.525 -202.785 90.695 ;
        RECT -202.495 90.525 -202.325 90.695 ;
        RECT -202.035 90.525 -201.865 90.695 ;
        RECT -201.575 90.525 -201.405 90.695 ;
        RECT -201.115 90.525 -200.945 90.695 ;
        RECT -200.655 90.525 -200.485 90.695 ;
        RECT -193.495 90.525 -193.325 90.695 ;
        RECT -193.035 90.525 -192.865 90.695 ;
        RECT -192.575 90.525 -192.405 90.695 ;
        RECT -192.115 90.525 -191.945 90.695 ;
        RECT -191.655 90.525 -191.485 90.695 ;
        RECT -191.195 90.525 -191.025 90.695 ;
        RECT -190.735 90.525 -190.565 90.695 ;
        RECT -183.575 90.525 -183.405 90.695 ;
        RECT -183.115 90.525 -182.945 90.695 ;
        RECT -182.655 90.525 -182.485 90.695 ;
        RECT -182.195 90.525 -182.025 90.695 ;
        RECT -181.735 90.525 -181.565 90.695 ;
        RECT -181.275 90.525 -181.105 90.695 ;
        RECT -180.815 90.525 -180.645 90.695 ;
        RECT -173.655 90.525 -173.485 90.695 ;
        RECT -173.195 90.525 -173.025 90.695 ;
        RECT -172.735 90.525 -172.565 90.695 ;
        RECT -172.275 90.525 -172.105 90.695 ;
        RECT -171.815 90.525 -171.645 90.695 ;
        RECT -171.355 90.525 -171.185 90.695 ;
        RECT -170.895 90.525 -170.725 90.695 ;
        RECT -163.735 90.525 -163.565 90.695 ;
        RECT -163.275 90.525 -163.105 90.695 ;
        RECT -162.815 90.525 -162.645 90.695 ;
        RECT -162.355 90.525 -162.185 90.695 ;
        RECT -161.895 90.525 -161.725 90.695 ;
        RECT -161.435 90.525 -161.265 90.695 ;
        RECT -160.975 90.525 -160.805 90.695 ;
        RECT -153.815 90.525 -153.645 90.695 ;
        RECT -153.355 90.525 -153.185 90.695 ;
        RECT -152.895 90.525 -152.725 90.695 ;
        RECT -152.435 90.525 -152.265 90.695 ;
        RECT -151.975 90.525 -151.805 90.695 ;
        RECT -151.515 90.525 -151.345 90.695 ;
        RECT -151.055 90.525 -150.885 90.695 ;
        RECT -143.895 90.525 -143.725 90.695 ;
        RECT -143.435 90.525 -143.265 90.695 ;
        RECT -142.975 90.525 -142.805 90.695 ;
        RECT -142.515 90.525 -142.345 90.695 ;
        RECT -142.055 90.525 -141.885 90.695 ;
        RECT -141.595 90.525 -141.425 90.695 ;
        RECT -141.135 90.525 -140.965 90.695 ;
        RECT -133.975 90.525 -133.805 90.695 ;
        RECT -133.515 90.525 -133.345 90.695 ;
        RECT -133.055 90.525 -132.885 90.695 ;
        RECT -132.595 90.525 -132.425 90.695 ;
        RECT -132.135 90.525 -131.965 90.695 ;
        RECT -131.675 90.525 -131.505 90.695 ;
        RECT -131.215 90.525 -131.045 90.695 ;
        RECT -124.055 90.525 -123.885 90.695 ;
        RECT -123.595 90.525 -123.425 90.695 ;
        RECT -123.135 90.525 -122.965 90.695 ;
        RECT -122.675 90.525 -122.505 90.695 ;
        RECT -122.215 90.525 -122.045 90.695 ;
        RECT -121.755 90.525 -121.585 90.695 ;
        RECT -121.295 90.525 -121.125 90.695 ;
        RECT -114.135 90.525 -113.965 90.695 ;
        RECT -113.675 90.525 -113.505 90.695 ;
        RECT -113.215 90.525 -113.045 90.695 ;
        RECT -112.755 90.525 -112.585 90.695 ;
        RECT -112.295 90.525 -112.125 90.695 ;
        RECT -111.835 90.525 -111.665 90.695 ;
        RECT -111.375 90.525 -111.205 90.695 ;
        RECT -104.215 90.525 -104.045 90.695 ;
        RECT -103.755 90.525 -103.585 90.695 ;
        RECT -103.295 90.525 -103.125 90.695 ;
        RECT -102.835 90.525 -102.665 90.695 ;
        RECT -102.375 90.525 -102.205 90.695 ;
        RECT -101.915 90.525 -101.745 90.695 ;
        RECT -101.455 90.525 -101.285 90.695 ;
        RECT -94.295 90.525 -94.125 90.695 ;
        RECT -93.835 90.525 -93.665 90.695 ;
        RECT -93.375 90.525 -93.205 90.695 ;
        RECT -92.915 90.525 -92.745 90.695 ;
        RECT -92.455 90.525 -92.285 90.695 ;
        RECT -91.995 90.525 -91.825 90.695 ;
        RECT -91.535 90.525 -91.365 90.695 ;
        RECT -84.375 90.525 -84.205 90.695 ;
        RECT -83.915 90.525 -83.745 90.695 ;
        RECT -83.455 90.525 -83.285 90.695 ;
        RECT -82.995 90.525 -82.825 90.695 ;
        RECT -82.535 90.525 -82.365 90.695 ;
        RECT -82.075 90.525 -81.905 90.695 ;
        RECT -81.615 90.525 -81.445 90.695 ;
        RECT -74.455 90.525 -74.285 90.695 ;
        RECT -73.995 90.525 -73.825 90.695 ;
        RECT -73.535 90.525 -73.365 90.695 ;
        RECT -73.075 90.525 -72.905 90.695 ;
        RECT -72.615 90.525 -72.445 90.695 ;
        RECT -72.155 90.525 -71.985 90.695 ;
        RECT -71.695 90.525 -71.525 90.695 ;
        RECT -64.535 90.525 -64.365 90.695 ;
        RECT -64.075 90.525 -63.905 90.695 ;
        RECT -63.615 90.525 -63.445 90.695 ;
        RECT -63.155 90.525 -62.985 90.695 ;
        RECT -62.695 90.525 -62.525 90.695 ;
        RECT -62.235 90.525 -62.065 90.695 ;
        RECT -61.775 90.525 -61.605 90.695 ;
        RECT -54.615 90.525 -54.445 90.695 ;
        RECT -54.155 90.525 -53.985 90.695 ;
        RECT -53.695 90.525 -53.525 90.695 ;
        RECT -53.235 90.525 -53.065 90.695 ;
        RECT -52.775 90.525 -52.605 90.695 ;
        RECT -52.315 90.525 -52.145 90.695 ;
        RECT -51.855 90.525 -51.685 90.695 ;
        RECT -44.695 90.525 -44.525 90.695 ;
        RECT -44.235 90.525 -44.065 90.695 ;
        RECT -43.775 90.525 -43.605 90.695 ;
        RECT -43.315 90.525 -43.145 90.695 ;
        RECT -42.855 90.525 -42.685 90.695 ;
        RECT -42.395 90.525 -42.225 90.695 ;
        RECT -41.935 90.525 -41.765 90.695 ;
        RECT -34.775 90.525 -34.605 90.695 ;
        RECT -34.315 90.525 -34.145 90.695 ;
        RECT -33.855 90.525 -33.685 90.695 ;
        RECT -33.395 90.525 -33.225 90.695 ;
        RECT -32.935 90.525 -32.765 90.695 ;
        RECT -32.475 90.525 -32.305 90.695 ;
        RECT -32.015 90.525 -31.845 90.695 ;
        RECT -24.855 90.525 -24.685 90.695 ;
        RECT -24.395 90.525 -24.225 90.695 ;
        RECT -23.935 90.525 -23.765 90.695 ;
        RECT -23.475 90.525 -23.305 90.695 ;
        RECT -23.015 90.525 -22.845 90.695 ;
        RECT -22.555 90.525 -22.385 90.695 ;
        RECT -22.095 90.525 -21.925 90.695 ;
        RECT -14.935 90.525 -14.765 90.695 ;
        RECT -14.475 90.525 -14.305 90.695 ;
        RECT -14.015 90.525 -13.845 90.695 ;
        RECT -13.555 90.525 -13.385 90.695 ;
        RECT -13.095 90.525 -12.925 90.695 ;
        RECT -12.635 90.525 -12.465 90.695 ;
        RECT -12.175 90.525 -12.005 90.695 ;
        RECT -5.015 90.525 -4.845 90.695 ;
        RECT -4.555 90.525 -4.385 90.695 ;
        RECT -4.095 90.525 -3.925 90.695 ;
        RECT -3.635 90.525 -3.465 90.695 ;
        RECT -3.175 90.525 -3.005 90.695 ;
        RECT -2.715 90.525 -2.545 90.695 ;
        RECT -2.255 90.525 -2.085 90.695 ;
        RECT 4.905 90.525 5.075 90.695 ;
        RECT 5.365 90.525 5.535 90.695 ;
        RECT 5.825 90.525 5.995 90.695 ;
        RECT 6.285 90.525 6.455 90.695 ;
        RECT 6.745 90.525 6.915 90.695 ;
        RECT 7.205 90.525 7.375 90.695 ;
        RECT 7.665 90.525 7.835 90.695 ;
        RECT 14.825 90.525 14.995 90.695 ;
        RECT 15.285 90.525 15.455 90.695 ;
        RECT 15.745 90.525 15.915 90.695 ;
        RECT 16.205 90.525 16.375 90.695 ;
        RECT 16.665 90.525 16.835 90.695 ;
        RECT 17.125 90.525 17.295 90.695 ;
        RECT 17.585 90.525 17.755 90.695 ;
        RECT 24.745 90.525 24.915 90.695 ;
        RECT 25.205 90.525 25.375 90.695 ;
        RECT 25.665 90.525 25.835 90.695 ;
        RECT 26.125 90.525 26.295 90.695 ;
        RECT -286.825 89.865 -286.655 90.035 ;
        RECT -286.355 89.940 -286.185 90.110 ;
        RECT -286.825 89.405 -286.655 89.575 ;
        RECT -286.825 88.945 -286.655 89.115 ;
        RECT -285.885 89.865 -285.715 90.035 ;
        RECT -276.905 89.865 -276.735 90.035 ;
        RECT -276.435 89.940 -276.265 90.110 ;
        RECT -285.885 89.405 -285.715 89.575 ;
        RECT -276.905 89.405 -276.735 89.575 ;
        RECT -285.885 88.945 -285.715 89.115 ;
        RECT -276.905 88.945 -276.735 89.115 ;
        RECT -275.965 89.865 -275.795 90.035 ;
        RECT -266.985 89.865 -266.815 90.035 ;
        RECT -266.515 89.940 -266.345 90.110 ;
        RECT -275.965 89.405 -275.795 89.575 ;
        RECT -266.985 89.405 -266.815 89.575 ;
        RECT -275.965 88.945 -275.795 89.115 ;
        RECT -266.985 88.945 -266.815 89.115 ;
        RECT -266.045 89.865 -265.875 90.035 ;
        RECT -257.065 89.865 -256.895 90.035 ;
        RECT -256.595 89.940 -256.425 90.110 ;
        RECT -266.045 89.405 -265.875 89.575 ;
        RECT -257.065 89.405 -256.895 89.575 ;
        RECT -266.045 88.945 -265.875 89.115 ;
        RECT -257.065 88.945 -256.895 89.115 ;
        RECT -256.125 89.865 -255.955 90.035 ;
        RECT -247.145 89.865 -246.975 90.035 ;
        RECT -246.675 89.940 -246.505 90.110 ;
        RECT -256.125 89.405 -255.955 89.575 ;
        RECT -247.145 89.405 -246.975 89.575 ;
        RECT -256.125 88.945 -255.955 89.115 ;
        RECT -247.145 88.945 -246.975 89.115 ;
        RECT -246.205 89.865 -246.035 90.035 ;
        RECT -237.225 89.865 -237.055 90.035 ;
        RECT -236.755 89.940 -236.585 90.110 ;
        RECT -246.205 89.405 -246.035 89.575 ;
        RECT -237.225 89.405 -237.055 89.575 ;
        RECT -246.205 88.945 -246.035 89.115 ;
        RECT -237.225 88.945 -237.055 89.115 ;
        RECT -236.285 89.865 -236.115 90.035 ;
        RECT -227.305 89.865 -227.135 90.035 ;
        RECT -226.835 89.940 -226.665 90.110 ;
        RECT -236.285 89.405 -236.115 89.575 ;
        RECT -227.305 89.405 -227.135 89.575 ;
        RECT -236.285 88.945 -236.115 89.115 ;
        RECT -227.305 88.945 -227.135 89.115 ;
        RECT -226.365 89.865 -226.195 90.035 ;
        RECT -217.385 89.865 -217.215 90.035 ;
        RECT -216.915 89.940 -216.745 90.110 ;
        RECT -226.365 89.405 -226.195 89.575 ;
        RECT -217.385 89.405 -217.215 89.575 ;
        RECT -226.365 88.945 -226.195 89.115 ;
        RECT -217.385 88.945 -217.215 89.115 ;
        RECT -216.445 89.865 -216.275 90.035 ;
        RECT -207.465 89.865 -207.295 90.035 ;
        RECT -206.995 89.940 -206.825 90.110 ;
        RECT -216.445 89.405 -216.275 89.575 ;
        RECT -207.465 89.405 -207.295 89.575 ;
        RECT -216.445 88.945 -216.275 89.115 ;
        RECT -207.465 88.945 -207.295 89.115 ;
        RECT -206.525 89.865 -206.355 90.035 ;
        RECT -197.545 89.865 -197.375 90.035 ;
        RECT -197.075 89.940 -196.905 90.110 ;
        RECT -206.525 89.405 -206.355 89.575 ;
        RECT -197.545 89.405 -197.375 89.575 ;
        RECT -206.525 88.945 -206.355 89.115 ;
        RECT -197.545 88.945 -197.375 89.115 ;
        RECT -196.605 89.865 -196.435 90.035 ;
        RECT -187.625 89.865 -187.455 90.035 ;
        RECT -187.155 89.940 -186.985 90.110 ;
        RECT -196.605 89.405 -196.435 89.575 ;
        RECT -187.625 89.405 -187.455 89.575 ;
        RECT -196.605 88.945 -196.435 89.115 ;
        RECT -187.625 88.945 -187.455 89.115 ;
        RECT -186.685 89.865 -186.515 90.035 ;
        RECT -177.705 89.865 -177.535 90.035 ;
        RECT -177.235 89.940 -177.065 90.110 ;
        RECT -186.685 89.405 -186.515 89.575 ;
        RECT -177.705 89.405 -177.535 89.575 ;
        RECT -186.685 88.945 -186.515 89.115 ;
        RECT -177.705 88.945 -177.535 89.115 ;
        RECT -176.765 89.865 -176.595 90.035 ;
        RECT -167.785 89.865 -167.615 90.035 ;
        RECT -167.315 89.940 -167.145 90.110 ;
        RECT -176.765 89.405 -176.595 89.575 ;
        RECT -167.785 89.405 -167.615 89.575 ;
        RECT -176.765 88.945 -176.595 89.115 ;
        RECT -167.785 88.945 -167.615 89.115 ;
        RECT -166.845 89.865 -166.675 90.035 ;
        RECT -157.865 89.865 -157.695 90.035 ;
        RECT -157.395 89.940 -157.225 90.110 ;
        RECT -166.845 89.405 -166.675 89.575 ;
        RECT -157.865 89.405 -157.695 89.575 ;
        RECT -166.845 88.945 -166.675 89.115 ;
        RECT -157.865 88.945 -157.695 89.115 ;
        RECT -156.925 89.865 -156.755 90.035 ;
        RECT -147.945 89.865 -147.775 90.035 ;
        RECT -147.475 89.940 -147.305 90.110 ;
        RECT -156.925 89.405 -156.755 89.575 ;
        RECT -147.945 89.405 -147.775 89.575 ;
        RECT -156.925 88.945 -156.755 89.115 ;
        RECT -147.945 88.945 -147.775 89.115 ;
        RECT -147.005 89.865 -146.835 90.035 ;
        RECT -138.025 89.865 -137.855 90.035 ;
        RECT -137.555 89.940 -137.385 90.110 ;
        RECT -147.005 89.405 -146.835 89.575 ;
        RECT -138.025 89.405 -137.855 89.575 ;
        RECT -147.005 88.945 -146.835 89.115 ;
        RECT -138.025 88.945 -137.855 89.115 ;
        RECT -137.085 89.865 -136.915 90.035 ;
        RECT -128.105 89.865 -127.935 90.035 ;
        RECT -127.635 89.940 -127.465 90.110 ;
        RECT -137.085 89.405 -136.915 89.575 ;
        RECT -128.105 89.405 -127.935 89.575 ;
        RECT -137.085 88.945 -136.915 89.115 ;
        RECT -128.105 88.945 -127.935 89.115 ;
        RECT -127.165 89.865 -126.995 90.035 ;
        RECT -118.185 89.865 -118.015 90.035 ;
        RECT -117.715 89.940 -117.545 90.110 ;
        RECT -127.165 89.405 -126.995 89.575 ;
        RECT -118.185 89.405 -118.015 89.575 ;
        RECT -127.165 88.945 -126.995 89.115 ;
        RECT -118.185 88.945 -118.015 89.115 ;
        RECT -117.245 89.865 -117.075 90.035 ;
        RECT -108.265 89.865 -108.095 90.035 ;
        RECT -107.795 89.940 -107.625 90.110 ;
        RECT -117.245 89.405 -117.075 89.575 ;
        RECT -108.265 89.405 -108.095 89.575 ;
        RECT -117.245 88.945 -117.075 89.115 ;
        RECT -108.265 88.945 -108.095 89.115 ;
        RECT -107.325 89.865 -107.155 90.035 ;
        RECT -98.345 89.865 -98.175 90.035 ;
        RECT -97.875 89.940 -97.705 90.110 ;
        RECT -107.325 89.405 -107.155 89.575 ;
        RECT -98.345 89.405 -98.175 89.575 ;
        RECT -107.325 88.945 -107.155 89.115 ;
        RECT -98.345 88.945 -98.175 89.115 ;
        RECT -97.405 89.865 -97.235 90.035 ;
        RECT -88.425 89.865 -88.255 90.035 ;
        RECT -87.955 89.940 -87.785 90.110 ;
        RECT -97.405 89.405 -97.235 89.575 ;
        RECT -88.425 89.405 -88.255 89.575 ;
        RECT -97.405 88.945 -97.235 89.115 ;
        RECT -88.425 88.945 -88.255 89.115 ;
        RECT -87.485 89.865 -87.315 90.035 ;
        RECT -78.505 89.865 -78.335 90.035 ;
        RECT -78.035 89.940 -77.865 90.110 ;
        RECT -87.485 89.405 -87.315 89.575 ;
        RECT -78.505 89.405 -78.335 89.575 ;
        RECT -87.485 88.945 -87.315 89.115 ;
        RECT -78.505 88.945 -78.335 89.115 ;
        RECT -77.565 89.865 -77.395 90.035 ;
        RECT -68.585 89.865 -68.415 90.035 ;
        RECT -68.115 89.940 -67.945 90.110 ;
        RECT -77.565 89.405 -77.395 89.575 ;
        RECT -68.585 89.405 -68.415 89.575 ;
        RECT -77.565 88.945 -77.395 89.115 ;
        RECT -68.585 88.945 -68.415 89.115 ;
        RECT -67.645 89.865 -67.475 90.035 ;
        RECT -58.665 89.865 -58.495 90.035 ;
        RECT -58.195 89.940 -58.025 90.110 ;
        RECT -67.645 89.405 -67.475 89.575 ;
        RECT -58.665 89.405 -58.495 89.575 ;
        RECT -67.645 88.945 -67.475 89.115 ;
        RECT -58.665 88.945 -58.495 89.115 ;
        RECT -57.725 89.865 -57.555 90.035 ;
        RECT -48.745 89.865 -48.575 90.035 ;
        RECT -48.275 89.940 -48.105 90.110 ;
        RECT -57.725 89.405 -57.555 89.575 ;
        RECT -48.745 89.405 -48.575 89.575 ;
        RECT -57.725 88.945 -57.555 89.115 ;
        RECT -48.745 88.945 -48.575 89.115 ;
        RECT -47.805 89.865 -47.635 90.035 ;
        RECT -38.825 89.865 -38.655 90.035 ;
        RECT -38.355 89.940 -38.185 90.110 ;
        RECT -47.805 89.405 -47.635 89.575 ;
        RECT -38.825 89.405 -38.655 89.575 ;
        RECT -47.805 88.945 -47.635 89.115 ;
        RECT -38.825 88.945 -38.655 89.115 ;
        RECT -37.885 89.865 -37.715 90.035 ;
        RECT -28.905 89.865 -28.735 90.035 ;
        RECT -28.435 89.940 -28.265 90.110 ;
        RECT -37.885 89.405 -37.715 89.575 ;
        RECT -28.905 89.405 -28.735 89.575 ;
        RECT -37.885 88.945 -37.715 89.115 ;
        RECT -28.905 88.945 -28.735 89.115 ;
        RECT -27.965 89.865 -27.795 90.035 ;
        RECT -18.985 89.865 -18.815 90.035 ;
        RECT -18.515 89.940 -18.345 90.110 ;
        RECT -27.965 89.405 -27.795 89.575 ;
        RECT -18.985 89.405 -18.815 89.575 ;
        RECT -27.965 88.945 -27.795 89.115 ;
        RECT -18.985 88.945 -18.815 89.115 ;
        RECT -18.045 89.865 -17.875 90.035 ;
        RECT -9.065 89.865 -8.895 90.035 ;
        RECT -8.595 89.940 -8.425 90.110 ;
        RECT -18.045 89.405 -17.875 89.575 ;
        RECT -9.065 89.405 -8.895 89.575 ;
        RECT -18.045 88.945 -17.875 89.115 ;
        RECT -9.065 88.945 -8.895 89.115 ;
        RECT -8.125 89.865 -7.955 90.035 ;
        RECT 0.855 89.865 1.025 90.035 ;
        RECT 1.325 89.940 1.495 90.110 ;
        RECT -8.125 89.405 -7.955 89.575 ;
        RECT 0.855 89.405 1.025 89.575 ;
        RECT -8.125 88.945 -7.955 89.115 ;
        RECT 0.855 88.945 1.025 89.115 ;
        RECT 1.795 89.865 1.965 90.035 ;
        RECT 10.775 89.865 10.945 90.035 ;
        RECT 11.245 89.940 11.415 90.110 ;
        RECT 1.795 89.405 1.965 89.575 ;
        RECT 10.775 89.405 10.945 89.575 ;
        RECT 1.795 88.945 1.965 89.115 ;
        RECT 10.775 88.945 10.945 89.115 ;
        RECT 11.715 89.865 11.885 90.035 ;
        RECT 20.695 89.865 20.865 90.035 ;
        RECT 21.165 89.940 21.335 90.110 ;
        RECT 11.715 89.405 11.885 89.575 ;
        RECT 20.695 89.405 20.865 89.575 ;
        RECT 11.715 88.945 11.885 89.115 ;
        RECT 20.695 88.945 20.865 89.115 ;
        RECT 21.635 89.865 21.805 90.035 ;
        RECT 21.635 89.405 21.805 89.575 ;
        RECT 21.635 88.945 21.805 89.115 ;
        RECT -281.615 7.115 -281.445 7.285 ;
        RECT -281.145 7.110 -280.975 7.280 ;
        RECT -280.675 7.115 -280.505 7.285 ;
        RECT -281.615 6.655 -281.445 6.825 ;
        RECT -281.615 6.195 -281.445 6.365 ;
        RECT -271.695 7.115 -271.525 7.285 ;
        RECT -271.225 7.110 -271.055 7.280 ;
        RECT -270.755 7.115 -270.585 7.285 ;
        RECT -280.675 6.655 -280.505 6.825 ;
        RECT -271.695 6.655 -271.525 6.825 ;
        RECT -280.675 6.195 -280.505 6.365 ;
        RECT -271.695 6.195 -271.525 6.365 ;
        RECT -261.775 7.115 -261.605 7.285 ;
        RECT -261.305 7.110 -261.135 7.280 ;
        RECT -260.835 7.115 -260.665 7.285 ;
        RECT -270.755 6.655 -270.585 6.825 ;
        RECT -261.775 6.655 -261.605 6.825 ;
        RECT -270.755 6.195 -270.585 6.365 ;
        RECT -261.775 6.195 -261.605 6.365 ;
        RECT -251.855 7.115 -251.685 7.285 ;
        RECT -251.385 7.110 -251.215 7.280 ;
        RECT -250.915 7.115 -250.745 7.285 ;
        RECT -260.835 6.655 -260.665 6.825 ;
        RECT -251.855 6.655 -251.685 6.825 ;
        RECT -260.835 6.195 -260.665 6.365 ;
        RECT -251.855 6.195 -251.685 6.365 ;
        RECT -241.935 7.115 -241.765 7.285 ;
        RECT -241.465 7.110 -241.295 7.280 ;
        RECT -240.995 7.115 -240.825 7.285 ;
        RECT -250.915 6.655 -250.745 6.825 ;
        RECT -241.935 6.655 -241.765 6.825 ;
        RECT -250.915 6.195 -250.745 6.365 ;
        RECT -241.935 6.195 -241.765 6.365 ;
        RECT -232.015 7.115 -231.845 7.285 ;
        RECT -231.545 7.110 -231.375 7.280 ;
        RECT -231.075 7.115 -230.905 7.285 ;
        RECT -240.995 6.655 -240.825 6.825 ;
        RECT -232.015 6.655 -231.845 6.825 ;
        RECT -240.995 6.195 -240.825 6.365 ;
        RECT -232.015 6.195 -231.845 6.365 ;
        RECT -222.095 7.115 -221.925 7.285 ;
        RECT -221.625 7.110 -221.455 7.280 ;
        RECT -221.155 7.115 -220.985 7.285 ;
        RECT -231.075 6.655 -230.905 6.825 ;
        RECT -222.095 6.655 -221.925 6.825 ;
        RECT -231.075 6.195 -230.905 6.365 ;
        RECT -222.095 6.195 -221.925 6.365 ;
        RECT -212.175 7.115 -212.005 7.285 ;
        RECT -211.705 7.110 -211.535 7.280 ;
        RECT -211.235 7.115 -211.065 7.285 ;
        RECT -221.155 6.655 -220.985 6.825 ;
        RECT -212.175 6.655 -212.005 6.825 ;
        RECT -221.155 6.195 -220.985 6.365 ;
        RECT -212.175 6.195 -212.005 6.365 ;
        RECT -202.255 7.115 -202.085 7.285 ;
        RECT -201.785 7.110 -201.615 7.280 ;
        RECT -201.315 7.115 -201.145 7.285 ;
        RECT -211.235 6.655 -211.065 6.825 ;
        RECT -202.255 6.655 -202.085 6.825 ;
        RECT -211.235 6.195 -211.065 6.365 ;
        RECT -202.255 6.195 -202.085 6.365 ;
        RECT -192.335 7.115 -192.165 7.285 ;
        RECT -191.865 7.110 -191.695 7.280 ;
        RECT -191.395 7.115 -191.225 7.285 ;
        RECT -201.315 6.655 -201.145 6.825 ;
        RECT -192.335 6.655 -192.165 6.825 ;
        RECT -201.315 6.195 -201.145 6.365 ;
        RECT -192.335 6.195 -192.165 6.365 ;
        RECT -182.415 7.115 -182.245 7.285 ;
        RECT -181.945 7.110 -181.775 7.280 ;
        RECT -181.475 7.115 -181.305 7.285 ;
        RECT -191.395 6.655 -191.225 6.825 ;
        RECT -182.415 6.655 -182.245 6.825 ;
        RECT -191.395 6.195 -191.225 6.365 ;
        RECT -182.415 6.195 -182.245 6.365 ;
        RECT -172.495 7.115 -172.325 7.285 ;
        RECT -172.025 7.110 -171.855 7.280 ;
        RECT -171.555 7.115 -171.385 7.285 ;
        RECT -181.475 6.655 -181.305 6.825 ;
        RECT -172.495 6.655 -172.325 6.825 ;
        RECT -181.475 6.195 -181.305 6.365 ;
        RECT -172.495 6.195 -172.325 6.365 ;
        RECT -162.575 7.115 -162.405 7.285 ;
        RECT -162.105 7.110 -161.935 7.280 ;
        RECT -161.635 7.115 -161.465 7.285 ;
        RECT -171.555 6.655 -171.385 6.825 ;
        RECT -162.575 6.655 -162.405 6.825 ;
        RECT -171.555 6.195 -171.385 6.365 ;
        RECT -162.575 6.195 -162.405 6.365 ;
        RECT -152.655 7.115 -152.485 7.285 ;
        RECT -152.185 7.110 -152.015 7.280 ;
        RECT -151.715 7.115 -151.545 7.285 ;
        RECT -161.635 6.655 -161.465 6.825 ;
        RECT -152.655 6.655 -152.485 6.825 ;
        RECT -161.635 6.195 -161.465 6.365 ;
        RECT -152.655 6.195 -152.485 6.365 ;
        RECT -142.735 7.115 -142.565 7.285 ;
        RECT -142.265 7.110 -142.095 7.280 ;
        RECT -141.795 7.115 -141.625 7.285 ;
        RECT -151.715 6.655 -151.545 6.825 ;
        RECT -142.735 6.655 -142.565 6.825 ;
        RECT -151.715 6.195 -151.545 6.365 ;
        RECT -142.735 6.195 -142.565 6.365 ;
        RECT -132.815 7.115 -132.645 7.285 ;
        RECT -132.345 7.110 -132.175 7.280 ;
        RECT -131.875 7.115 -131.705 7.285 ;
        RECT -141.795 6.655 -141.625 6.825 ;
        RECT -132.815 6.655 -132.645 6.825 ;
        RECT -141.795 6.195 -141.625 6.365 ;
        RECT -132.815 6.195 -132.645 6.365 ;
        RECT -122.895 7.115 -122.725 7.285 ;
        RECT -122.425 7.110 -122.255 7.280 ;
        RECT -121.955 7.115 -121.785 7.285 ;
        RECT -131.875 6.655 -131.705 6.825 ;
        RECT -122.895 6.655 -122.725 6.825 ;
        RECT -131.875 6.195 -131.705 6.365 ;
        RECT -122.895 6.195 -122.725 6.365 ;
        RECT -112.975 7.115 -112.805 7.285 ;
        RECT -112.505 7.110 -112.335 7.280 ;
        RECT -112.035 7.115 -111.865 7.285 ;
        RECT -121.955 6.655 -121.785 6.825 ;
        RECT -112.975 6.655 -112.805 6.825 ;
        RECT -121.955 6.195 -121.785 6.365 ;
        RECT -112.975 6.195 -112.805 6.365 ;
        RECT -103.055 7.115 -102.885 7.285 ;
        RECT -102.585 7.110 -102.415 7.280 ;
        RECT -102.115 7.115 -101.945 7.285 ;
        RECT -112.035 6.655 -111.865 6.825 ;
        RECT -103.055 6.655 -102.885 6.825 ;
        RECT -112.035 6.195 -111.865 6.365 ;
        RECT -103.055 6.195 -102.885 6.365 ;
        RECT -93.135 7.115 -92.965 7.285 ;
        RECT -92.665 7.110 -92.495 7.280 ;
        RECT -92.195 7.115 -92.025 7.285 ;
        RECT -102.115 6.655 -101.945 6.825 ;
        RECT -93.135 6.655 -92.965 6.825 ;
        RECT -102.115 6.195 -101.945 6.365 ;
        RECT -93.135 6.195 -92.965 6.365 ;
        RECT -83.215 7.115 -83.045 7.285 ;
        RECT -82.745 7.110 -82.575 7.280 ;
        RECT -82.275 7.115 -82.105 7.285 ;
        RECT -92.195 6.655 -92.025 6.825 ;
        RECT -83.215 6.655 -83.045 6.825 ;
        RECT -92.195 6.195 -92.025 6.365 ;
        RECT -83.215 6.195 -83.045 6.365 ;
        RECT -73.295 7.115 -73.125 7.285 ;
        RECT -72.825 7.110 -72.655 7.280 ;
        RECT -72.355 7.115 -72.185 7.285 ;
        RECT -82.275 6.655 -82.105 6.825 ;
        RECT -73.295 6.655 -73.125 6.825 ;
        RECT -82.275 6.195 -82.105 6.365 ;
        RECT -73.295 6.195 -73.125 6.365 ;
        RECT -63.375 7.115 -63.205 7.285 ;
        RECT -62.905 7.110 -62.735 7.280 ;
        RECT -62.435 7.115 -62.265 7.285 ;
        RECT -72.355 6.655 -72.185 6.825 ;
        RECT -63.375 6.655 -63.205 6.825 ;
        RECT -72.355 6.195 -72.185 6.365 ;
        RECT -63.375 6.195 -63.205 6.365 ;
        RECT -53.455 7.115 -53.285 7.285 ;
        RECT -52.985 7.110 -52.815 7.280 ;
        RECT -52.515 7.115 -52.345 7.285 ;
        RECT -62.435 6.655 -62.265 6.825 ;
        RECT -53.455 6.655 -53.285 6.825 ;
        RECT -62.435 6.195 -62.265 6.365 ;
        RECT -53.455 6.195 -53.285 6.365 ;
        RECT -43.535 7.115 -43.365 7.285 ;
        RECT -43.065 7.110 -42.895 7.280 ;
        RECT -42.595 7.115 -42.425 7.285 ;
        RECT -52.515 6.655 -52.345 6.825 ;
        RECT -43.535 6.655 -43.365 6.825 ;
        RECT -52.515 6.195 -52.345 6.365 ;
        RECT -43.535 6.195 -43.365 6.365 ;
        RECT -33.615 7.115 -33.445 7.285 ;
        RECT -33.145 7.110 -32.975 7.280 ;
        RECT -32.675 7.115 -32.505 7.285 ;
        RECT -42.595 6.655 -42.425 6.825 ;
        RECT -33.615 6.655 -33.445 6.825 ;
        RECT -42.595 6.195 -42.425 6.365 ;
        RECT -33.615 6.195 -33.445 6.365 ;
        RECT -23.695 7.115 -23.525 7.285 ;
        RECT -23.225 7.110 -23.055 7.280 ;
        RECT -22.755 7.115 -22.585 7.285 ;
        RECT -32.675 6.655 -32.505 6.825 ;
        RECT -23.695 6.655 -23.525 6.825 ;
        RECT -32.675 6.195 -32.505 6.365 ;
        RECT -23.695 6.195 -23.525 6.365 ;
        RECT -13.775 7.115 -13.605 7.285 ;
        RECT -13.305 7.110 -13.135 7.280 ;
        RECT -12.835 7.115 -12.665 7.285 ;
        RECT -22.755 6.655 -22.585 6.825 ;
        RECT -13.775 6.655 -13.605 6.825 ;
        RECT -22.755 6.195 -22.585 6.365 ;
        RECT -13.775 6.195 -13.605 6.365 ;
        RECT -3.855 7.115 -3.685 7.285 ;
        RECT -3.385 7.110 -3.215 7.280 ;
        RECT -2.915 7.115 -2.745 7.285 ;
        RECT -12.835 6.655 -12.665 6.825 ;
        RECT -3.855 6.655 -3.685 6.825 ;
        RECT -12.835 6.195 -12.665 6.365 ;
        RECT -3.855 6.195 -3.685 6.365 ;
        RECT 6.065 7.115 6.235 7.285 ;
        RECT 6.535 7.110 6.705 7.280 ;
        RECT 7.005 7.115 7.175 7.285 ;
        RECT -2.915 6.655 -2.745 6.825 ;
        RECT 6.065 6.655 6.235 6.825 ;
        RECT -2.915 6.195 -2.745 6.365 ;
        RECT 6.065 6.195 6.235 6.365 ;
        RECT 15.985 7.115 16.155 7.285 ;
        RECT 16.455 7.110 16.625 7.280 ;
        RECT 16.925 7.115 17.095 7.285 ;
        RECT 7.005 6.655 7.175 6.825 ;
        RECT 15.985 6.655 16.155 6.825 ;
        RECT 7.005 6.195 7.175 6.365 ;
        RECT 15.985 6.195 16.155 6.365 ;
        RECT 25.905 7.115 26.075 7.285 ;
        RECT 26.375 7.110 26.545 7.280 ;
        RECT 16.925 6.655 17.095 6.825 ;
        RECT 25.905 6.655 26.075 6.825 ;
        RECT 16.925 6.195 17.095 6.365 ;
        RECT 25.905 6.195 26.075 6.365 ;
        RECT -287.485 5.535 -287.315 5.705 ;
        RECT -287.025 5.535 -286.855 5.705 ;
        RECT -286.565 5.535 -286.395 5.705 ;
        RECT -286.105 5.535 -285.935 5.705 ;
        RECT -285.645 5.535 -285.475 5.705 ;
        RECT -285.185 5.535 -285.015 5.705 ;
        RECT -284.725 5.535 -284.555 5.705 ;
        RECT -277.565 5.535 -277.395 5.705 ;
        RECT -277.105 5.535 -276.935 5.705 ;
        RECT -276.645 5.535 -276.475 5.705 ;
        RECT -276.185 5.535 -276.015 5.705 ;
        RECT -275.725 5.535 -275.555 5.705 ;
        RECT -275.265 5.535 -275.095 5.705 ;
        RECT -274.805 5.535 -274.635 5.705 ;
        RECT -267.645 5.535 -267.475 5.705 ;
        RECT -267.185 5.535 -267.015 5.705 ;
        RECT -266.725 5.535 -266.555 5.705 ;
        RECT -266.265 5.535 -266.095 5.705 ;
        RECT -265.805 5.535 -265.635 5.705 ;
        RECT -265.345 5.535 -265.175 5.705 ;
        RECT -264.885 5.535 -264.715 5.705 ;
        RECT -257.725 5.535 -257.555 5.705 ;
        RECT -257.265 5.535 -257.095 5.705 ;
        RECT -256.805 5.535 -256.635 5.705 ;
        RECT -256.345 5.535 -256.175 5.705 ;
        RECT -255.885 5.535 -255.715 5.705 ;
        RECT -255.425 5.535 -255.255 5.705 ;
        RECT -254.965 5.535 -254.795 5.705 ;
        RECT -247.805 5.535 -247.635 5.705 ;
        RECT -247.345 5.535 -247.175 5.705 ;
        RECT -246.885 5.535 -246.715 5.705 ;
        RECT -246.425 5.535 -246.255 5.705 ;
        RECT -245.965 5.535 -245.795 5.705 ;
        RECT -245.505 5.535 -245.335 5.705 ;
        RECT -245.045 5.535 -244.875 5.705 ;
        RECT -237.885 5.535 -237.715 5.705 ;
        RECT -237.425 5.535 -237.255 5.705 ;
        RECT -236.965 5.535 -236.795 5.705 ;
        RECT -236.505 5.535 -236.335 5.705 ;
        RECT -236.045 5.535 -235.875 5.705 ;
        RECT -235.585 5.535 -235.415 5.705 ;
        RECT -235.125 5.535 -234.955 5.705 ;
        RECT -227.965 5.535 -227.795 5.705 ;
        RECT -227.505 5.535 -227.335 5.705 ;
        RECT -227.045 5.535 -226.875 5.705 ;
        RECT -226.585 5.535 -226.415 5.705 ;
        RECT -226.125 5.535 -225.955 5.705 ;
        RECT -225.665 5.535 -225.495 5.705 ;
        RECT -225.205 5.535 -225.035 5.705 ;
        RECT -218.045 5.535 -217.875 5.705 ;
        RECT -217.585 5.535 -217.415 5.705 ;
        RECT -217.125 5.535 -216.955 5.705 ;
        RECT -216.665 5.535 -216.495 5.705 ;
        RECT -216.205 5.535 -216.035 5.705 ;
        RECT -215.745 5.535 -215.575 5.705 ;
        RECT -215.285 5.535 -215.115 5.705 ;
        RECT -208.125 5.535 -207.955 5.705 ;
        RECT -207.665 5.535 -207.495 5.705 ;
        RECT -207.205 5.535 -207.035 5.705 ;
        RECT -206.745 5.535 -206.575 5.705 ;
        RECT -206.285 5.535 -206.115 5.705 ;
        RECT -205.825 5.535 -205.655 5.705 ;
        RECT -205.365 5.535 -205.195 5.705 ;
        RECT -198.205 5.535 -198.035 5.705 ;
        RECT -197.745 5.535 -197.575 5.705 ;
        RECT -197.285 5.535 -197.115 5.705 ;
        RECT -196.825 5.535 -196.655 5.705 ;
        RECT -196.365 5.535 -196.195 5.705 ;
        RECT -195.905 5.535 -195.735 5.705 ;
        RECT -195.445 5.535 -195.275 5.705 ;
        RECT -188.285 5.535 -188.115 5.705 ;
        RECT -187.825 5.535 -187.655 5.705 ;
        RECT -187.365 5.535 -187.195 5.705 ;
        RECT -186.905 5.535 -186.735 5.705 ;
        RECT -186.445 5.535 -186.275 5.705 ;
        RECT -185.985 5.535 -185.815 5.705 ;
        RECT -185.525 5.535 -185.355 5.705 ;
        RECT -178.365 5.535 -178.195 5.705 ;
        RECT -177.905 5.535 -177.735 5.705 ;
        RECT -177.445 5.535 -177.275 5.705 ;
        RECT -176.985 5.535 -176.815 5.705 ;
        RECT -176.525 5.535 -176.355 5.705 ;
        RECT -176.065 5.535 -175.895 5.705 ;
        RECT -175.605 5.535 -175.435 5.705 ;
        RECT -168.445 5.535 -168.275 5.705 ;
        RECT -167.985 5.535 -167.815 5.705 ;
        RECT -167.525 5.535 -167.355 5.705 ;
        RECT -167.065 5.535 -166.895 5.705 ;
        RECT -166.605 5.535 -166.435 5.705 ;
        RECT -166.145 5.535 -165.975 5.705 ;
        RECT -165.685 5.535 -165.515 5.705 ;
        RECT -158.525 5.535 -158.355 5.705 ;
        RECT -158.065 5.535 -157.895 5.705 ;
        RECT -157.605 5.535 -157.435 5.705 ;
        RECT -157.145 5.535 -156.975 5.705 ;
        RECT -156.685 5.535 -156.515 5.705 ;
        RECT -156.225 5.535 -156.055 5.705 ;
        RECT -155.765 5.535 -155.595 5.705 ;
        RECT -148.605 5.535 -148.435 5.705 ;
        RECT -148.145 5.535 -147.975 5.705 ;
        RECT -147.685 5.535 -147.515 5.705 ;
        RECT -147.225 5.535 -147.055 5.705 ;
        RECT -146.765 5.535 -146.595 5.705 ;
        RECT -146.305 5.535 -146.135 5.705 ;
        RECT -145.845 5.535 -145.675 5.705 ;
        RECT -138.685 5.535 -138.515 5.705 ;
        RECT -138.225 5.535 -138.055 5.705 ;
        RECT -137.765 5.535 -137.595 5.705 ;
        RECT -137.305 5.535 -137.135 5.705 ;
        RECT -136.845 5.535 -136.675 5.705 ;
        RECT -136.385 5.535 -136.215 5.705 ;
        RECT -135.925 5.535 -135.755 5.705 ;
        RECT -128.765 5.535 -128.595 5.705 ;
        RECT -128.305 5.535 -128.135 5.705 ;
        RECT -127.845 5.535 -127.675 5.705 ;
        RECT -127.385 5.535 -127.215 5.705 ;
        RECT -126.925 5.535 -126.755 5.705 ;
        RECT -126.465 5.535 -126.295 5.705 ;
        RECT -126.005 5.535 -125.835 5.705 ;
        RECT -118.845 5.535 -118.675 5.705 ;
        RECT -118.385 5.535 -118.215 5.705 ;
        RECT -117.925 5.535 -117.755 5.705 ;
        RECT -117.465 5.535 -117.295 5.705 ;
        RECT -117.005 5.535 -116.835 5.705 ;
        RECT -116.545 5.535 -116.375 5.705 ;
        RECT -116.085 5.535 -115.915 5.705 ;
        RECT -108.925 5.535 -108.755 5.705 ;
        RECT -108.465 5.535 -108.295 5.705 ;
        RECT -108.005 5.535 -107.835 5.705 ;
        RECT -107.545 5.535 -107.375 5.705 ;
        RECT -107.085 5.535 -106.915 5.705 ;
        RECT -106.625 5.535 -106.455 5.705 ;
        RECT -106.165 5.535 -105.995 5.705 ;
        RECT -99.005 5.535 -98.835 5.705 ;
        RECT -98.545 5.535 -98.375 5.705 ;
        RECT -98.085 5.535 -97.915 5.705 ;
        RECT -97.625 5.535 -97.455 5.705 ;
        RECT -97.165 5.535 -96.995 5.705 ;
        RECT -96.705 5.535 -96.535 5.705 ;
        RECT -96.245 5.535 -96.075 5.705 ;
        RECT -89.085 5.535 -88.915 5.705 ;
        RECT -88.625 5.535 -88.455 5.705 ;
        RECT -88.165 5.535 -87.995 5.705 ;
        RECT -87.705 5.535 -87.535 5.705 ;
        RECT -87.245 5.535 -87.075 5.705 ;
        RECT -86.785 5.535 -86.615 5.705 ;
        RECT -86.325 5.535 -86.155 5.705 ;
        RECT -79.165 5.535 -78.995 5.705 ;
        RECT -78.705 5.535 -78.535 5.705 ;
        RECT -78.245 5.535 -78.075 5.705 ;
        RECT -77.785 5.535 -77.615 5.705 ;
        RECT -77.325 5.535 -77.155 5.705 ;
        RECT -76.865 5.535 -76.695 5.705 ;
        RECT -76.405 5.535 -76.235 5.705 ;
        RECT -69.245 5.535 -69.075 5.705 ;
        RECT -68.785 5.535 -68.615 5.705 ;
        RECT -68.325 5.535 -68.155 5.705 ;
        RECT -67.865 5.535 -67.695 5.705 ;
        RECT -67.405 5.535 -67.235 5.705 ;
        RECT -66.945 5.535 -66.775 5.705 ;
        RECT -66.485 5.535 -66.315 5.705 ;
        RECT -59.325 5.535 -59.155 5.705 ;
        RECT -58.865 5.535 -58.695 5.705 ;
        RECT -58.405 5.535 -58.235 5.705 ;
        RECT -57.945 5.535 -57.775 5.705 ;
        RECT -57.485 5.535 -57.315 5.705 ;
        RECT -57.025 5.535 -56.855 5.705 ;
        RECT -56.565 5.535 -56.395 5.705 ;
        RECT -49.405 5.535 -49.235 5.705 ;
        RECT -48.945 5.535 -48.775 5.705 ;
        RECT -48.485 5.535 -48.315 5.705 ;
        RECT -48.025 5.535 -47.855 5.705 ;
        RECT -47.565 5.535 -47.395 5.705 ;
        RECT -47.105 5.535 -46.935 5.705 ;
        RECT -46.645 5.535 -46.475 5.705 ;
        RECT -39.485 5.535 -39.315 5.705 ;
        RECT -39.025 5.535 -38.855 5.705 ;
        RECT -38.565 5.535 -38.395 5.705 ;
        RECT -38.105 5.535 -37.935 5.705 ;
        RECT -37.645 5.535 -37.475 5.705 ;
        RECT -37.185 5.535 -37.015 5.705 ;
        RECT -36.725 5.535 -36.555 5.705 ;
        RECT -29.565 5.535 -29.395 5.705 ;
        RECT -29.105 5.535 -28.935 5.705 ;
        RECT -28.645 5.535 -28.475 5.705 ;
        RECT -28.185 5.535 -28.015 5.705 ;
        RECT -27.725 5.535 -27.555 5.705 ;
        RECT -27.265 5.535 -27.095 5.705 ;
        RECT -26.805 5.535 -26.635 5.705 ;
        RECT -19.645 5.535 -19.475 5.705 ;
        RECT -19.185 5.535 -19.015 5.705 ;
        RECT -18.725 5.535 -18.555 5.705 ;
        RECT -18.265 5.535 -18.095 5.705 ;
        RECT -17.805 5.535 -17.635 5.705 ;
        RECT -17.345 5.535 -17.175 5.705 ;
        RECT -16.885 5.535 -16.715 5.705 ;
        RECT -9.725 5.535 -9.555 5.705 ;
        RECT -9.265 5.535 -9.095 5.705 ;
        RECT -8.805 5.535 -8.635 5.705 ;
        RECT -8.345 5.535 -8.175 5.705 ;
        RECT -7.885 5.535 -7.715 5.705 ;
        RECT -7.425 5.535 -7.255 5.705 ;
        RECT -6.965 5.535 -6.795 5.705 ;
        RECT 0.195 5.535 0.365 5.705 ;
        RECT 0.655 5.535 0.825 5.705 ;
        RECT 1.115 5.535 1.285 5.705 ;
        RECT 1.575 5.535 1.745 5.705 ;
        RECT 2.035 5.535 2.205 5.705 ;
        RECT 2.495 5.535 2.665 5.705 ;
        RECT 2.955 5.535 3.125 5.705 ;
        RECT 10.115 5.535 10.285 5.705 ;
        RECT 10.575 5.535 10.745 5.705 ;
        RECT 11.035 5.535 11.205 5.705 ;
        RECT 11.495 5.535 11.665 5.705 ;
        RECT 11.955 5.535 12.125 5.705 ;
        RECT 12.415 5.535 12.585 5.705 ;
        RECT 12.875 5.535 13.045 5.705 ;
        RECT 20.035 5.535 20.205 5.705 ;
        RECT 20.495 5.535 20.665 5.705 ;
        RECT 20.955 5.535 21.125 5.705 ;
        RECT 21.415 5.535 21.585 5.705 ;
        RECT 21.875 5.535 22.045 5.705 ;
        RECT 22.335 5.535 22.505 5.705 ;
        RECT 22.795 5.535 22.965 5.705 ;
        RECT -282.525 2.815 -282.355 2.985 ;
        RECT -282.065 2.815 -281.895 2.985 ;
        RECT -281.605 2.815 -281.435 2.985 ;
        RECT -281.145 2.815 -280.975 2.985 ;
        RECT -280.685 2.815 -280.515 2.985 ;
        RECT -280.225 2.815 -280.055 2.985 ;
        RECT -279.765 2.815 -279.595 2.985 ;
        RECT -272.605 2.815 -272.435 2.985 ;
        RECT -272.145 2.815 -271.975 2.985 ;
        RECT -271.685 2.815 -271.515 2.985 ;
        RECT -271.225 2.815 -271.055 2.985 ;
        RECT -270.765 2.815 -270.595 2.985 ;
        RECT -270.305 2.815 -270.135 2.985 ;
        RECT -269.845 2.815 -269.675 2.985 ;
        RECT -262.685 2.815 -262.515 2.985 ;
        RECT -262.225 2.815 -262.055 2.985 ;
        RECT -261.765 2.815 -261.595 2.985 ;
        RECT -261.305 2.815 -261.135 2.985 ;
        RECT -260.845 2.815 -260.675 2.985 ;
        RECT -260.385 2.815 -260.215 2.985 ;
        RECT -259.925 2.815 -259.755 2.985 ;
        RECT -252.765 2.815 -252.595 2.985 ;
        RECT -252.305 2.815 -252.135 2.985 ;
        RECT -251.845 2.815 -251.675 2.985 ;
        RECT -251.385 2.815 -251.215 2.985 ;
        RECT -250.925 2.815 -250.755 2.985 ;
        RECT -250.465 2.815 -250.295 2.985 ;
        RECT -250.005 2.815 -249.835 2.985 ;
        RECT -242.845 2.815 -242.675 2.985 ;
        RECT -242.385 2.815 -242.215 2.985 ;
        RECT -241.925 2.815 -241.755 2.985 ;
        RECT -241.465 2.815 -241.295 2.985 ;
        RECT -241.005 2.815 -240.835 2.985 ;
        RECT -240.545 2.815 -240.375 2.985 ;
        RECT -240.085 2.815 -239.915 2.985 ;
        RECT -232.925 2.815 -232.755 2.985 ;
        RECT -232.465 2.815 -232.295 2.985 ;
        RECT -232.005 2.815 -231.835 2.985 ;
        RECT -231.545 2.815 -231.375 2.985 ;
        RECT -231.085 2.815 -230.915 2.985 ;
        RECT -230.625 2.815 -230.455 2.985 ;
        RECT -230.165 2.815 -229.995 2.985 ;
        RECT -223.005 2.815 -222.835 2.985 ;
        RECT -222.545 2.815 -222.375 2.985 ;
        RECT -222.085 2.815 -221.915 2.985 ;
        RECT -221.625 2.815 -221.455 2.985 ;
        RECT -221.165 2.815 -220.995 2.985 ;
        RECT -220.705 2.815 -220.535 2.985 ;
        RECT -220.245 2.815 -220.075 2.985 ;
        RECT -213.085 2.815 -212.915 2.985 ;
        RECT -212.625 2.815 -212.455 2.985 ;
        RECT -212.165 2.815 -211.995 2.985 ;
        RECT -211.705 2.815 -211.535 2.985 ;
        RECT -211.245 2.815 -211.075 2.985 ;
        RECT -210.785 2.815 -210.615 2.985 ;
        RECT -210.325 2.815 -210.155 2.985 ;
        RECT -203.165 2.815 -202.995 2.985 ;
        RECT -202.705 2.815 -202.535 2.985 ;
        RECT -202.245 2.815 -202.075 2.985 ;
        RECT -201.785 2.815 -201.615 2.985 ;
        RECT -201.325 2.815 -201.155 2.985 ;
        RECT -200.865 2.815 -200.695 2.985 ;
        RECT -200.405 2.815 -200.235 2.985 ;
        RECT -193.245 2.815 -193.075 2.985 ;
        RECT -192.785 2.815 -192.615 2.985 ;
        RECT -192.325 2.815 -192.155 2.985 ;
        RECT -191.865 2.815 -191.695 2.985 ;
        RECT -191.405 2.815 -191.235 2.985 ;
        RECT -190.945 2.815 -190.775 2.985 ;
        RECT -190.485 2.815 -190.315 2.985 ;
        RECT -183.325 2.815 -183.155 2.985 ;
        RECT -182.865 2.815 -182.695 2.985 ;
        RECT -182.405 2.815 -182.235 2.985 ;
        RECT -181.945 2.815 -181.775 2.985 ;
        RECT -181.485 2.815 -181.315 2.985 ;
        RECT -181.025 2.815 -180.855 2.985 ;
        RECT -180.565 2.815 -180.395 2.985 ;
        RECT -173.405 2.815 -173.235 2.985 ;
        RECT -172.945 2.815 -172.775 2.985 ;
        RECT -172.485 2.815 -172.315 2.985 ;
        RECT -172.025 2.815 -171.855 2.985 ;
        RECT -171.565 2.815 -171.395 2.985 ;
        RECT -171.105 2.815 -170.935 2.985 ;
        RECT -170.645 2.815 -170.475 2.985 ;
        RECT -163.485 2.815 -163.315 2.985 ;
        RECT -163.025 2.815 -162.855 2.985 ;
        RECT -162.565 2.815 -162.395 2.985 ;
        RECT -162.105 2.815 -161.935 2.985 ;
        RECT -161.645 2.815 -161.475 2.985 ;
        RECT -161.185 2.815 -161.015 2.985 ;
        RECT -160.725 2.815 -160.555 2.985 ;
        RECT -153.565 2.815 -153.395 2.985 ;
        RECT -153.105 2.815 -152.935 2.985 ;
        RECT -152.645 2.815 -152.475 2.985 ;
        RECT -152.185 2.815 -152.015 2.985 ;
        RECT -151.725 2.815 -151.555 2.985 ;
        RECT -151.265 2.815 -151.095 2.985 ;
        RECT -150.805 2.815 -150.635 2.985 ;
        RECT -143.645 2.815 -143.475 2.985 ;
        RECT -143.185 2.815 -143.015 2.985 ;
        RECT -142.725 2.815 -142.555 2.985 ;
        RECT -142.265 2.815 -142.095 2.985 ;
        RECT -141.805 2.815 -141.635 2.985 ;
        RECT -141.345 2.815 -141.175 2.985 ;
        RECT -140.885 2.815 -140.715 2.985 ;
        RECT -133.725 2.815 -133.555 2.985 ;
        RECT -133.265 2.815 -133.095 2.985 ;
        RECT -132.805 2.815 -132.635 2.985 ;
        RECT -132.345 2.815 -132.175 2.985 ;
        RECT -131.885 2.815 -131.715 2.985 ;
        RECT -131.425 2.815 -131.255 2.985 ;
        RECT -130.965 2.815 -130.795 2.985 ;
        RECT -123.805 2.815 -123.635 2.985 ;
        RECT -123.345 2.815 -123.175 2.985 ;
        RECT -122.885 2.815 -122.715 2.985 ;
        RECT -122.425 2.815 -122.255 2.985 ;
        RECT -121.965 2.815 -121.795 2.985 ;
        RECT -121.505 2.815 -121.335 2.985 ;
        RECT -121.045 2.815 -120.875 2.985 ;
        RECT -113.885 2.815 -113.715 2.985 ;
        RECT -113.425 2.815 -113.255 2.985 ;
        RECT -112.965 2.815 -112.795 2.985 ;
        RECT -112.505 2.815 -112.335 2.985 ;
        RECT -112.045 2.815 -111.875 2.985 ;
        RECT -111.585 2.815 -111.415 2.985 ;
        RECT -111.125 2.815 -110.955 2.985 ;
        RECT -103.965 2.815 -103.795 2.985 ;
        RECT -103.505 2.815 -103.335 2.985 ;
        RECT -103.045 2.815 -102.875 2.985 ;
        RECT -102.585 2.815 -102.415 2.985 ;
        RECT -102.125 2.815 -101.955 2.985 ;
        RECT -101.665 2.815 -101.495 2.985 ;
        RECT -101.205 2.815 -101.035 2.985 ;
        RECT -94.045 2.815 -93.875 2.985 ;
        RECT -93.585 2.815 -93.415 2.985 ;
        RECT -93.125 2.815 -92.955 2.985 ;
        RECT -92.665 2.815 -92.495 2.985 ;
        RECT -92.205 2.815 -92.035 2.985 ;
        RECT -91.745 2.815 -91.575 2.985 ;
        RECT -91.285 2.815 -91.115 2.985 ;
        RECT -84.125 2.815 -83.955 2.985 ;
        RECT -83.665 2.815 -83.495 2.985 ;
        RECT -83.205 2.815 -83.035 2.985 ;
        RECT -82.745 2.815 -82.575 2.985 ;
        RECT -82.285 2.815 -82.115 2.985 ;
        RECT -81.825 2.815 -81.655 2.985 ;
        RECT -81.365 2.815 -81.195 2.985 ;
        RECT -74.205 2.815 -74.035 2.985 ;
        RECT -73.745 2.815 -73.575 2.985 ;
        RECT -73.285 2.815 -73.115 2.985 ;
        RECT -72.825 2.815 -72.655 2.985 ;
        RECT -72.365 2.815 -72.195 2.985 ;
        RECT -71.905 2.815 -71.735 2.985 ;
        RECT -71.445 2.815 -71.275 2.985 ;
        RECT -64.285 2.815 -64.115 2.985 ;
        RECT -63.825 2.815 -63.655 2.985 ;
        RECT -63.365 2.815 -63.195 2.985 ;
        RECT -62.905 2.815 -62.735 2.985 ;
        RECT -62.445 2.815 -62.275 2.985 ;
        RECT -61.985 2.815 -61.815 2.985 ;
        RECT -61.525 2.815 -61.355 2.985 ;
        RECT -54.365 2.815 -54.195 2.985 ;
        RECT -53.905 2.815 -53.735 2.985 ;
        RECT -53.445 2.815 -53.275 2.985 ;
        RECT -52.985 2.815 -52.815 2.985 ;
        RECT -52.525 2.815 -52.355 2.985 ;
        RECT -52.065 2.815 -51.895 2.985 ;
        RECT -51.605 2.815 -51.435 2.985 ;
        RECT -44.445 2.815 -44.275 2.985 ;
        RECT -43.985 2.815 -43.815 2.985 ;
        RECT -43.525 2.815 -43.355 2.985 ;
        RECT -43.065 2.815 -42.895 2.985 ;
        RECT -42.605 2.815 -42.435 2.985 ;
        RECT -42.145 2.815 -41.975 2.985 ;
        RECT -41.685 2.815 -41.515 2.985 ;
        RECT -34.525 2.815 -34.355 2.985 ;
        RECT -34.065 2.815 -33.895 2.985 ;
        RECT -33.605 2.815 -33.435 2.985 ;
        RECT -33.145 2.815 -32.975 2.985 ;
        RECT -32.685 2.815 -32.515 2.985 ;
        RECT -32.225 2.815 -32.055 2.985 ;
        RECT -31.765 2.815 -31.595 2.985 ;
        RECT -24.605 2.815 -24.435 2.985 ;
        RECT -24.145 2.815 -23.975 2.985 ;
        RECT -23.685 2.815 -23.515 2.985 ;
        RECT -23.225 2.815 -23.055 2.985 ;
        RECT -22.765 2.815 -22.595 2.985 ;
        RECT -22.305 2.815 -22.135 2.985 ;
        RECT -21.845 2.815 -21.675 2.985 ;
        RECT -14.685 2.815 -14.515 2.985 ;
        RECT -14.225 2.815 -14.055 2.985 ;
        RECT -13.765 2.815 -13.595 2.985 ;
        RECT -13.305 2.815 -13.135 2.985 ;
        RECT -12.845 2.815 -12.675 2.985 ;
        RECT -12.385 2.815 -12.215 2.985 ;
        RECT -11.925 2.815 -11.755 2.985 ;
        RECT -4.765 2.815 -4.595 2.985 ;
        RECT -4.305 2.815 -4.135 2.985 ;
        RECT -3.845 2.815 -3.675 2.985 ;
        RECT -3.385 2.815 -3.215 2.985 ;
        RECT -2.925 2.815 -2.755 2.985 ;
        RECT -2.465 2.815 -2.295 2.985 ;
        RECT -2.005 2.815 -1.835 2.985 ;
        RECT 5.155 2.815 5.325 2.985 ;
        RECT 5.615 2.815 5.785 2.985 ;
        RECT 6.075 2.815 6.245 2.985 ;
        RECT 6.535 2.815 6.705 2.985 ;
        RECT 6.995 2.815 7.165 2.985 ;
        RECT 7.455 2.815 7.625 2.985 ;
        RECT 7.915 2.815 8.085 2.985 ;
        RECT 15.075 2.815 15.245 2.985 ;
        RECT 15.535 2.815 15.705 2.985 ;
        RECT 15.995 2.815 16.165 2.985 ;
        RECT 16.455 2.815 16.625 2.985 ;
        RECT 16.915 2.815 17.085 2.985 ;
        RECT 17.375 2.815 17.545 2.985 ;
        RECT 17.835 2.815 18.005 2.985 ;
        RECT 24.995 2.815 25.165 2.985 ;
        RECT 25.455 2.815 25.625 2.985 ;
        RECT 25.915 2.815 26.085 2.985 ;
        RECT 26.375 2.815 26.545 2.985 ;
        RECT -286.575 2.155 -286.405 2.325 ;
        RECT -286.105 2.230 -285.935 2.400 ;
        RECT -286.575 1.695 -286.405 1.865 ;
        RECT -286.575 1.235 -286.405 1.405 ;
        RECT -285.635 2.155 -285.465 2.325 ;
        RECT -276.655 2.155 -276.485 2.325 ;
        RECT -276.185 2.230 -276.015 2.400 ;
        RECT -285.635 1.695 -285.465 1.865 ;
        RECT -276.655 1.695 -276.485 1.865 ;
        RECT -285.635 1.235 -285.465 1.405 ;
        RECT -276.655 1.235 -276.485 1.405 ;
        RECT -275.715 2.155 -275.545 2.325 ;
        RECT -266.735 2.155 -266.565 2.325 ;
        RECT -266.265 2.230 -266.095 2.400 ;
        RECT -275.715 1.695 -275.545 1.865 ;
        RECT -266.735 1.695 -266.565 1.865 ;
        RECT -275.715 1.235 -275.545 1.405 ;
        RECT -266.735 1.235 -266.565 1.405 ;
        RECT -265.795 2.155 -265.625 2.325 ;
        RECT -256.815 2.155 -256.645 2.325 ;
        RECT -256.345 2.230 -256.175 2.400 ;
        RECT -265.795 1.695 -265.625 1.865 ;
        RECT -256.815 1.695 -256.645 1.865 ;
        RECT -265.795 1.235 -265.625 1.405 ;
        RECT -256.815 1.235 -256.645 1.405 ;
        RECT -255.875 2.155 -255.705 2.325 ;
        RECT -246.895 2.155 -246.725 2.325 ;
        RECT -246.425 2.230 -246.255 2.400 ;
        RECT -255.875 1.695 -255.705 1.865 ;
        RECT -246.895 1.695 -246.725 1.865 ;
        RECT -255.875 1.235 -255.705 1.405 ;
        RECT -246.895 1.235 -246.725 1.405 ;
        RECT -245.955 2.155 -245.785 2.325 ;
        RECT -236.975 2.155 -236.805 2.325 ;
        RECT -236.505 2.230 -236.335 2.400 ;
        RECT -245.955 1.695 -245.785 1.865 ;
        RECT -236.975 1.695 -236.805 1.865 ;
        RECT -245.955 1.235 -245.785 1.405 ;
        RECT -236.975 1.235 -236.805 1.405 ;
        RECT -236.035 2.155 -235.865 2.325 ;
        RECT -227.055 2.155 -226.885 2.325 ;
        RECT -226.585 2.230 -226.415 2.400 ;
        RECT -236.035 1.695 -235.865 1.865 ;
        RECT -227.055 1.695 -226.885 1.865 ;
        RECT -236.035 1.235 -235.865 1.405 ;
        RECT -227.055 1.235 -226.885 1.405 ;
        RECT -226.115 2.155 -225.945 2.325 ;
        RECT -217.135 2.155 -216.965 2.325 ;
        RECT -216.665 2.230 -216.495 2.400 ;
        RECT -226.115 1.695 -225.945 1.865 ;
        RECT -217.135 1.695 -216.965 1.865 ;
        RECT -226.115 1.235 -225.945 1.405 ;
        RECT -217.135 1.235 -216.965 1.405 ;
        RECT -216.195 2.155 -216.025 2.325 ;
        RECT -207.215 2.155 -207.045 2.325 ;
        RECT -206.745 2.230 -206.575 2.400 ;
        RECT -216.195 1.695 -216.025 1.865 ;
        RECT -207.215 1.695 -207.045 1.865 ;
        RECT -216.195 1.235 -216.025 1.405 ;
        RECT -207.215 1.235 -207.045 1.405 ;
        RECT -206.275 2.155 -206.105 2.325 ;
        RECT -197.295 2.155 -197.125 2.325 ;
        RECT -196.825 2.230 -196.655 2.400 ;
        RECT -206.275 1.695 -206.105 1.865 ;
        RECT -197.295 1.695 -197.125 1.865 ;
        RECT -206.275 1.235 -206.105 1.405 ;
        RECT -197.295 1.235 -197.125 1.405 ;
        RECT -196.355 2.155 -196.185 2.325 ;
        RECT -187.375 2.155 -187.205 2.325 ;
        RECT -186.905 2.230 -186.735 2.400 ;
        RECT -196.355 1.695 -196.185 1.865 ;
        RECT -187.375 1.695 -187.205 1.865 ;
        RECT -196.355 1.235 -196.185 1.405 ;
        RECT -187.375 1.235 -187.205 1.405 ;
        RECT -186.435 2.155 -186.265 2.325 ;
        RECT -177.455 2.155 -177.285 2.325 ;
        RECT -176.985 2.230 -176.815 2.400 ;
        RECT -186.435 1.695 -186.265 1.865 ;
        RECT -177.455 1.695 -177.285 1.865 ;
        RECT -186.435 1.235 -186.265 1.405 ;
        RECT -177.455 1.235 -177.285 1.405 ;
        RECT -176.515 2.155 -176.345 2.325 ;
        RECT -167.535 2.155 -167.365 2.325 ;
        RECT -167.065 2.230 -166.895 2.400 ;
        RECT -176.515 1.695 -176.345 1.865 ;
        RECT -167.535 1.695 -167.365 1.865 ;
        RECT -176.515 1.235 -176.345 1.405 ;
        RECT -167.535 1.235 -167.365 1.405 ;
        RECT -166.595 2.155 -166.425 2.325 ;
        RECT -157.615 2.155 -157.445 2.325 ;
        RECT -157.145 2.230 -156.975 2.400 ;
        RECT -166.595 1.695 -166.425 1.865 ;
        RECT -157.615 1.695 -157.445 1.865 ;
        RECT -166.595 1.235 -166.425 1.405 ;
        RECT -157.615 1.235 -157.445 1.405 ;
        RECT -156.675 2.155 -156.505 2.325 ;
        RECT -147.695 2.155 -147.525 2.325 ;
        RECT -147.225 2.230 -147.055 2.400 ;
        RECT -156.675 1.695 -156.505 1.865 ;
        RECT -147.695 1.695 -147.525 1.865 ;
        RECT -156.675 1.235 -156.505 1.405 ;
        RECT -147.695 1.235 -147.525 1.405 ;
        RECT -146.755 2.155 -146.585 2.325 ;
        RECT -137.775 2.155 -137.605 2.325 ;
        RECT -137.305 2.230 -137.135 2.400 ;
        RECT -146.755 1.695 -146.585 1.865 ;
        RECT -137.775 1.695 -137.605 1.865 ;
        RECT -146.755 1.235 -146.585 1.405 ;
        RECT -137.775 1.235 -137.605 1.405 ;
        RECT -136.835 2.155 -136.665 2.325 ;
        RECT -127.855 2.155 -127.685 2.325 ;
        RECT -127.385 2.230 -127.215 2.400 ;
        RECT -136.835 1.695 -136.665 1.865 ;
        RECT -127.855 1.695 -127.685 1.865 ;
        RECT -136.835 1.235 -136.665 1.405 ;
        RECT -127.855 1.235 -127.685 1.405 ;
        RECT -126.915 2.155 -126.745 2.325 ;
        RECT -117.935 2.155 -117.765 2.325 ;
        RECT -117.465 2.230 -117.295 2.400 ;
        RECT -126.915 1.695 -126.745 1.865 ;
        RECT -117.935 1.695 -117.765 1.865 ;
        RECT -126.915 1.235 -126.745 1.405 ;
        RECT -117.935 1.235 -117.765 1.405 ;
        RECT -116.995 2.155 -116.825 2.325 ;
        RECT -108.015 2.155 -107.845 2.325 ;
        RECT -107.545 2.230 -107.375 2.400 ;
        RECT -116.995 1.695 -116.825 1.865 ;
        RECT -108.015 1.695 -107.845 1.865 ;
        RECT -116.995 1.235 -116.825 1.405 ;
        RECT -108.015 1.235 -107.845 1.405 ;
        RECT -107.075 2.155 -106.905 2.325 ;
        RECT -98.095 2.155 -97.925 2.325 ;
        RECT -97.625 2.230 -97.455 2.400 ;
        RECT -107.075 1.695 -106.905 1.865 ;
        RECT -98.095 1.695 -97.925 1.865 ;
        RECT -107.075 1.235 -106.905 1.405 ;
        RECT -98.095 1.235 -97.925 1.405 ;
        RECT -97.155 2.155 -96.985 2.325 ;
        RECT -88.175 2.155 -88.005 2.325 ;
        RECT -87.705 2.230 -87.535 2.400 ;
        RECT -97.155 1.695 -96.985 1.865 ;
        RECT -88.175 1.695 -88.005 1.865 ;
        RECT -97.155 1.235 -96.985 1.405 ;
        RECT -88.175 1.235 -88.005 1.405 ;
        RECT -87.235 2.155 -87.065 2.325 ;
        RECT -78.255 2.155 -78.085 2.325 ;
        RECT -77.785 2.230 -77.615 2.400 ;
        RECT -87.235 1.695 -87.065 1.865 ;
        RECT -78.255 1.695 -78.085 1.865 ;
        RECT -87.235 1.235 -87.065 1.405 ;
        RECT -78.255 1.235 -78.085 1.405 ;
        RECT -77.315 2.155 -77.145 2.325 ;
        RECT -68.335 2.155 -68.165 2.325 ;
        RECT -67.865 2.230 -67.695 2.400 ;
        RECT -77.315 1.695 -77.145 1.865 ;
        RECT -68.335 1.695 -68.165 1.865 ;
        RECT -77.315 1.235 -77.145 1.405 ;
        RECT -68.335 1.235 -68.165 1.405 ;
        RECT -67.395 2.155 -67.225 2.325 ;
        RECT -58.415 2.155 -58.245 2.325 ;
        RECT -57.945 2.230 -57.775 2.400 ;
        RECT -67.395 1.695 -67.225 1.865 ;
        RECT -58.415 1.695 -58.245 1.865 ;
        RECT -67.395 1.235 -67.225 1.405 ;
        RECT -58.415 1.235 -58.245 1.405 ;
        RECT -57.475 2.155 -57.305 2.325 ;
        RECT -48.495 2.155 -48.325 2.325 ;
        RECT -48.025 2.230 -47.855 2.400 ;
        RECT -57.475 1.695 -57.305 1.865 ;
        RECT -48.495 1.695 -48.325 1.865 ;
        RECT -57.475 1.235 -57.305 1.405 ;
        RECT -48.495 1.235 -48.325 1.405 ;
        RECT -47.555 2.155 -47.385 2.325 ;
        RECT -38.575 2.155 -38.405 2.325 ;
        RECT -38.105 2.230 -37.935 2.400 ;
        RECT -47.555 1.695 -47.385 1.865 ;
        RECT -38.575 1.695 -38.405 1.865 ;
        RECT -47.555 1.235 -47.385 1.405 ;
        RECT -38.575 1.235 -38.405 1.405 ;
        RECT -37.635 2.155 -37.465 2.325 ;
        RECT -28.655 2.155 -28.485 2.325 ;
        RECT -28.185 2.230 -28.015 2.400 ;
        RECT -37.635 1.695 -37.465 1.865 ;
        RECT -28.655 1.695 -28.485 1.865 ;
        RECT -37.635 1.235 -37.465 1.405 ;
        RECT -28.655 1.235 -28.485 1.405 ;
        RECT -27.715 2.155 -27.545 2.325 ;
        RECT -18.735 2.155 -18.565 2.325 ;
        RECT -18.265 2.230 -18.095 2.400 ;
        RECT -27.715 1.695 -27.545 1.865 ;
        RECT -18.735 1.695 -18.565 1.865 ;
        RECT -27.715 1.235 -27.545 1.405 ;
        RECT -18.735 1.235 -18.565 1.405 ;
        RECT -17.795 2.155 -17.625 2.325 ;
        RECT -8.815 2.155 -8.645 2.325 ;
        RECT -8.345 2.230 -8.175 2.400 ;
        RECT -17.795 1.695 -17.625 1.865 ;
        RECT -8.815 1.695 -8.645 1.865 ;
        RECT -17.795 1.235 -17.625 1.405 ;
        RECT -8.815 1.235 -8.645 1.405 ;
        RECT -7.875 2.155 -7.705 2.325 ;
        RECT 1.105 2.155 1.275 2.325 ;
        RECT 1.575 2.230 1.745 2.400 ;
        RECT -7.875 1.695 -7.705 1.865 ;
        RECT 1.105 1.695 1.275 1.865 ;
        RECT -7.875 1.235 -7.705 1.405 ;
        RECT 1.105 1.235 1.275 1.405 ;
        RECT 2.045 2.155 2.215 2.325 ;
        RECT 11.025 2.155 11.195 2.325 ;
        RECT 11.495 2.230 11.665 2.400 ;
        RECT 2.045 1.695 2.215 1.865 ;
        RECT 11.025 1.695 11.195 1.865 ;
        RECT 2.045 1.235 2.215 1.405 ;
        RECT 11.025 1.235 11.195 1.405 ;
        RECT 11.965 2.155 12.135 2.325 ;
        RECT 20.945 2.155 21.115 2.325 ;
        RECT 21.415 2.230 21.585 2.400 ;
        RECT 11.965 1.695 12.135 1.865 ;
        RECT 20.945 1.695 21.115 1.865 ;
        RECT 11.965 1.235 12.135 1.405 ;
        RECT 20.945 1.235 21.115 1.405 ;
        RECT 21.885 2.155 22.055 2.325 ;
        RECT 21.885 1.695 22.055 1.865 ;
        RECT 21.885 1.235 22.055 1.405 ;
        RECT -279.855 -86.235 -279.685 -86.065 ;
        RECT -279.385 -86.240 -279.215 -86.070 ;
        RECT -278.915 -86.235 -278.745 -86.065 ;
        RECT -279.855 -86.695 -279.685 -86.525 ;
        RECT -279.855 -87.155 -279.685 -86.985 ;
        RECT -269.935 -86.235 -269.765 -86.065 ;
        RECT -269.465 -86.240 -269.295 -86.070 ;
        RECT -268.995 -86.235 -268.825 -86.065 ;
        RECT -278.915 -86.695 -278.745 -86.525 ;
        RECT -269.935 -86.695 -269.765 -86.525 ;
        RECT -278.915 -87.155 -278.745 -86.985 ;
        RECT -269.935 -87.155 -269.765 -86.985 ;
        RECT -260.015 -86.235 -259.845 -86.065 ;
        RECT -259.545 -86.240 -259.375 -86.070 ;
        RECT -259.075 -86.235 -258.905 -86.065 ;
        RECT -268.995 -86.695 -268.825 -86.525 ;
        RECT -260.015 -86.695 -259.845 -86.525 ;
        RECT -268.995 -87.155 -268.825 -86.985 ;
        RECT -260.015 -87.155 -259.845 -86.985 ;
        RECT -250.095 -86.235 -249.925 -86.065 ;
        RECT -249.625 -86.240 -249.455 -86.070 ;
        RECT -249.155 -86.235 -248.985 -86.065 ;
        RECT -259.075 -86.695 -258.905 -86.525 ;
        RECT -250.095 -86.695 -249.925 -86.525 ;
        RECT -259.075 -87.155 -258.905 -86.985 ;
        RECT -250.095 -87.155 -249.925 -86.985 ;
        RECT -240.175 -86.235 -240.005 -86.065 ;
        RECT -239.705 -86.240 -239.535 -86.070 ;
        RECT -239.235 -86.235 -239.065 -86.065 ;
        RECT -249.155 -86.695 -248.985 -86.525 ;
        RECT -240.175 -86.695 -240.005 -86.525 ;
        RECT -249.155 -87.155 -248.985 -86.985 ;
        RECT -240.175 -87.155 -240.005 -86.985 ;
        RECT -230.255 -86.235 -230.085 -86.065 ;
        RECT -229.785 -86.240 -229.615 -86.070 ;
        RECT -229.315 -86.235 -229.145 -86.065 ;
        RECT -239.235 -86.695 -239.065 -86.525 ;
        RECT -230.255 -86.695 -230.085 -86.525 ;
        RECT -239.235 -87.155 -239.065 -86.985 ;
        RECT -230.255 -87.155 -230.085 -86.985 ;
        RECT -220.335 -86.235 -220.165 -86.065 ;
        RECT -219.865 -86.240 -219.695 -86.070 ;
        RECT -219.395 -86.235 -219.225 -86.065 ;
        RECT -229.315 -86.695 -229.145 -86.525 ;
        RECT -220.335 -86.695 -220.165 -86.525 ;
        RECT -229.315 -87.155 -229.145 -86.985 ;
        RECT -220.335 -87.155 -220.165 -86.985 ;
        RECT -210.415 -86.235 -210.245 -86.065 ;
        RECT -209.945 -86.240 -209.775 -86.070 ;
        RECT -209.475 -86.235 -209.305 -86.065 ;
        RECT -219.395 -86.695 -219.225 -86.525 ;
        RECT -210.415 -86.695 -210.245 -86.525 ;
        RECT -219.395 -87.155 -219.225 -86.985 ;
        RECT -210.415 -87.155 -210.245 -86.985 ;
        RECT -200.495 -86.235 -200.325 -86.065 ;
        RECT -200.025 -86.240 -199.855 -86.070 ;
        RECT -199.555 -86.235 -199.385 -86.065 ;
        RECT -209.475 -86.695 -209.305 -86.525 ;
        RECT -200.495 -86.695 -200.325 -86.525 ;
        RECT -209.475 -87.155 -209.305 -86.985 ;
        RECT -200.495 -87.155 -200.325 -86.985 ;
        RECT -190.575 -86.235 -190.405 -86.065 ;
        RECT -190.105 -86.240 -189.935 -86.070 ;
        RECT -189.635 -86.235 -189.465 -86.065 ;
        RECT -199.555 -86.695 -199.385 -86.525 ;
        RECT -190.575 -86.695 -190.405 -86.525 ;
        RECT -199.555 -87.155 -199.385 -86.985 ;
        RECT -190.575 -87.155 -190.405 -86.985 ;
        RECT -180.655 -86.235 -180.485 -86.065 ;
        RECT -180.185 -86.240 -180.015 -86.070 ;
        RECT -179.715 -86.235 -179.545 -86.065 ;
        RECT -189.635 -86.695 -189.465 -86.525 ;
        RECT -180.655 -86.695 -180.485 -86.525 ;
        RECT -189.635 -87.155 -189.465 -86.985 ;
        RECT -180.655 -87.155 -180.485 -86.985 ;
        RECT -170.735 -86.235 -170.565 -86.065 ;
        RECT -170.265 -86.240 -170.095 -86.070 ;
        RECT -169.795 -86.235 -169.625 -86.065 ;
        RECT -179.715 -86.695 -179.545 -86.525 ;
        RECT -170.735 -86.695 -170.565 -86.525 ;
        RECT -179.715 -87.155 -179.545 -86.985 ;
        RECT -170.735 -87.155 -170.565 -86.985 ;
        RECT -160.815 -86.235 -160.645 -86.065 ;
        RECT -160.345 -86.240 -160.175 -86.070 ;
        RECT -159.875 -86.235 -159.705 -86.065 ;
        RECT -169.795 -86.695 -169.625 -86.525 ;
        RECT -160.815 -86.695 -160.645 -86.525 ;
        RECT -169.795 -87.155 -169.625 -86.985 ;
        RECT -160.815 -87.155 -160.645 -86.985 ;
        RECT -150.895 -86.235 -150.725 -86.065 ;
        RECT -150.425 -86.240 -150.255 -86.070 ;
        RECT -149.955 -86.235 -149.785 -86.065 ;
        RECT -159.875 -86.695 -159.705 -86.525 ;
        RECT -150.895 -86.695 -150.725 -86.525 ;
        RECT -159.875 -87.155 -159.705 -86.985 ;
        RECT -150.895 -87.155 -150.725 -86.985 ;
        RECT -140.975 -86.235 -140.805 -86.065 ;
        RECT -140.505 -86.240 -140.335 -86.070 ;
        RECT -140.035 -86.235 -139.865 -86.065 ;
        RECT -149.955 -86.695 -149.785 -86.525 ;
        RECT -140.975 -86.695 -140.805 -86.525 ;
        RECT -149.955 -87.155 -149.785 -86.985 ;
        RECT -140.975 -87.155 -140.805 -86.985 ;
        RECT -131.055 -86.235 -130.885 -86.065 ;
        RECT -130.585 -86.240 -130.415 -86.070 ;
        RECT -130.115 -86.235 -129.945 -86.065 ;
        RECT -140.035 -86.695 -139.865 -86.525 ;
        RECT -131.055 -86.695 -130.885 -86.525 ;
        RECT -140.035 -87.155 -139.865 -86.985 ;
        RECT -131.055 -87.155 -130.885 -86.985 ;
        RECT -121.135 -86.235 -120.965 -86.065 ;
        RECT -120.665 -86.240 -120.495 -86.070 ;
        RECT -120.195 -86.235 -120.025 -86.065 ;
        RECT -130.115 -86.695 -129.945 -86.525 ;
        RECT -121.135 -86.695 -120.965 -86.525 ;
        RECT -130.115 -87.155 -129.945 -86.985 ;
        RECT -121.135 -87.155 -120.965 -86.985 ;
        RECT -111.215 -86.235 -111.045 -86.065 ;
        RECT -110.745 -86.240 -110.575 -86.070 ;
        RECT -110.275 -86.235 -110.105 -86.065 ;
        RECT -120.195 -86.695 -120.025 -86.525 ;
        RECT -111.215 -86.695 -111.045 -86.525 ;
        RECT -120.195 -87.155 -120.025 -86.985 ;
        RECT -111.215 -87.155 -111.045 -86.985 ;
        RECT -101.295 -86.235 -101.125 -86.065 ;
        RECT -100.825 -86.240 -100.655 -86.070 ;
        RECT -100.355 -86.235 -100.185 -86.065 ;
        RECT -110.275 -86.695 -110.105 -86.525 ;
        RECT -101.295 -86.695 -101.125 -86.525 ;
        RECT -110.275 -87.155 -110.105 -86.985 ;
        RECT -101.295 -87.155 -101.125 -86.985 ;
        RECT -91.375 -86.235 -91.205 -86.065 ;
        RECT -90.905 -86.240 -90.735 -86.070 ;
        RECT -90.435 -86.235 -90.265 -86.065 ;
        RECT -100.355 -86.695 -100.185 -86.525 ;
        RECT -91.375 -86.695 -91.205 -86.525 ;
        RECT -100.355 -87.155 -100.185 -86.985 ;
        RECT -91.375 -87.155 -91.205 -86.985 ;
        RECT -81.455 -86.235 -81.285 -86.065 ;
        RECT -80.985 -86.240 -80.815 -86.070 ;
        RECT -80.515 -86.235 -80.345 -86.065 ;
        RECT -90.435 -86.695 -90.265 -86.525 ;
        RECT -81.455 -86.695 -81.285 -86.525 ;
        RECT -90.435 -87.155 -90.265 -86.985 ;
        RECT -81.455 -87.155 -81.285 -86.985 ;
        RECT -71.535 -86.235 -71.365 -86.065 ;
        RECT -71.065 -86.240 -70.895 -86.070 ;
        RECT -70.595 -86.235 -70.425 -86.065 ;
        RECT -80.515 -86.695 -80.345 -86.525 ;
        RECT -71.535 -86.695 -71.365 -86.525 ;
        RECT -80.515 -87.155 -80.345 -86.985 ;
        RECT -71.535 -87.155 -71.365 -86.985 ;
        RECT -61.615 -86.235 -61.445 -86.065 ;
        RECT -61.145 -86.240 -60.975 -86.070 ;
        RECT -60.675 -86.235 -60.505 -86.065 ;
        RECT -70.595 -86.695 -70.425 -86.525 ;
        RECT -61.615 -86.695 -61.445 -86.525 ;
        RECT -70.595 -87.155 -70.425 -86.985 ;
        RECT -61.615 -87.155 -61.445 -86.985 ;
        RECT -51.695 -86.235 -51.525 -86.065 ;
        RECT -51.225 -86.240 -51.055 -86.070 ;
        RECT -50.755 -86.235 -50.585 -86.065 ;
        RECT -60.675 -86.695 -60.505 -86.525 ;
        RECT -51.695 -86.695 -51.525 -86.525 ;
        RECT -60.675 -87.155 -60.505 -86.985 ;
        RECT -51.695 -87.155 -51.525 -86.985 ;
        RECT -41.775 -86.235 -41.605 -86.065 ;
        RECT -41.305 -86.240 -41.135 -86.070 ;
        RECT -40.835 -86.235 -40.665 -86.065 ;
        RECT -50.755 -86.695 -50.585 -86.525 ;
        RECT -41.775 -86.695 -41.605 -86.525 ;
        RECT -50.755 -87.155 -50.585 -86.985 ;
        RECT -41.775 -87.155 -41.605 -86.985 ;
        RECT -31.855 -86.235 -31.685 -86.065 ;
        RECT -31.385 -86.240 -31.215 -86.070 ;
        RECT -30.915 -86.235 -30.745 -86.065 ;
        RECT -40.835 -86.695 -40.665 -86.525 ;
        RECT -31.855 -86.695 -31.685 -86.525 ;
        RECT -40.835 -87.155 -40.665 -86.985 ;
        RECT -31.855 -87.155 -31.685 -86.985 ;
        RECT -21.935 -86.235 -21.765 -86.065 ;
        RECT -21.465 -86.240 -21.295 -86.070 ;
        RECT -20.995 -86.235 -20.825 -86.065 ;
        RECT -30.915 -86.695 -30.745 -86.525 ;
        RECT -21.935 -86.695 -21.765 -86.525 ;
        RECT -30.915 -87.155 -30.745 -86.985 ;
        RECT -21.935 -87.155 -21.765 -86.985 ;
        RECT -12.015 -86.235 -11.845 -86.065 ;
        RECT -11.545 -86.240 -11.375 -86.070 ;
        RECT -11.075 -86.235 -10.905 -86.065 ;
        RECT -20.995 -86.695 -20.825 -86.525 ;
        RECT -12.015 -86.695 -11.845 -86.525 ;
        RECT -20.995 -87.155 -20.825 -86.985 ;
        RECT -12.015 -87.155 -11.845 -86.985 ;
        RECT -2.095 -86.235 -1.925 -86.065 ;
        RECT -1.625 -86.240 -1.455 -86.070 ;
        RECT -1.155 -86.235 -0.985 -86.065 ;
        RECT -11.075 -86.695 -10.905 -86.525 ;
        RECT -2.095 -86.695 -1.925 -86.525 ;
        RECT -11.075 -87.155 -10.905 -86.985 ;
        RECT -2.095 -87.155 -1.925 -86.985 ;
        RECT 7.825 -86.235 7.995 -86.065 ;
        RECT 8.295 -86.240 8.465 -86.070 ;
        RECT 8.765 -86.235 8.935 -86.065 ;
        RECT -1.155 -86.695 -0.985 -86.525 ;
        RECT 7.825 -86.695 7.995 -86.525 ;
        RECT -1.155 -87.155 -0.985 -86.985 ;
        RECT 7.825 -87.155 7.995 -86.985 ;
        RECT 17.745 -86.235 17.915 -86.065 ;
        RECT 18.215 -86.240 18.385 -86.070 ;
        RECT 18.685 -86.235 18.855 -86.065 ;
        RECT 8.765 -86.695 8.935 -86.525 ;
        RECT 17.745 -86.695 17.915 -86.525 ;
        RECT 8.765 -87.155 8.935 -86.985 ;
        RECT 17.745 -87.155 17.915 -86.985 ;
        RECT 27.665 -86.235 27.835 -86.065 ;
        RECT 28.135 -86.240 28.305 -86.070 ;
        RECT 18.685 -86.695 18.855 -86.525 ;
        RECT 27.665 -86.695 27.835 -86.525 ;
        RECT 18.685 -87.155 18.855 -86.985 ;
        RECT 27.665 -87.155 27.835 -86.985 ;
        RECT -285.725 -87.815 -285.555 -87.645 ;
        RECT -285.265 -87.815 -285.095 -87.645 ;
        RECT -284.805 -87.815 -284.635 -87.645 ;
        RECT -284.345 -87.815 -284.175 -87.645 ;
        RECT -283.885 -87.815 -283.715 -87.645 ;
        RECT -283.425 -87.815 -283.255 -87.645 ;
        RECT -282.965 -87.815 -282.795 -87.645 ;
        RECT -275.805 -87.815 -275.635 -87.645 ;
        RECT -275.345 -87.815 -275.175 -87.645 ;
        RECT -274.885 -87.815 -274.715 -87.645 ;
        RECT -274.425 -87.815 -274.255 -87.645 ;
        RECT -273.965 -87.815 -273.795 -87.645 ;
        RECT -273.505 -87.815 -273.335 -87.645 ;
        RECT -273.045 -87.815 -272.875 -87.645 ;
        RECT -265.885 -87.815 -265.715 -87.645 ;
        RECT -265.425 -87.815 -265.255 -87.645 ;
        RECT -264.965 -87.815 -264.795 -87.645 ;
        RECT -264.505 -87.815 -264.335 -87.645 ;
        RECT -264.045 -87.815 -263.875 -87.645 ;
        RECT -263.585 -87.815 -263.415 -87.645 ;
        RECT -263.125 -87.815 -262.955 -87.645 ;
        RECT -255.965 -87.815 -255.795 -87.645 ;
        RECT -255.505 -87.815 -255.335 -87.645 ;
        RECT -255.045 -87.815 -254.875 -87.645 ;
        RECT -254.585 -87.815 -254.415 -87.645 ;
        RECT -254.125 -87.815 -253.955 -87.645 ;
        RECT -253.665 -87.815 -253.495 -87.645 ;
        RECT -253.205 -87.815 -253.035 -87.645 ;
        RECT -246.045 -87.815 -245.875 -87.645 ;
        RECT -245.585 -87.815 -245.415 -87.645 ;
        RECT -245.125 -87.815 -244.955 -87.645 ;
        RECT -244.665 -87.815 -244.495 -87.645 ;
        RECT -244.205 -87.815 -244.035 -87.645 ;
        RECT -243.745 -87.815 -243.575 -87.645 ;
        RECT -243.285 -87.815 -243.115 -87.645 ;
        RECT -236.125 -87.815 -235.955 -87.645 ;
        RECT -235.665 -87.815 -235.495 -87.645 ;
        RECT -235.205 -87.815 -235.035 -87.645 ;
        RECT -234.745 -87.815 -234.575 -87.645 ;
        RECT -234.285 -87.815 -234.115 -87.645 ;
        RECT -233.825 -87.815 -233.655 -87.645 ;
        RECT -233.365 -87.815 -233.195 -87.645 ;
        RECT -226.205 -87.815 -226.035 -87.645 ;
        RECT -225.745 -87.815 -225.575 -87.645 ;
        RECT -225.285 -87.815 -225.115 -87.645 ;
        RECT -224.825 -87.815 -224.655 -87.645 ;
        RECT -224.365 -87.815 -224.195 -87.645 ;
        RECT -223.905 -87.815 -223.735 -87.645 ;
        RECT -223.445 -87.815 -223.275 -87.645 ;
        RECT -216.285 -87.815 -216.115 -87.645 ;
        RECT -215.825 -87.815 -215.655 -87.645 ;
        RECT -215.365 -87.815 -215.195 -87.645 ;
        RECT -214.905 -87.815 -214.735 -87.645 ;
        RECT -214.445 -87.815 -214.275 -87.645 ;
        RECT -213.985 -87.815 -213.815 -87.645 ;
        RECT -213.525 -87.815 -213.355 -87.645 ;
        RECT -206.365 -87.815 -206.195 -87.645 ;
        RECT -205.905 -87.815 -205.735 -87.645 ;
        RECT -205.445 -87.815 -205.275 -87.645 ;
        RECT -204.985 -87.815 -204.815 -87.645 ;
        RECT -204.525 -87.815 -204.355 -87.645 ;
        RECT -204.065 -87.815 -203.895 -87.645 ;
        RECT -203.605 -87.815 -203.435 -87.645 ;
        RECT -196.445 -87.815 -196.275 -87.645 ;
        RECT -195.985 -87.815 -195.815 -87.645 ;
        RECT -195.525 -87.815 -195.355 -87.645 ;
        RECT -195.065 -87.815 -194.895 -87.645 ;
        RECT -194.605 -87.815 -194.435 -87.645 ;
        RECT -194.145 -87.815 -193.975 -87.645 ;
        RECT -193.685 -87.815 -193.515 -87.645 ;
        RECT -186.525 -87.815 -186.355 -87.645 ;
        RECT -186.065 -87.815 -185.895 -87.645 ;
        RECT -185.605 -87.815 -185.435 -87.645 ;
        RECT -185.145 -87.815 -184.975 -87.645 ;
        RECT -184.685 -87.815 -184.515 -87.645 ;
        RECT -184.225 -87.815 -184.055 -87.645 ;
        RECT -183.765 -87.815 -183.595 -87.645 ;
        RECT -176.605 -87.815 -176.435 -87.645 ;
        RECT -176.145 -87.815 -175.975 -87.645 ;
        RECT -175.685 -87.815 -175.515 -87.645 ;
        RECT -175.225 -87.815 -175.055 -87.645 ;
        RECT -174.765 -87.815 -174.595 -87.645 ;
        RECT -174.305 -87.815 -174.135 -87.645 ;
        RECT -173.845 -87.815 -173.675 -87.645 ;
        RECT -166.685 -87.815 -166.515 -87.645 ;
        RECT -166.225 -87.815 -166.055 -87.645 ;
        RECT -165.765 -87.815 -165.595 -87.645 ;
        RECT -165.305 -87.815 -165.135 -87.645 ;
        RECT -164.845 -87.815 -164.675 -87.645 ;
        RECT -164.385 -87.815 -164.215 -87.645 ;
        RECT -163.925 -87.815 -163.755 -87.645 ;
        RECT -156.765 -87.815 -156.595 -87.645 ;
        RECT -156.305 -87.815 -156.135 -87.645 ;
        RECT -155.845 -87.815 -155.675 -87.645 ;
        RECT -155.385 -87.815 -155.215 -87.645 ;
        RECT -154.925 -87.815 -154.755 -87.645 ;
        RECT -154.465 -87.815 -154.295 -87.645 ;
        RECT -154.005 -87.815 -153.835 -87.645 ;
        RECT -146.845 -87.815 -146.675 -87.645 ;
        RECT -146.385 -87.815 -146.215 -87.645 ;
        RECT -145.925 -87.815 -145.755 -87.645 ;
        RECT -145.465 -87.815 -145.295 -87.645 ;
        RECT -145.005 -87.815 -144.835 -87.645 ;
        RECT -144.545 -87.815 -144.375 -87.645 ;
        RECT -144.085 -87.815 -143.915 -87.645 ;
        RECT -136.925 -87.815 -136.755 -87.645 ;
        RECT -136.465 -87.815 -136.295 -87.645 ;
        RECT -136.005 -87.815 -135.835 -87.645 ;
        RECT -135.545 -87.815 -135.375 -87.645 ;
        RECT -135.085 -87.815 -134.915 -87.645 ;
        RECT -134.625 -87.815 -134.455 -87.645 ;
        RECT -134.165 -87.815 -133.995 -87.645 ;
        RECT -127.005 -87.815 -126.835 -87.645 ;
        RECT -126.545 -87.815 -126.375 -87.645 ;
        RECT -126.085 -87.815 -125.915 -87.645 ;
        RECT -125.625 -87.815 -125.455 -87.645 ;
        RECT -125.165 -87.815 -124.995 -87.645 ;
        RECT -124.705 -87.815 -124.535 -87.645 ;
        RECT -124.245 -87.815 -124.075 -87.645 ;
        RECT -117.085 -87.815 -116.915 -87.645 ;
        RECT -116.625 -87.815 -116.455 -87.645 ;
        RECT -116.165 -87.815 -115.995 -87.645 ;
        RECT -115.705 -87.815 -115.535 -87.645 ;
        RECT -115.245 -87.815 -115.075 -87.645 ;
        RECT -114.785 -87.815 -114.615 -87.645 ;
        RECT -114.325 -87.815 -114.155 -87.645 ;
        RECT -107.165 -87.815 -106.995 -87.645 ;
        RECT -106.705 -87.815 -106.535 -87.645 ;
        RECT -106.245 -87.815 -106.075 -87.645 ;
        RECT -105.785 -87.815 -105.615 -87.645 ;
        RECT -105.325 -87.815 -105.155 -87.645 ;
        RECT -104.865 -87.815 -104.695 -87.645 ;
        RECT -104.405 -87.815 -104.235 -87.645 ;
        RECT -97.245 -87.815 -97.075 -87.645 ;
        RECT -96.785 -87.815 -96.615 -87.645 ;
        RECT -96.325 -87.815 -96.155 -87.645 ;
        RECT -95.865 -87.815 -95.695 -87.645 ;
        RECT -95.405 -87.815 -95.235 -87.645 ;
        RECT -94.945 -87.815 -94.775 -87.645 ;
        RECT -94.485 -87.815 -94.315 -87.645 ;
        RECT -87.325 -87.815 -87.155 -87.645 ;
        RECT -86.865 -87.815 -86.695 -87.645 ;
        RECT -86.405 -87.815 -86.235 -87.645 ;
        RECT -85.945 -87.815 -85.775 -87.645 ;
        RECT -85.485 -87.815 -85.315 -87.645 ;
        RECT -85.025 -87.815 -84.855 -87.645 ;
        RECT -84.565 -87.815 -84.395 -87.645 ;
        RECT -77.405 -87.815 -77.235 -87.645 ;
        RECT -76.945 -87.815 -76.775 -87.645 ;
        RECT -76.485 -87.815 -76.315 -87.645 ;
        RECT -76.025 -87.815 -75.855 -87.645 ;
        RECT -75.565 -87.815 -75.395 -87.645 ;
        RECT -75.105 -87.815 -74.935 -87.645 ;
        RECT -74.645 -87.815 -74.475 -87.645 ;
        RECT -67.485 -87.815 -67.315 -87.645 ;
        RECT -67.025 -87.815 -66.855 -87.645 ;
        RECT -66.565 -87.815 -66.395 -87.645 ;
        RECT -66.105 -87.815 -65.935 -87.645 ;
        RECT -65.645 -87.815 -65.475 -87.645 ;
        RECT -65.185 -87.815 -65.015 -87.645 ;
        RECT -64.725 -87.815 -64.555 -87.645 ;
        RECT -57.565 -87.815 -57.395 -87.645 ;
        RECT -57.105 -87.815 -56.935 -87.645 ;
        RECT -56.645 -87.815 -56.475 -87.645 ;
        RECT -56.185 -87.815 -56.015 -87.645 ;
        RECT -55.725 -87.815 -55.555 -87.645 ;
        RECT -55.265 -87.815 -55.095 -87.645 ;
        RECT -54.805 -87.815 -54.635 -87.645 ;
        RECT -47.645 -87.815 -47.475 -87.645 ;
        RECT -47.185 -87.815 -47.015 -87.645 ;
        RECT -46.725 -87.815 -46.555 -87.645 ;
        RECT -46.265 -87.815 -46.095 -87.645 ;
        RECT -45.805 -87.815 -45.635 -87.645 ;
        RECT -45.345 -87.815 -45.175 -87.645 ;
        RECT -44.885 -87.815 -44.715 -87.645 ;
        RECT -37.725 -87.815 -37.555 -87.645 ;
        RECT -37.265 -87.815 -37.095 -87.645 ;
        RECT -36.805 -87.815 -36.635 -87.645 ;
        RECT -36.345 -87.815 -36.175 -87.645 ;
        RECT -35.885 -87.815 -35.715 -87.645 ;
        RECT -35.425 -87.815 -35.255 -87.645 ;
        RECT -34.965 -87.815 -34.795 -87.645 ;
        RECT -27.805 -87.815 -27.635 -87.645 ;
        RECT -27.345 -87.815 -27.175 -87.645 ;
        RECT -26.885 -87.815 -26.715 -87.645 ;
        RECT -26.425 -87.815 -26.255 -87.645 ;
        RECT -25.965 -87.815 -25.795 -87.645 ;
        RECT -25.505 -87.815 -25.335 -87.645 ;
        RECT -25.045 -87.815 -24.875 -87.645 ;
        RECT -17.885 -87.815 -17.715 -87.645 ;
        RECT -17.425 -87.815 -17.255 -87.645 ;
        RECT -16.965 -87.815 -16.795 -87.645 ;
        RECT -16.505 -87.815 -16.335 -87.645 ;
        RECT -16.045 -87.815 -15.875 -87.645 ;
        RECT -15.585 -87.815 -15.415 -87.645 ;
        RECT -15.125 -87.815 -14.955 -87.645 ;
        RECT -7.965 -87.815 -7.795 -87.645 ;
        RECT -7.505 -87.815 -7.335 -87.645 ;
        RECT -7.045 -87.815 -6.875 -87.645 ;
        RECT -6.585 -87.815 -6.415 -87.645 ;
        RECT -6.125 -87.815 -5.955 -87.645 ;
        RECT -5.665 -87.815 -5.495 -87.645 ;
        RECT -5.205 -87.815 -5.035 -87.645 ;
        RECT 1.955 -87.815 2.125 -87.645 ;
        RECT 2.415 -87.815 2.585 -87.645 ;
        RECT 2.875 -87.815 3.045 -87.645 ;
        RECT 3.335 -87.815 3.505 -87.645 ;
        RECT 3.795 -87.815 3.965 -87.645 ;
        RECT 4.255 -87.815 4.425 -87.645 ;
        RECT 4.715 -87.815 4.885 -87.645 ;
        RECT 11.875 -87.815 12.045 -87.645 ;
        RECT 12.335 -87.815 12.505 -87.645 ;
        RECT 12.795 -87.815 12.965 -87.645 ;
        RECT 13.255 -87.815 13.425 -87.645 ;
        RECT 13.715 -87.815 13.885 -87.645 ;
        RECT 14.175 -87.815 14.345 -87.645 ;
        RECT 14.635 -87.815 14.805 -87.645 ;
        RECT 21.795 -87.815 21.965 -87.645 ;
        RECT 22.255 -87.815 22.425 -87.645 ;
        RECT 22.715 -87.815 22.885 -87.645 ;
        RECT 23.175 -87.815 23.345 -87.645 ;
        RECT 23.635 -87.815 23.805 -87.645 ;
        RECT 24.095 -87.815 24.265 -87.645 ;
        RECT 24.555 -87.815 24.725 -87.645 ;
        RECT -280.765 -90.535 -280.595 -90.365 ;
        RECT -280.305 -90.535 -280.135 -90.365 ;
        RECT -279.845 -90.535 -279.675 -90.365 ;
        RECT -279.385 -90.535 -279.215 -90.365 ;
        RECT -278.925 -90.535 -278.755 -90.365 ;
        RECT -278.465 -90.535 -278.295 -90.365 ;
        RECT -278.005 -90.535 -277.835 -90.365 ;
        RECT -270.845 -90.535 -270.675 -90.365 ;
        RECT -270.385 -90.535 -270.215 -90.365 ;
        RECT -269.925 -90.535 -269.755 -90.365 ;
        RECT -269.465 -90.535 -269.295 -90.365 ;
        RECT -269.005 -90.535 -268.835 -90.365 ;
        RECT -268.545 -90.535 -268.375 -90.365 ;
        RECT -268.085 -90.535 -267.915 -90.365 ;
        RECT -260.925 -90.535 -260.755 -90.365 ;
        RECT -260.465 -90.535 -260.295 -90.365 ;
        RECT -260.005 -90.535 -259.835 -90.365 ;
        RECT -259.545 -90.535 -259.375 -90.365 ;
        RECT -259.085 -90.535 -258.915 -90.365 ;
        RECT -258.625 -90.535 -258.455 -90.365 ;
        RECT -258.165 -90.535 -257.995 -90.365 ;
        RECT -251.005 -90.535 -250.835 -90.365 ;
        RECT -250.545 -90.535 -250.375 -90.365 ;
        RECT -250.085 -90.535 -249.915 -90.365 ;
        RECT -249.625 -90.535 -249.455 -90.365 ;
        RECT -249.165 -90.535 -248.995 -90.365 ;
        RECT -248.705 -90.535 -248.535 -90.365 ;
        RECT -248.245 -90.535 -248.075 -90.365 ;
        RECT -241.085 -90.535 -240.915 -90.365 ;
        RECT -240.625 -90.535 -240.455 -90.365 ;
        RECT -240.165 -90.535 -239.995 -90.365 ;
        RECT -239.705 -90.535 -239.535 -90.365 ;
        RECT -239.245 -90.535 -239.075 -90.365 ;
        RECT -238.785 -90.535 -238.615 -90.365 ;
        RECT -238.325 -90.535 -238.155 -90.365 ;
        RECT -231.165 -90.535 -230.995 -90.365 ;
        RECT -230.705 -90.535 -230.535 -90.365 ;
        RECT -230.245 -90.535 -230.075 -90.365 ;
        RECT -229.785 -90.535 -229.615 -90.365 ;
        RECT -229.325 -90.535 -229.155 -90.365 ;
        RECT -228.865 -90.535 -228.695 -90.365 ;
        RECT -228.405 -90.535 -228.235 -90.365 ;
        RECT -221.245 -90.535 -221.075 -90.365 ;
        RECT -220.785 -90.535 -220.615 -90.365 ;
        RECT -220.325 -90.535 -220.155 -90.365 ;
        RECT -219.865 -90.535 -219.695 -90.365 ;
        RECT -219.405 -90.535 -219.235 -90.365 ;
        RECT -218.945 -90.535 -218.775 -90.365 ;
        RECT -218.485 -90.535 -218.315 -90.365 ;
        RECT -211.325 -90.535 -211.155 -90.365 ;
        RECT -210.865 -90.535 -210.695 -90.365 ;
        RECT -210.405 -90.535 -210.235 -90.365 ;
        RECT -209.945 -90.535 -209.775 -90.365 ;
        RECT -209.485 -90.535 -209.315 -90.365 ;
        RECT -209.025 -90.535 -208.855 -90.365 ;
        RECT -208.565 -90.535 -208.395 -90.365 ;
        RECT -201.405 -90.535 -201.235 -90.365 ;
        RECT -200.945 -90.535 -200.775 -90.365 ;
        RECT -200.485 -90.535 -200.315 -90.365 ;
        RECT -200.025 -90.535 -199.855 -90.365 ;
        RECT -199.565 -90.535 -199.395 -90.365 ;
        RECT -199.105 -90.535 -198.935 -90.365 ;
        RECT -198.645 -90.535 -198.475 -90.365 ;
        RECT -191.485 -90.535 -191.315 -90.365 ;
        RECT -191.025 -90.535 -190.855 -90.365 ;
        RECT -190.565 -90.535 -190.395 -90.365 ;
        RECT -190.105 -90.535 -189.935 -90.365 ;
        RECT -189.645 -90.535 -189.475 -90.365 ;
        RECT -189.185 -90.535 -189.015 -90.365 ;
        RECT -188.725 -90.535 -188.555 -90.365 ;
        RECT -181.565 -90.535 -181.395 -90.365 ;
        RECT -181.105 -90.535 -180.935 -90.365 ;
        RECT -180.645 -90.535 -180.475 -90.365 ;
        RECT -180.185 -90.535 -180.015 -90.365 ;
        RECT -179.725 -90.535 -179.555 -90.365 ;
        RECT -179.265 -90.535 -179.095 -90.365 ;
        RECT -178.805 -90.535 -178.635 -90.365 ;
        RECT -171.645 -90.535 -171.475 -90.365 ;
        RECT -171.185 -90.535 -171.015 -90.365 ;
        RECT -170.725 -90.535 -170.555 -90.365 ;
        RECT -170.265 -90.535 -170.095 -90.365 ;
        RECT -169.805 -90.535 -169.635 -90.365 ;
        RECT -169.345 -90.535 -169.175 -90.365 ;
        RECT -168.885 -90.535 -168.715 -90.365 ;
        RECT -161.725 -90.535 -161.555 -90.365 ;
        RECT -161.265 -90.535 -161.095 -90.365 ;
        RECT -160.805 -90.535 -160.635 -90.365 ;
        RECT -160.345 -90.535 -160.175 -90.365 ;
        RECT -159.885 -90.535 -159.715 -90.365 ;
        RECT -159.425 -90.535 -159.255 -90.365 ;
        RECT -158.965 -90.535 -158.795 -90.365 ;
        RECT -151.805 -90.535 -151.635 -90.365 ;
        RECT -151.345 -90.535 -151.175 -90.365 ;
        RECT -150.885 -90.535 -150.715 -90.365 ;
        RECT -150.425 -90.535 -150.255 -90.365 ;
        RECT -149.965 -90.535 -149.795 -90.365 ;
        RECT -149.505 -90.535 -149.335 -90.365 ;
        RECT -149.045 -90.535 -148.875 -90.365 ;
        RECT -141.885 -90.535 -141.715 -90.365 ;
        RECT -141.425 -90.535 -141.255 -90.365 ;
        RECT -140.965 -90.535 -140.795 -90.365 ;
        RECT -140.505 -90.535 -140.335 -90.365 ;
        RECT -140.045 -90.535 -139.875 -90.365 ;
        RECT -139.585 -90.535 -139.415 -90.365 ;
        RECT -139.125 -90.535 -138.955 -90.365 ;
        RECT -131.965 -90.535 -131.795 -90.365 ;
        RECT -131.505 -90.535 -131.335 -90.365 ;
        RECT -131.045 -90.535 -130.875 -90.365 ;
        RECT -130.585 -90.535 -130.415 -90.365 ;
        RECT -130.125 -90.535 -129.955 -90.365 ;
        RECT -129.665 -90.535 -129.495 -90.365 ;
        RECT -129.205 -90.535 -129.035 -90.365 ;
        RECT -122.045 -90.535 -121.875 -90.365 ;
        RECT -121.585 -90.535 -121.415 -90.365 ;
        RECT -121.125 -90.535 -120.955 -90.365 ;
        RECT -120.665 -90.535 -120.495 -90.365 ;
        RECT -120.205 -90.535 -120.035 -90.365 ;
        RECT -119.745 -90.535 -119.575 -90.365 ;
        RECT -119.285 -90.535 -119.115 -90.365 ;
        RECT -112.125 -90.535 -111.955 -90.365 ;
        RECT -111.665 -90.535 -111.495 -90.365 ;
        RECT -111.205 -90.535 -111.035 -90.365 ;
        RECT -110.745 -90.535 -110.575 -90.365 ;
        RECT -110.285 -90.535 -110.115 -90.365 ;
        RECT -109.825 -90.535 -109.655 -90.365 ;
        RECT -109.365 -90.535 -109.195 -90.365 ;
        RECT -102.205 -90.535 -102.035 -90.365 ;
        RECT -101.745 -90.535 -101.575 -90.365 ;
        RECT -101.285 -90.535 -101.115 -90.365 ;
        RECT -100.825 -90.535 -100.655 -90.365 ;
        RECT -100.365 -90.535 -100.195 -90.365 ;
        RECT -99.905 -90.535 -99.735 -90.365 ;
        RECT -99.445 -90.535 -99.275 -90.365 ;
        RECT -92.285 -90.535 -92.115 -90.365 ;
        RECT -91.825 -90.535 -91.655 -90.365 ;
        RECT -91.365 -90.535 -91.195 -90.365 ;
        RECT -90.905 -90.535 -90.735 -90.365 ;
        RECT -90.445 -90.535 -90.275 -90.365 ;
        RECT -89.985 -90.535 -89.815 -90.365 ;
        RECT -89.525 -90.535 -89.355 -90.365 ;
        RECT -82.365 -90.535 -82.195 -90.365 ;
        RECT -81.905 -90.535 -81.735 -90.365 ;
        RECT -81.445 -90.535 -81.275 -90.365 ;
        RECT -80.985 -90.535 -80.815 -90.365 ;
        RECT -80.525 -90.535 -80.355 -90.365 ;
        RECT -80.065 -90.535 -79.895 -90.365 ;
        RECT -79.605 -90.535 -79.435 -90.365 ;
        RECT -72.445 -90.535 -72.275 -90.365 ;
        RECT -71.985 -90.535 -71.815 -90.365 ;
        RECT -71.525 -90.535 -71.355 -90.365 ;
        RECT -71.065 -90.535 -70.895 -90.365 ;
        RECT -70.605 -90.535 -70.435 -90.365 ;
        RECT -70.145 -90.535 -69.975 -90.365 ;
        RECT -69.685 -90.535 -69.515 -90.365 ;
        RECT -62.525 -90.535 -62.355 -90.365 ;
        RECT -62.065 -90.535 -61.895 -90.365 ;
        RECT -61.605 -90.535 -61.435 -90.365 ;
        RECT -61.145 -90.535 -60.975 -90.365 ;
        RECT -60.685 -90.535 -60.515 -90.365 ;
        RECT -60.225 -90.535 -60.055 -90.365 ;
        RECT -59.765 -90.535 -59.595 -90.365 ;
        RECT -52.605 -90.535 -52.435 -90.365 ;
        RECT -52.145 -90.535 -51.975 -90.365 ;
        RECT -51.685 -90.535 -51.515 -90.365 ;
        RECT -51.225 -90.535 -51.055 -90.365 ;
        RECT -50.765 -90.535 -50.595 -90.365 ;
        RECT -50.305 -90.535 -50.135 -90.365 ;
        RECT -49.845 -90.535 -49.675 -90.365 ;
        RECT -42.685 -90.535 -42.515 -90.365 ;
        RECT -42.225 -90.535 -42.055 -90.365 ;
        RECT -41.765 -90.535 -41.595 -90.365 ;
        RECT -41.305 -90.535 -41.135 -90.365 ;
        RECT -40.845 -90.535 -40.675 -90.365 ;
        RECT -40.385 -90.535 -40.215 -90.365 ;
        RECT -39.925 -90.535 -39.755 -90.365 ;
        RECT -32.765 -90.535 -32.595 -90.365 ;
        RECT -32.305 -90.535 -32.135 -90.365 ;
        RECT -31.845 -90.535 -31.675 -90.365 ;
        RECT -31.385 -90.535 -31.215 -90.365 ;
        RECT -30.925 -90.535 -30.755 -90.365 ;
        RECT -30.465 -90.535 -30.295 -90.365 ;
        RECT -30.005 -90.535 -29.835 -90.365 ;
        RECT -22.845 -90.535 -22.675 -90.365 ;
        RECT -22.385 -90.535 -22.215 -90.365 ;
        RECT -21.925 -90.535 -21.755 -90.365 ;
        RECT -21.465 -90.535 -21.295 -90.365 ;
        RECT -21.005 -90.535 -20.835 -90.365 ;
        RECT -20.545 -90.535 -20.375 -90.365 ;
        RECT -20.085 -90.535 -19.915 -90.365 ;
        RECT -12.925 -90.535 -12.755 -90.365 ;
        RECT -12.465 -90.535 -12.295 -90.365 ;
        RECT -12.005 -90.535 -11.835 -90.365 ;
        RECT -11.545 -90.535 -11.375 -90.365 ;
        RECT -11.085 -90.535 -10.915 -90.365 ;
        RECT -10.625 -90.535 -10.455 -90.365 ;
        RECT -10.165 -90.535 -9.995 -90.365 ;
        RECT -3.005 -90.535 -2.835 -90.365 ;
        RECT -2.545 -90.535 -2.375 -90.365 ;
        RECT -2.085 -90.535 -1.915 -90.365 ;
        RECT -1.625 -90.535 -1.455 -90.365 ;
        RECT -1.165 -90.535 -0.995 -90.365 ;
        RECT -0.705 -90.535 -0.535 -90.365 ;
        RECT -0.245 -90.535 -0.075 -90.365 ;
        RECT 6.915 -90.535 7.085 -90.365 ;
        RECT 7.375 -90.535 7.545 -90.365 ;
        RECT 7.835 -90.535 8.005 -90.365 ;
        RECT 8.295 -90.535 8.465 -90.365 ;
        RECT 8.755 -90.535 8.925 -90.365 ;
        RECT 9.215 -90.535 9.385 -90.365 ;
        RECT 9.675 -90.535 9.845 -90.365 ;
        RECT 16.835 -90.535 17.005 -90.365 ;
        RECT 17.295 -90.535 17.465 -90.365 ;
        RECT 17.755 -90.535 17.925 -90.365 ;
        RECT 18.215 -90.535 18.385 -90.365 ;
        RECT 18.675 -90.535 18.845 -90.365 ;
        RECT 19.135 -90.535 19.305 -90.365 ;
        RECT 19.595 -90.535 19.765 -90.365 ;
        RECT 26.755 -90.535 26.925 -90.365 ;
        RECT 27.215 -90.535 27.385 -90.365 ;
        RECT 27.675 -90.535 27.845 -90.365 ;
        RECT 28.135 -90.535 28.305 -90.365 ;
        RECT -284.815 -91.195 -284.645 -91.025 ;
        RECT -284.345 -91.120 -284.175 -90.950 ;
        RECT -284.815 -91.655 -284.645 -91.485 ;
        RECT -284.815 -92.115 -284.645 -91.945 ;
        RECT -283.875 -91.195 -283.705 -91.025 ;
        RECT -274.895 -91.195 -274.725 -91.025 ;
        RECT -274.425 -91.120 -274.255 -90.950 ;
        RECT -283.875 -91.655 -283.705 -91.485 ;
        RECT -274.895 -91.655 -274.725 -91.485 ;
        RECT -283.875 -92.115 -283.705 -91.945 ;
        RECT -274.895 -92.115 -274.725 -91.945 ;
        RECT -273.955 -91.195 -273.785 -91.025 ;
        RECT -264.975 -91.195 -264.805 -91.025 ;
        RECT -264.505 -91.120 -264.335 -90.950 ;
        RECT -273.955 -91.655 -273.785 -91.485 ;
        RECT -264.975 -91.655 -264.805 -91.485 ;
        RECT -273.955 -92.115 -273.785 -91.945 ;
        RECT -264.975 -92.115 -264.805 -91.945 ;
        RECT -264.035 -91.195 -263.865 -91.025 ;
        RECT -255.055 -91.195 -254.885 -91.025 ;
        RECT -254.585 -91.120 -254.415 -90.950 ;
        RECT -264.035 -91.655 -263.865 -91.485 ;
        RECT -255.055 -91.655 -254.885 -91.485 ;
        RECT -264.035 -92.115 -263.865 -91.945 ;
        RECT -255.055 -92.115 -254.885 -91.945 ;
        RECT -254.115 -91.195 -253.945 -91.025 ;
        RECT -245.135 -91.195 -244.965 -91.025 ;
        RECT -244.665 -91.120 -244.495 -90.950 ;
        RECT -254.115 -91.655 -253.945 -91.485 ;
        RECT -245.135 -91.655 -244.965 -91.485 ;
        RECT -254.115 -92.115 -253.945 -91.945 ;
        RECT -245.135 -92.115 -244.965 -91.945 ;
        RECT -244.195 -91.195 -244.025 -91.025 ;
        RECT -235.215 -91.195 -235.045 -91.025 ;
        RECT -234.745 -91.120 -234.575 -90.950 ;
        RECT -244.195 -91.655 -244.025 -91.485 ;
        RECT -235.215 -91.655 -235.045 -91.485 ;
        RECT -244.195 -92.115 -244.025 -91.945 ;
        RECT -235.215 -92.115 -235.045 -91.945 ;
        RECT -234.275 -91.195 -234.105 -91.025 ;
        RECT -225.295 -91.195 -225.125 -91.025 ;
        RECT -224.825 -91.120 -224.655 -90.950 ;
        RECT -234.275 -91.655 -234.105 -91.485 ;
        RECT -225.295 -91.655 -225.125 -91.485 ;
        RECT -234.275 -92.115 -234.105 -91.945 ;
        RECT -225.295 -92.115 -225.125 -91.945 ;
        RECT -224.355 -91.195 -224.185 -91.025 ;
        RECT -215.375 -91.195 -215.205 -91.025 ;
        RECT -214.905 -91.120 -214.735 -90.950 ;
        RECT -224.355 -91.655 -224.185 -91.485 ;
        RECT -215.375 -91.655 -215.205 -91.485 ;
        RECT -224.355 -92.115 -224.185 -91.945 ;
        RECT -215.375 -92.115 -215.205 -91.945 ;
        RECT -214.435 -91.195 -214.265 -91.025 ;
        RECT -205.455 -91.195 -205.285 -91.025 ;
        RECT -204.985 -91.120 -204.815 -90.950 ;
        RECT -214.435 -91.655 -214.265 -91.485 ;
        RECT -205.455 -91.655 -205.285 -91.485 ;
        RECT -214.435 -92.115 -214.265 -91.945 ;
        RECT -205.455 -92.115 -205.285 -91.945 ;
        RECT -204.515 -91.195 -204.345 -91.025 ;
        RECT -195.535 -91.195 -195.365 -91.025 ;
        RECT -195.065 -91.120 -194.895 -90.950 ;
        RECT -204.515 -91.655 -204.345 -91.485 ;
        RECT -195.535 -91.655 -195.365 -91.485 ;
        RECT -204.515 -92.115 -204.345 -91.945 ;
        RECT -195.535 -92.115 -195.365 -91.945 ;
        RECT -194.595 -91.195 -194.425 -91.025 ;
        RECT -185.615 -91.195 -185.445 -91.025 ;
        RECT -185.145 -91.120 -184.975 -90.950 ;
        RECT -194.595 -91.655 -194.425 -91.485 ;
        RECT -185.615 -91.655 -185.445 -91.485 ;
        RECT -194.595 -92.115 -194.425 -91.945 ;
        RECT -185.615 -92.115 -185.445 -91.945 ;
        RECT -184.675 -91.195 -184.505 -91.025 ;
        RECT -175.695 -91.195 -175.525 -91.025 ;
        RECT -175.225 -91.120 -175.055 -90.950 ;
        RECT -184.675 -91.655 -184.505 -91.485 ;
        RECT -175.695 -91.655 -175.525 -91.485 ;
        RECT -184.675 -92.115 -184.505 -91.945 ;
        RECT -175.695 -92.115 -175.525 -91.945 ;
        RECT -174.755 -91.195 -174.585 -91.025 ;
        RECT -165.775 -91.195 -165.605 -91.025 ;
        RECT -165.305 -91.120 -165.135 -90.950 ;
        RECT -174.755 -91.655 -174.585 -91.485 ;
        RECT -165.775 -91.655 -165.605 -91.485 ;
        RECT -174.755 -92.115 -174.585 -91.945 ;
        RECT -165.775 -92.115 -165.605 -91.945 ;
        RECT -164.835 -91.195 -164.665 -91.025 ;
        RECT -155.855 -91.195 -155.685 -91.025 ;
        RECT -155.385 -91.120 -155.215 -90.950 ;
        RECT -164.835 -91.655 -164.665 -91.485 ;
        RECT -155.855 -91.655 -155.685 -91.485 ;
        RECT -164.835 -92.115 -164.665 -91.945 ;
        RECT -155.855 -92.115 -155.685 -91.945 ;
        RECT -154.915 -91.195 -154.745 -91.025 ;
        RECT -145.935 -91.195 -145.765 -91.025 ;
        RECT -145.465 -91.120 -145.295 -90.950 ;
        RECT -154.915 -91.655 -154.745 -91.485 ;
        RECT -145.935 -91.655 -145.765 -91.485 ;
        RECT -154.915 -92.115 -154.745 -91.945 ;
        RECT -145.935 -92.115 -145.765 -91.945 ;
        RECT -144.995 -91.195 -144.825 -91.025 ;
        RECT -136.015 -91.195 -135.845 -91.025 ;
        RECT -135.545 -91.120 -135.375 -90.950 ;
        RECT -144.995 -91.655 -144.825 -91.485 ;
        RECT -136.015 -91.655 -135.845 -91.485 ;
        RECT -144.995 -92.115 -144.825 -91.945 ;
        RECT -136.015 -92.115 -135.845 -91.945 ;
        RECT -135.075 -91.195 -134.905 -91.025 ;
        RECT -126.095 -91.195 -125.925 -91.025 ;
        RECT -125.625 -91.120 -125.455 -90.950 ;
        RECT -135.075 -91.655 -134.905 -91.485 ;
        RECT -126.095 -91.655 -125.925 -91.485 ;
        RECT -135.075 -92.115 -134.905 -91.945 ;
        RECT -126.095 -92.115 -125.925 -91.945 ;
        RECT -125.155 -91.195 -124.985 -91.025 ;
        RECT -116.175 -91.195 -116.005 -91.025 ;
        RECT -115.705 -91.120 -115.535 -90.950 ;
        RECT -125.155 -91.655 -124.985 -91.485 ;
        RECT -116.175 -91.655 -116.005 -91.485 ;
        RECT -125.155 -92.115 -124.985 -91.945 ;
        RECT -116.175 -92.115 -116.005 -91.945 ;
        RECT -115.235 -91.195 -115.065 -91.025 ;
        RECT -106.255 -91.195 -106.085 -91.025 ;
        RECT -105.785 -91.120 -105.615 -90.950 ;
        RECT -115.235 -91.655 -115.065 -91.485 ;
        RECT -106.255 -91.655 -106.085 -91.485 ;
        RECT -115.235 -92.115 -115.065 -91.945 ;
        RECT -106.255 -92.115 -106.085 -91.945 ;
        RECT -105.315 -91.195 -105.145 -91.025 ;
        RECT -96.335 -91.195 -96.165 -91.025 ;
        RECT -95.865 -91.120 -95.695 -90.950 ;
        RECT -105.315 -91.655 -105.145 -91.485 ;
        RECT -96.335 -91.655 -96.165 -91.485 ;
        RECT -105.315 -92.115 -105.145 -91.945 ;
        RECT -96.335 -92.115 -96.165 -91.945 ;
        RECT -95.395 -91.195 -95.225 -91.025 ;
        RECT -86.415 -91.195 -86.245 -91.025 ;
        RECT -85.945 -91.120 -85.775 -90.950 ;
        RECT -95.395 -91.655 -95.225 -91.485 ;
        RECT -86.415 -91.655 -86.245 -91.485 ;
        RECT -95.395 -92.115 -95.225 -91.945 ;
        RECT -86.415 -92.115 -86.245 -91.945 ;
        RECT -85.475 -91.195 -85.305 -91.025 ;
        RECT -76.495 -91.195 -76.325 -91.025 ;
        RECT -76.025 -91.120 -75.855 -90.950 ;
        RECT -85.475 -91.655 -85.305 -91.485 ;
        RECT -76.495 -91.655 -76.325 -91.485 ;
        RECT -85.475 -92.115 -85.305 -91.945 ;
        RECT -76.495 -92.115 -76.325 -91.945 ;
        RECT -75.555 -91.195 -75.385 -91.025 ;
        RECT -66.575 -91.195 -66.405 -91.025 ;
        RECT -66.105 -91.120 -65.935 -90.950 ;
        RECT -75.555 -91.655 -75.385 -91.485 ;
        RECT -66.575 -91.655 -66.405 -91.485 ;
        RECT -75.555 -92.115 -75.385 -91.945 ;
        RECT -66.575 -92.115 -66.405 -91.945 ;
        RECT -65.635 -91.195 -65.465 -91.025 ;
        RECT -56.655 -91.195 -56.485 -91.025 ;
        RECT -56.185 -91.120 -56.015 -90.950 ;
        RECT -65.635 -91.655 -65.465 -91.485 ;
        RECT -56.655 -91.655 -56.485 -91.485 ;
        RECT -65.635 -92.115 -65.465 -91.945 ;
        RECT -56.655 -92.115 -56.485 -91.945 ;
        RECT -55.715 -91.195 -55.545 -91.025 ;
        RECT -46.735 -91.195 -46.565 -91.025 ;
        RECT -46.265 -91.120 -46.095 -90.950 ;
        RECT -55.715 -91.655 -55.545 -91.485 ;
        RECT -46.735 -91.655 -46.565 -91.485 ;
        RECT -55.715 -92.115 -55.545 -91.945 ;
        RECT -46.735 -92.115 -46.565 -91.945 ;
        RECT -45.795 -91.195 -45.625 -91.025 ;
        RECT -36.815 -91.195 -36.645 -91.025 ;
        RECT -36.345 -91.120 -36.175 -90.950 ;
        RECT -45.795 -91.655 -45.625 -91.485 ;
        RECT -36.815 -91.655 -36.645 -91.485 ;
        RECT -45.795 -92.115 -45.625 -91.945 ;
        RECT -36.815 -92.115 -36.645 -91.945 ;
        RECT -35.875 -91.195 -35.705 -91.025 ;
        RECT -26.895 -91.195 -26.725 -91.025 ;
        RECT -26.425 -91.120 -26.255 -90.950 ;
        RECT -35.875 -91.655 -35.705 -91.485 ;
        RECT -26.895 -91.655 -26.725 -91.485 ;
        RECT -35.875 -92.115 -35.705 -91.945 ;
        RECT -26.895 -92.115 -26.725 -91.945 ;
        RECT -25.955 -91.195 -25.785 -91.025 ;
        RECT -16.975 -91.195 -16.805 -91.025 ;
        RECT -16.505 -91.120 -16.335 -90.950 ;
        RECT -25.955 -91.655 -25.785 -91.485 ;
        RECT -16.975 -91.655 -16.805 -91.485 ;
        RECT -25.955 -92.115 -25.785 -91.945 ;
        RECT -16.975 -92.115 -16.805 -91.945 ;
        RECT -16.035 -91.195 -15.865 -91.025 ;
        RECT -7.055 -91.195 -6.885 -91.025 ;
        RECT -6.585 -91.120 -6.415 -90.950 ;
        RECT -16.035 -91.655 -15.865 -91.485 ;
        RECT -7.055 -91.655 -6.885 -91.485 ;
        RECT -16.035 -92.115 -15.865 -91.945 ;
        RECT -7.055 -92.115 -6.885 -91.945 ;
        RECT -6.115 -91.195 -5.945 -91.025 ;
        RECT 2.865 -91.195 3.035 -91.025 ;
        RECT 3.335 -91.120 3.505 -90.950 ;
        RECT -6.115 -91.655 -5.945 -91.485 ;
        RECT 2.865 -91.655 3.035 -91.485 ;
        RECT -6.115 -92.115 -5.945 -91.945 ;
        RECT 2.865 -92.115 3.035 -91.945 ;
        RECT 3.805 -91.195 3.975 -91.025 ;
        RECT 12.785 -91.195 12.955 -91.025 ;
        RECT 13.255 -91.120 13.425 -90.950 ;
        RECT 3.805 -91.655 3.975 -91.485 ;
        RECT 12.785 -91.655 12.955 -91.485 ;
        RECT 3.805 -92.115 3.975 -91.945 ;
        RECT 12.785 -92.115 12.955 -91.945 ;
        RECT 13.725 -91.195 13.895 -91.025 ;
        RECT 22.705 -91.195 22.875 -91.025 ;
        RECT 23.175 -91.120 23.345 -90.950 ;
        RECT 13.725 -91.655 13.895 -91.485 ;
        RECT 22.705 -91.655 22.875 -91.485 ;
        RECT 13.725 -92.115 13.895 -91.945 ;
        RECT 22.705 -92.115 22.875 -91.945 ;
        RECT 23.645 -91.195 23.815 -91.025 ;
        RECT 23.645 -91.655 23.815 -91.485 ;
        RECT 23.645 -92.115 23.815 -91.945 ;
        RECT -279.605 -173.945 -279.435 -173.775 ;
        RECT -279.135 -173.950 -278.965 -173.780 ;
        RECT -278.665 -173.945 -278.495 -173.775 ;
        RECT -279.605 -174.405 -279.435 -174.235 ;
        RECT -279.605 -174.865 -279.435 -174.695 ;
        RECT -269.685 -173.945 -269.515 -173.775 ;
        RECT -269.215 -173.950 -269.045 -173.780 ;
        RECT -268.745 -173.945 -268.575 -173.775 ;
        RECT -278.665 -174.405 -278.495 -174.235 ;
        RECT -269.685 -174.405 -269.515 -174.235 ;
        RECT -278.665 -174.865 -278.495 -174.695 ;
        RECT -269.685 -174.865 -269.515 -174.695 ;
        RECT -259.765 -173.945 -259.595 -173.775 ;
        RECT -259.295 -173.950 -259.125 -173.780 ;
        RECT -258.825 -173.945 -258.655 -173.775 ;
        RECT -268.745 -174.405 -268.575 -174.235 ;
        RECT -259.765 -174.405 -259.595 -174.235 ;
        RECT -268.745 -174.865 -268.575 -174.695 ;
        RECT -259.765 -174.865 -259.595 -174.695 ;
        RECT -249.845 -173.945 -249.675 -173.775 ;
        RECT -249.375 -173.950 -249.205 -173.780 ;
        RECT -248.905 -173.945 -248.735 -173.775 ;
        RECT -258.825 -174.405 -258.655 -174.235 ;
        RECT -249.845 -174.405 -249.675 -174.235 ;
        RECT -258.825 -174.865 -258.655 -174.695 ;
        RECT -249.845 -174.865 -249.675 -174.695 ;
        RECT -239.925 -173.945 -239.755 -173.775 ;
        RECT -239.455 -173.950 -239.285 -173.780 ;
        RECT -238.985 -173.945 -238.815 -173.775 ;
        RECT -248.905 -174.405 -248.735 -174.235 ;
        RECT -239.925 -174.405 -239.755 -174.235 ;
        RECT -248.905 -174.865 -248.735 -174.695 ;
        RECT -239.925 -174.865 -239.755 -174.695 ;
        RECT -230.005 -173.945 -229.835 -173.775 ;
        RECT -229.535 -173.950 -229.365 -173.780 ;
        RECT -229.065 -173.945 -228.895 -173.775 ;
        RECT -238.985 -174.405 -238.815 -174.235 ;
        RECT -230.005 -174.405 -229.835 -174.235 ;
        RECT -238.985 -174.865 -238.815 -174.695 ;
        RECT -230.005 -174.865 -229.835 -174.695 ;
        RECT -220.085 -173.945 -219.915 -173.775 ;
        RECT -219.615 -173.950 -219.445 -173.780 ;
        RECT -219.145 -173.945 -218.975 -173.775 ;
        RECT -229.065 -174.405 -228.895 -174.235 ;
        RECT -220.085 -174.405 -219.915 -174.235 ;
        RECT -229.065 -174.865 -228.895 -174.695 ;
        RECT -220.085 -174.865 -219.915 -174.695 ;
        RECT -210.165 -173.945 -209.995 -173.775 ;
        RECT -209.695 -173.950 -209.525 -173.780 ;
        RECT -209.225 -173.945 -209.055 -173.775 ;
        RECT -219.145 -174.405 -218.975 -174.235 ;
        RECT -210.165 -174.405 -209.995 -174.235 ;
        RECT -219.145 -174.865 -218.975 -174.695 ;
        RECT -210.165 -174.865 -209.995 -174.695 ;
        RECT -200.245 -173.945 -200.075 -173.775 ;
        RECT -199.775 -173.950 -199.605 -173.780 ;
        RECT -199.305 -173.945 -199.135 -173.775 ;
        RECT -209.225 -174.405 -209.055 -174.235 ;
        RECT -200.245 -174.405 -200.075 -174.235 ;
        RECT -209.225 -174.865 -209.055 -174.695 ;
        RECT -200.245 -174.865 -200.075 -174.695 ;
        RECT -190.325 -173.945 -190.155 -173.775 ;
        RECT -189.855 -173.950 -189.685 -173.780 ;
        RECT -189.385 -173.945 -189.215 -173.775 ;
        RECT -199.305 -174.405 -199.135 -174.235 ;
        RECT -190.325 -174.405 -190.155 -174.235 ;
        RECT -199.305 -174.865 -199.135 -174.695 ;
        RECT -190.325 -174.865 -190.155 -174.695 ;
        RECT -180.405 -173.945 -180.235 -173.775 ;
        RECT -179.935 -173.950 -179.765 -173.780 ;
        RECT -179.465 -173.945 -179.295 -173.775 ;
        RECT -189.385 -174.405 -189.215 -174.235 ;
        RECT -180.405 -174.405 -180.235 -174.235 ;
        RECT -189.385 -174.865 -189.215 -174.695 ;
        RECT -180.405 -174.865 -180.235 -174.695 ;
        RECT -170.485 -173.945 -170.315 -173.775 ;
        RECT -170.015 -173.950 -169.845 -173.780 ;
        RECT -169.545 -173.945 -169.375 -173.775 ;
        RECT -179.465 -174.405 -179.295 -174.235 ;
        RECT -170.485 -174.405 -170.315 -174.235 ;
        RECT -179.465 -174.865 -179.295 -174.695 ;
        RECT -170.485 -174.865 -170.315 -174.695 ;
        RECT -160.565 -173.945 -160.395 -173.775 ;
        RECT -160.095 -173.950 -159.925 -173.780 ;
        RECT -159.625 -173.945 -159.455 -173.775 ;
        RECT -169.545 -174.405 -169.375 -174.235 ;
        RECT -160.565 -174.405 -160.395 -174.235 ;
        RECT -169.545 -174.865 -169.375 -174.695 ;
        RECT -160.565 -174.865 -160.395 -174.695 ;
        RECT -150.645 -173.945 -150.475 -173.775 ;
        RECT -150.175 -173.950 -150.005 -173.780 ;
        RECT -149.705 -173.945 -149.535 -173.775 ;
        RECT -159.625 -174.405 -159.455 -174.235 ;
        RECT -150.645 -174.405 -150.475 -174.235 ;
        RECT -159.625 -174.865 -159.455 -174.695 ;
        RECT -150.645 -174.865 -150.475 -174.695 ;
        RECT -140.725 -173.945 -140.555 -173.775 ;
        RECT -140.255 -173.950 -140.085 -173.780 ;
        RECT -139.785 -173.945 -139.615 -173.775 ;
        RECT -149.705 -174.405 -149.535 -174.235 ;
        RECT -140.725 -174.405 -140.555 -174.235 ;
        RECT -149.705 -174.865 -149.535 -174.695 ;
        RECT -140.725 -174.865 -140.555 -174.695 ;
        RECT -130.805 -173.945 -130.635 -173.775 ;
        RECT -130.335 -173.950 -130.165 -173.780 ;
        RECT -129.865 -173.945 -129.695 -173.775 ;
        RECT -139.785 -174.405 -139.615 -174.235 ;
        RECT -130.805 -174.405 -130.635 -174.235 ;
        RECT -139.785 -174.865 -139.615 -174.695 ;
        RECT -130.805 -174.865 -130.635 -174.695 ;
        RECT -120.885 -173.945 -120.715 -173.775 ;
        RECT -120.415 -173.950 -120.245 -173.780 ;
        RECT -119.945 -173.945 -119.775 -173.775 ;
        RECT -129.865 -174.405 -129.695 -174.235 ;
        RECT -120.885 -174.405 -120.715 -174.235 ;
        RECT -129.865 -174.865 -129.695 -174.695 ;
        RECT -120.885 -174.865 -120.715 -174.695 ;
        RECT -110.965 -173.945 -110.795 -173.775 ;
        RECT -110.495 -173.950 -110.325 -173.780 ;
        RECT -110.025 -173.945 -109.855 -173.775 ;
        RECT -119.945 -174.405 -119.775 -174.235 ;
        RECT -110.965 -174.405 -110.795 -174.235 ;
        RECT -119.945 -174.865 -119.775 -174.695 ;
        RECT -110.965 -174.865 -110.795 -174.695 ;
        RECT -101.045 -173.945 -100.875 -173.775 ;
        RECT -100.575 -173.950 -100.405 -173.780 ;
        RECT -100.105 -173.945 -99.935 -173.775 ;
        RECT -110.025 -174.405 -109.855 -174.235 ;
        RECT -101.045 -174.405 -100.875 -174.235 ;
        RECT -110.025 -174.865 -109.855 -174.695 ;
        RECT -101.045 -174.865 -100.875 -174.695 ;
        RECT -91.125 -173.945 -90.955 -173.775 ;
        RECT -90.655 -173.950 -90.485 -173.780 ;
        RECT -90.185 -173.945 -90.015 -173.775 ;
        RECT -100.105 -174.405 -99.935 -174.235 ;
        RECT -91.125 -174.405 -90.955 -174.235 ;
        RECT -100.105 -174.865 -99.935 -174.695 ;
        RECT -91.125 -174.865 -90.955 -174.695 ;
        RECT -81.205 -173.945 -81.035 -173.775 ;
        RECT -80.735 -173.950 -80.565 -173.780 ;
        RECT -80.265 -173.945 -80.095 -173.775 ;
        RECT -90.185 -174.405 -90.015 -174.235 ;
        RECT -81.205 -174.405 -81.035 -174.235 ;
        RECT -90.185 -174.865 -90.015 -174.695 ;
        RECT -81.205 -174.865 -81.035 -174.695 ;
        RECT -71.285 -173.945 -71.115 -173.775 ;
        RECT -70.815 -173.950 -70.645 -173.780 ;
        RECT -70.345 -173.945 -70.175 -173.775 ;
        RECT -80.265 -174.405 -80.095 -174.235 ;
        RECT -71.285 -174.405 -71.115 -174.235 ;
        RECT -80.265 -174.865 -80.095 -174.695 ;
        RECT -71.285 -174.865 -71.115 -174.695 ;
        RECT -61.365 -173.945 -61.195 -173.775 ;
        RECT -60.895 -173.950 -60.725 -173.780 ;
        RECT -60.425 -173.945 -60.255 -173.775 ;
        RECT -70.345 -174.405 -70.175 -174.235 ;
        RECT -61.365 -174.405 -61.195 -174.235 ;
        RECT -70.345 -174.865 -70.175 -174.695 ;
        RECT -61.365 -174.865 -61.195 -174.695 ;
        RECT -51.445 -173.945 -51.275 -173.775 ;
        RECT -50.975 -173.950 -50.805 -173.780 ;
        RECT -50.505 -173.945 -50.335 -173.775 ;
        RECT -60.425 -174.405 -60.255 -174.235 ;
        RECT -51.445 -174.405 -51.275 -174.235 ;
        RECT -60.425 -174.865 -60.255 -174.695 ;
        RECT -51.445 -174.865 -51.275 -174.695 ;
        RECT -41.525 -173.945 -41.355 -173.775 ;
        RECT -41.055 -173.950 -40.885 -173.780 ;
        RECT -40.585 -173.945 -40.415 -173.775 ;
        RECT -50.505 -174.405 -50.335 -174.235 ;
        RECT -41.525 -174.405 -41.355 -174.235 ;
        RECT -50.505 -174.865 -50.335 -174.695 ;
        RECT -41.525 -174.865 -41.355 -174.695 ;
        RECT -31.605 -173.945 -31.435 -173.775 ;
        RECT -31.135 -173.950 -30.965 -173.780 ;
        RECT -30.665 -173.945 -30.495 -173.775 ;
        RECT -40.585 -174.405 -40.415 -174.235 ;
        RECT -31.605 -174.405 -31.435 -174.235 ;
        RECT -40.585 -174.865 -40.415 -174.695 ;
        RECT -31.605 -174.865 -31.435 -174.695 ;
        RECT -21.685 -173.945 -21.515 -173.775 ;
        RECT -21.215 -173.950 -21.045 -173.780 ;
        RECT -20.745 -173.945 -20.575 -173.775 ;
        RECT -30.665 -174.405 -30.495 -174.235 ;
        RECT -21.685 -174.405 -21.515 -174.235 ;
        RECT -30.665 -174.865 -30.495 -174.695 ;
        RECT -21.685 -174.865 -21.515 -174.695 ;
        RECT -11.765 -173.945 -11.595 -173.775 ;
        RECT -11.295 -173.950 -11.125 -173.780 ;
        RECT -10.825 -173.945 -10.655 -173.775 ;
        RECT -20.745 -174.405 -20.575 -174.235 ;
        RECT -11.765 -174.405 -11.595 -174.235 ;
        RECT -20.745 -174.865 -20.575 -174.695 ;
        RECT -11.765 -174.865 -11.595 -174.695 ;
        RECT -1.845 -173.945 -1.675 -173.775 ;
        RECT -1.375 -173.950 -1.205 -173.780 ;
        RECT -0.905 -173.945 -0.735 -173.775 ;
        RECT -10.825 -174.405 -10.655 -174.235 ;
        RECT -1.845 -174.405 -1.675 -174.235 ;
        RECT -10.825 -174.865 -10.655 -174.695 ;
        RECT -1.845 -174.865 -1.675 -174.695 ;
        RECT 8.075 -173.945 8.245 -173.775 ;
        RECT 8.545 -173.950 8.715 -173.780 ;
        RECT 9.015 -173.945 9.185 -173.775 ;
        RECT -0.905 -174.405 -0.735 -174.235 ;
        RECT 8.075 -174.405 8.245 -174.235 ;
        RECT -0.905 -174.865 -0.735 -174.695 ;
        RECT 8.075 -174.865 8.245 -174.695 ;
        RECT 17.995 -173.945 18.165 -173.775 ;
        RECT 18.465 -173.950 18.635 -173.780 ;
        RECT 18.935 -173.945 19.105 -173.775 ;
        RECT 9.015 -174.405 9.185 -174.235 ;
        RECT 17.995 -174.405 18.165 -174.235 ;
        RECT 9.015 -174.865 9.185 -174.695 ;
        RECT 17.995 -174.865 18.165 -174.695 ;
        RECT 27.915 -173.945 28.085 -173.775 ;
        RECT 28.385 -173.950 28.555 -173.780 ;
        RECT 18.935 -174.405 19.105 -174.235 ;
        RECT 27.915 -174.405 28.085 -174.235 ;
        RECT 18.935 -174.865 19.105 -174.695 ;
        RECT 27.915 -174.865 28.085 -174.695 ;
        RECT -285.475 -175.525 -285.305 -175.355 ;
        RECT -285.015 -175.525 -284.845 -175.355 ;
        RECT -284.555 -175.525 -284.385 -175.355 ;
        RECT -284.095 -175.525 -283.925 -175.355 ;
        RECT -283.635 -175.525 -283.465 -175.355 ;
        RECT -283.175 -175.525 -283.005 -175.355 ;
        RECT -282.715 -175.525 -282.545 -175.355 ;
        RECT -275.555 -175.525 -275.385 -175.355 ;
        RECT -275.095 -175.525 -274.925 -175.355 ;
        RECT -274.635 -175.525 -274.465 -175.355 ;
        RECT -274.175 -175.525 -274.005 -175.355 ;
        RECT -273.715 -175.525 -273.545 -175.355 ;
        RECT -273.255 -175.525 -273.085 -175.355 ;
        RECT -272.795 -175.525 -272.625 -175.355 ;
        RECT -265.635 -175.525 -265.465 -175.355 ;
        RECT -265.175 -175.525 -265.005 -175.355 ;
        RECT -264.715 -175.525 -264.545 -175.355 ;
        RECT -264.255 -175.525 -264.085 -175.355 ;
        RECT -263.795 -175.525 -263.625 -175.355 ;
        RECT -263.335 -175.525 -263.165 -175.355 ;
        RECT -262.875 -175.525 -262.705 -175.355 ;
        RECT -255.715 -175.525 -255.545 -175.355 ;
        RECT -255.255 -175.525 -255.085 -175.355 ;
        RECT -254.795 -175.525 -254.625 -175.355 ;
        RECT -254.335 -175.525 -254.165 -175.355 ;
        RECT -253.875 -175.525 -253.705 -175.355 ;
        RECT -253.415 -175.525 -253.245 -175.355 ;
        RECT -252.955 -175.525 -252.785 -175.355 ;
        RECT -245.795 -175.525 -245.625 -175.355 ;
        RECT -245.335 -175.525 -245.165 -175.355 ;
        RECT -244.875 -175.525 -244.705 -175.355 ;
        RECT -244.415 -175.525 -244.245 -175.355 ;
        RECT -243.955 -175.525 -243.785 -175.355 ;
        RECT -243.495 -175.525 -243.325 -175.355 ;
        RECT -243.035 -175.525 -242.865 -175.355 ;
        RECT -235.875 -175.525 -235.705 -175.355 ;
        RECT -235.415 -175.525 -235.245 -175.355 ;
        RECT -234.955 -175.525 -234.785 -175.355 ;
        RECT -234.495 -175.525 -234.325 -175.355 ;
        RECT -234.035 -175.525 -233.865 -175.355 ;
        RECT -233.575 -175.525 -233.405 -175.355 ;
        RECT -233.115 -175.525 -232.945 -175.355 ;
        RECT -225.955 -175.525 -225.785 -175.355 ;
        RECT -225.495 -175.525 -225.325 -175.355 ;
        RECT -225.035 -175.525 -224.865 -175.355 ;
        RECT -224.575 -175.525 -224.405 -175.355 ;
        RECT -224.115 -175.525 -223.945 -175.355 ;
        RECT -223.655 -175.525 -223.485 -175.355 ;
        RECT -223.195 -175.525 -223.025 -175.355 ;
        RECT -216.035 -175.525 -215.865 -175.355 ;
        RECT -215.575 -175.525 -215.405 -175.355 ;
        RECT -215.115 -175.525 -214.945 -175.355 ;
        RECT -214.655 -175.525 -214.485 -175.355 ;
        RECT -214.195 -175.525 -214.025 -175.355 ;
        RECT -213.735 -175.525 -213.565 -175.355 ;
        RECT -213.275 -175.525 -213.105 -175.355 ;
        RECT -206.115 -175.525 -205.945 -175.355 ;
        RECT -205.655 -175.525 -205.485 -175.355 ;
        RECT -205.195 -175.525 -205.025 -175.355 ;
        RECT -204.735 -175.525 -204.565 -175.355 ;
        RECT -204.275 -175.525 -204.105 -175.355 ;
        RECT -203.815 -175.525 -203.645 -175.355 ;
        RECT -203.355 -175.525 -203.185 -175.355 ;
        RECT -196.195 -175.525 -196.025 -175.355 ;
        RECT -195.735 -175.525 -195.565 -175.355 ;
        RECT -195.275 -175.525 -195.105 -175.355 ;
        RECT -194.815 -175.525 -194.645 -175.355 ;
        RECT -194.355 -175.525 -194.185 -175.355 ;
        RECT -193.895 -175.525 -193.725 -175.355 ;
        RECT -193.435 -175.525 -193.265 -175.355 ;
        RECT -186.275 -175.525 -186.105 -175.355 ;
        RECT -185.815 -175.525 -185.645 -175.355 ;
        RECT -185.355 -175.525 -185.185 -175.355 ;
        RECT -184.895 -175.525 -184.725 -175.355 ;
        RECT -184.435 -175.525 -184.265 -175.355 ;
        RECT -183.975 -175.525 -183.805 -175.355 ;
        RECT -183.515 -175.525 -183.345 -175.355 ;
        RECT -176.355 -175.525 -176.185 -175.355 ;
        RECT -175.895 -175.525 -175.725 -175.355 ;
        RECT -175.435 -175.525 -175.265 -175.355 ;
        RECT -174.975 -175.525 -174.805 -175.355 ;
        RECT -174.515 -175.525 -174.345 -175.355 ;
        RECT -174.055 -175.525 -173.885 -175.355 ;
        RECT -173.595 -175.525 -173.425 -175.355 ;
        RECT -166.435 -175.525 -166.265 -175.355 ;
        RECT -165.975 -175.525 -165.805 -175.355 ;
        RECT -165.515 -175.525 -165.345 -175.355 ;
        RECT -165.055 -175.525 -164.885 -175.355 ;
        RECT -164.595 -175.525 -164.425 -175.355 ;
        RECT -164.135 -175.525 -163.965 -175.355 ;
        RECT -163.675 -175.525 -163.505 -175.355 ;
        RECT -156.515 -175.525 -156.345 -175.355 ;
        RECT -156.055 -175.525 -155.885 -175.355 ;
        RECT -155.595 -175.525 -155.425 -175.355 ;
        RECT -155.135 -175.525 -154.965 -175.355 ;
        RECT -154.675 -175.525 -154.505 -175.355 ;
        RECT -154.215 -175.525 -154.045 -175.355 ;
        RECT -153.755 -175.525 -153.585 -175.355 ;
        RECT -146.595 -175.525 -146.425 -175.355 ;
        RECT -146.135 -175.525 -145.965 -175.355 ;
        RECT -145.675 -175.525 -145.505 -175.355 ;
        RECT -145.215 -175.525 -145.045 -175.355 ;
        RECT -144.755 -175.525 -144.585 -175.355 ;
        RECT -144.295 -175.525 -144.125 -175.355 ;
        RECT -143.835 -175.525 -143.665 -175.355 ;
        RECT -136.675 -175.525 -136.505 -175.355 ;
        RECT -136.215 -175.525 -136.045 -175.355 ;
        RECT -135.755 -175.525 -135.585 -175.355 ;
        RECT -135.295 -175.525 -135.125 -175.355 ;
        RECT -134.835 -175.525 -134.665 -175.355 ;
        RECT -134.375 -175.525 -134.205 -175.355 ;
        RECT -133.915 -175.525 -133.745 -175.355 ;
        RECT -126.755 -175.525 -126.585 -175.355 ;
        RECT -126.295 -175.525 -126.125 -175.355 ;
        RECT -125.835 -175.525 -125.665 -175.355 ;
        RECT -125.375 -175.525 -125.205 -175.355 ;
        RECT -124.915 -175.525 -124.745 -175.355 ;
        RECT -124.455 -175.525 -124.285 -175.355 ;
        RECT -123.995 -175.525 -123.825 -175.355 ;
        RECT -116.835 -175.525 -116.665 -175.355 ;
        RECT -116.375 -175.525 -116.205 -175.355 ;
        RECT -115.915 -175.525 -115.745 -175.355 ;
        RECT -115.455 -175.525 -115.285 -175.355 ;
        RECT -114.995 -175.525 -114.825 -175.355 ;
        RECT -114.535 -175.525 -114.365 -175.355 ;
        RECT -114.075 -175.525 -113.905 -175.355 ;
        RECT -106.915 -175.525 -106.745 -175.355 ;
        RECT -106.455 -175.525 -106.285 -175.355 ;
        RECT -105.995 -175.525 -105.825 -175.355 ;
        RECT -105.535 -175.525 -105.365 -175.355 ;
        RECT -105.075 -175.525 -104.905 -175.355 ;
        RECT -104.615 -175.525 -104.445 -175.355 ;
        RECT -104.155 -175.525 -103.985 -175.355 ;
        RECT -96.995 -175.525 -96.825 -175.355 ;
        RECT -96.535 -175.525 -96.365 -175.355 ;
        RECT -96.075 -175.525 -95.905 -175.355 ;
        RECT -95.615 -175.525 -95.445 -175.355 ;
        RECT -95.155 -175.525 -94.985 -175.355 ;
        RECT -94.695 -175.525 -94.525 -175.355 ;
        RECT -94.235 -175.525 -94.065 -175.355 ;
        RECT -87.075 -175.525 -86.905 -175.355 ;
        RECT -86.615 -175.525 -86.445 -175.355 ;
        RECT -86.155 -175.525 -85.985 -175.355 ;
        RECT -85.695 -175.525 -85.525 -175.355 ;
        RECT -85.235 -175.525 -85.065 -175.355 ;
        RECT -84.775 -175.525 -84.605 -175.355 ;
        RECT -84.315 -175.525 -84.145 -175.355 ;
        RECT -77.155 -175.525 -76.985 -175.355 ;
        RECT -76.695 -175.525 -76.525 -175.355 ;
        RECT -76.235 -175.525 -76.065 -175.355 ;
        RECT -75.775 -175.525 -75.605 -175.355 ;
        RECT -75.315 -175.525 -75.145 -175.355 ;
        RECT -74.855 -175.525 -74.685 -175.355 ;
        RECT -74.395 -175.525 -74.225 -175.355 ;
        RECT -67.235 -175.525 -67.065 -175.355 ;
        RECT -66.775 -175.525 -66.605 -175.355 ;
        RECT -66.315 -175.525 -66.145 -175.355 ;
        RECT -65.855 -175.525 -65.685 -175.355 ;
        RECT -65.395 -175.525 -65.225 -175.355 ;
        RECT -64.935 -175.525 -64.765 -175.355 ;
        RECT -64.475 -175.525 -64.305 -175.355 ;
        RECT -57.315 -175.525 -57.145 -175.355 ;
        RECT -56.855 -175.525 -56.685 -175.355 ;
        RECT -56.395 -175.525 -56.225 -175.355 ;
        RECT -55.935 -175.525 -55.765 -175.355 ;
        RECT -55.475 -175.525 -55.305 -175.355 ;
        RECT -55.015 -175.525 -54.845 -175.355 ;
        RECT -54.555 -175.525 -54.385 -175.355 ;
        RECT -47.395 -175.525 -47.225 -175.355 ;
        RECT -46.935 -175.525 -46.765 -175.355 ;
        RECT -46.475 -175.525 -46.305 -175.355 ;
        RECT -46.015 -175.525 -45.845 -175.355 ;
        RECT -45.555 -175.525 -45.385 -175.355 ;
        RECT -45.095 -175.525 -44.925 -175.355 ;
        RECT -44.635 -175.525 -44.465 -175.355 ;
        RECT -37.475 -175.525 -37.305 -175.355 ;
        RECT -37.015 -175.525 -36.845 -175.355 ;
        RECT -36.555 -175.525 -36.385 -175.355 ;
        RECT -36.095 -175.525 -35.925 -175.355 ;
        RECT -35.635 -175.525 -35.465 -175.355 ;
        RECT -35.175 -175.525 -35.005 -175.355 ;
        RECT -34.715 -175.525 -34.545 -175.355 ;
        RECT -27.555 -175.525 -27.385 -175.355 ;
        RECT -27.095 -175.525 -26.925 -175.355 ;
        RECT -26.635 -175.525 -26.465 -175.355 ;
        RECT -26.175 -175.525 -26.005 -175.355 ;
        RECT -25.715 -175.525 -25.545 -175.355 ;
        RECT -25.255 -175.525 -25.085 -175.355 ;
        RECT -24.795 -175.525 -24.625 -175.355 ;
        RECT -17.635 -175.525 -17.465 -175.355 ;
        RECT -17.175 -175.525 -17.005 -175.355 ;
        RECT -16.715 -175.525 -16.545 -175.355 ;
        RECT -16.255 -175.525 -16.085 -175.355 ;
        RECT -15.795 -175.525 -15.625 -175.355 ;
        RECT -15.335 -175.525 -15.165 -175.355 ;
        RECT -14.875 -175.525 -14.705 -175.355 ;
        RECT -7.715 -175.525 -7.545 -175.355 ;
        RECT -7.255 -175.525 -7.085 -175.355 ;
        RECT -6.795 -175.525 -6.625 -175.355 ;
        RECT -6.335 -175.525 -6.165 -175.355 ;
        RECT -5.875 -175.525 -5.705 -175.355 ;
        RECT -5.415 -175.525 -5.245 -175.355 ;
        RECT -4.955 -175.525 -4.785 -175.355 ;
        RECT 2.205 -175.525 2.375 -175.355 ;
        RECT 2.665 -175.525 2.835 -175.355 ;
        RECT 3.125 -175.525 3.295 -175.355 ;
        RECT 3.585 -175.525 3.755 -175.355 ;
        RECT 4.045 -175.525 4.215 -175.355 ;
        RECT 4.505 -175.525 4.675 -175.355 ;
        RECT 4.965 -175.525 5.135 -175.355 ;
        RECT 12.125 -175.525 12.295 -175.355 ;
        RECT 12.585 -175.525 12.755 -175.355 ;
        RECT 13.045 -175.525 13.215 -175.355 ;
        RECT 13.505 -175.525 13.675 -175.355 ;
        RECT 13.965 -175.525 14.135 -175.355 ;
        RECT 14.425 -175.525 14.595 -175.355 ;
        RECT 14.885 -175.525 15.055 -175.355 ;
        RECT 22.045 -175.525 22.215 -175.355 ;
        RECT 22.505 -175.525 22.675 -175.355 ;
        RECT 22.965 -175.525 23.135 -175.355 ;
        RECT 23.425 -175.525 23.595 -175.355 ;
        RECT 23.885 -175.525 24.055 -175.355 ;
        RECT 24.345 -175.525 24.515 -175.355 ;
        RECT 24.805 -175.525 24.975 -175.355 ;
        RECT -280.515 -178.245 -280.345 -178.075 ;
        RECT -280.055 -178.245 -279.885 -178.075 ;
        RECT -279.595 -178.245 -279.425 -178.075 ;
        RECT -279.135 -178.245 -278.965 -178.075 ;
        RECT -278.675 -178.245 -278.505 -178.075 ;
        RECT -278.215 -178.245 -278.045 -178.075 ;
        RECT -277.755 -178.245 -277.585 -178.075 ;
        RECT -270.595 -178.245 -270.425 -178.075 ;
        RECT -270.135 -178.245 -269.965 -178.075 ;
        RECT -269.675 -178.245 -269.505 -178.075 ;
        RECT -269.215 -178.245 -269.045 -178.075 ;
        RECT -268.755 -178.245 -268.585 -178.075 ;
        RECT -268.295 -178.245 -268.125 -178.075 ;
        RECT -267.835 -178.245 -267.665 -178.075 ;
        RECT -260.675 -178.245 -260.505 -178.075 ;
        RECT -260.215 -178.245 -260.045 -178.075 ;
        RECT -259.755 -178.245 -259.585 -178.075 ;
        RECT -259.295 -178.245 -259.125 -178.075 ;
        RECT -258.835 -178.245 -258.665 -178.075 ;
        RECT -258.375 -178.245 -258.205 -178.075 ;
        RECT -257.915 -178.245 -257.745 -178.075 ;
        RECT -250.755 -178.245 -250.585 -178.075 ;
        RECT -250.295 -178.245 -250.125 -178.075 ;
        RECT -249.835 -178.245 -249.665 -178.075 ;
        RECT -249.375 -178.245 -249.205 -178.075 ;
        RECT -248.915 -178.245 -248.745 -178.075 ;
        RECT -248.455 -178.245 -248.285 -178.075 ;
        RECT -247.995 -178.245 -247.825 -178.075 ;
        RECT -240.835 -178.245 -240.665 -178.075 ;
        RECT -240.375 -178.245 -240.205 -178.075 ;
        RECT -239.915 -178.245 -239.745 -178.075 ;
        RECT -239.455 -178.245 -239.285 -178.075 ;
        RECT -238.995 -178.245 -238.825 -178.075 ;
        RECT -238.535 -178.245 -238.365 -178.075 ;
        RECT -238.075 -178.245 -237.905 -178.075 ;
        RECT -230.915 -178.245 -230.745 -178.075 ;
        RECT -230.455 -178.245 -230.285 -178.075 ;
        RECT -229.995 -178.245 -229.825 -178.075 ;
        RECT -229.535 -178.245 -229.365 -178.075 ;
        RECT -229.075 -178.245 -228.905 -178.075 ;
        RECT -228.615 -178.245 -228.445 -178.075 ;
        RECT -228.155 -178.245 -227.985 -178.075 ;
        RECT -220.995 -178.245 -220.825 -178.075 ;
        RECT -220.535 -178.245 -220.365 -178.075 ;
        RECT -220.075 -178.245 -219.905 -178.075 ;
        RECT -219.615 -178.245 -219.445 -178.075 ;
        RECT -219.155 -178.245 -218.985 -178.075 ;
        RECT -218.695 -178.245 -218.525 -178.075 ;
        RECT -218.235 -178.245 -218.065 -178.075 ;
        RECT -211.075 -178.245 -210.905 -178.075 ;
        RECT -210.615 -178.245 -210.445 -178.075 ;
        RECT -210.155 -178.245 -209.985 -178.075 ;
        RECT -209.695 -178.245 -209.525 -178.075 ;
        RECT -209.235 -178.245 -209.065 -178.075 ;
        RECT -208.775 -178.245 -208.605 -178.075 ;
        RECT -208.315 -178.245 -208.145 -178.075 ;
        RECT -201.155 -178.245 -200.985 -178.075 ;
        RECT -200.695 -178.245 -200.525 -178.075 ;
        RECT -200.235 -178.245 -200.065 -178.075 ;
        RECT -199.775 -178.245 -199.605 -178.075 ;
        RECT -199.315 -178.245 -199.145 -178.075 ;
        RECT -198.855 -178.245 -198.685 -178.075 ;
        RECT -198.395 -178.245 -198.225 -178.075 ;
        RECT -191.235 -178.245 -191.065 -178.075 ;
        RECT -190.775 -178.245 -190.605 -178.075 ;
        RECT -190.315 -178.245 -190.145 -178.075 ;
        RECT -189.855 -178.245 -189.685 -178.075 ;
        RECT -189.395 -178.245 -189.225 -178.075 ;
        RECT -188.935 -178.245 -188.765 -178.075 ;
        RECT -188.475 -178.245 -188.305 -178.075 ;
        RECT -181.315 -178.245 -181.145 -178.075 ;
        RECT -180.855 -178.245 -180.685 -178.075 ;
        RECT -180.395 -178.245 -180.225 -178.075 ;
        RECT -179.935 -178.245 -179.765 -178.075 ;
        RECT -179.475 -178.245 -179.305 -178.075 ;
        RECT -179.015 -178.245 -178.845 -178.075 ;
        RECT -178.555 -178.245 -178.385 -178.075 ;
        RECT -171.395 -178.245 -171.225 -178.075 ;
        RECT -170.935 -178.245 -170.765 -178.075 ;
        RECT -170.475 -178.245 -170.305 -178.075 ;
        RECT -170.015 -178.245 -169.845 -178.075 ;
        RECT -169.555 -178.245 -169.385 -178.075 ;
        RECT -169.095 -178.245 -168.925 -178.075 ;
        RECT -168.635 -178.245 -168.465 -178.075 ;
        RECT -161.475 -178.245 -161.305 -178.075 ;
        RECT -161.015 -178.245 -160.845 -178.075 ;
        RECT -160.555 -178.245 -160.385 -178.075 ;
        RECT -160.095 -178.245 -159.925 -178.075 ;
        RECT -159.635 -178.245 -159.465 -178.075 ;
        RECT -159.175 -178.245 -159.005 -178.075 ;
        RECT -158.715 -178.245 -158.545 -178.075 ;
        RECT -151.555 -178.245 -151.385 -178.075 ;
        RECT -151.095 -178.245 -150.925 -178.075 ;
        RECT -150.635 -178.245 -150.465 -178.075 ;
        RECT -150.175 -178.245 -150.005 -178.075 ;
        RECT -149.715 -178.245 -149.545 -178.075 ;
        RECT -149.255 -178.245 -149.085 -178.075 ;
        RECT -148.795 -178.245 -148.625 -178.075 ;
        RECT -141.635 -178.245 -141.465 -178.075 ;
        RECT -141.175 -178.245 -141.005 -178.075 ;
        RECT -140.715 -178.245 -140.545 -178.075 ;
        RECT -140.255 -178.245 -140.085 -178.075 ;
        RECT -139.795 -178.245 -139.625 -178.075 ;
        RECT -139.335 -178.245 -139.165 -178.075 ;
        RECT -138.875 -178.245 -138.705 -178.075 ;
        RECT -131.715 -178.245 -131.545 -178.075 ;
        RECT -131.255 -178.245 -131.085 -178.075 ;
        RECT -130.795 -178.245 -130.625 -178.075 ;
        RECT -130.335 -178.245 -130.165 -178.075 ;
        RECT -129.875 -178.245 -129.705 -178.075 ;
        RECT -129.415 -178.245 -129.245 -178.075 ;
        RECT -128.955 -178.245 -128.785 -178.075 ;
        RECT -121.795 -178.245 -121.625 -178.075 ;
        RECT -121.335 -178.245 -121.165 -178.075 ;
        RECT -120.875 -178.245 -120.705 -178.075 ;
        RECT -120.415 -178.245 -120.245 -178.075 ;
        RECT -119.955 -178.245 -119.785 -178.075 ;
        RECT -119.495 -178.245 -119.325 -178.075 ;
        RECT -119.035 -178.245 -118.865 -178.075 ;
        RECT -111.875 -178.245 -111.705 -178.075 ;
        RECT -111.415 -178.245 -111.245 -178.075 ;
        RECT -110.955 -178.245 -110.785 -178.075 ;
        RECT -110.495 -178.245 -110.325 -178.075 ;
        RECT -110.035 -178.245 -109.865 -178.075 ;
        RECT -109.575 -178.245 -109.405 -178.075 ;
        RECT -109.115 -178.245 -108.945 -178.075 ;
        RECT -101.955 -178.245 -101.785 -178.075 ;
        RECT -101.495 -178.245 -101.325 -178.075 ;
        RECT -101.035 -178.245 -100.865 -178.075 ;
        RECT -100.575 -178.245 -100.405 -178.075 ;
        RECT -100.115 -178.245 -99.945 -178.075 ;
        RECT -99.655 -178.245 -99.485 -178.075 ;
        RECT -99.195 -178.245 -99.025 -178.075 ;
        RECT -92.035 -178.245 -91.865 -178.075 ;
        RECT -91.575 -178.245 -91.405 -178.075 ;
        RECT -91.115 -178.245 -90.945 -178.075 ;
        RECT -90.655 -178.245 -90.485 -178.075 ;
        RECT -90.195 -178.245 -90.025 -178.075 ;
        RECT -89.735 -178.245 -89.565 -178.075 ;
        RECT -89.275 -178.245 -89.105 -178.075 ;
        RECT -82.115 -178.245 -81.945 -178.075 ;
        RECT -81.655 -178.245 -81.485 -178.075 ;
        RECT -81.195 -178.245 -81.025 -178.075 ;
        RECT -80.735 -178.245 -80.565 -178.075 ;
        RECT -80.275 -178.245 -80.105 -178.075 ;
        RECT -79.815 -178.245 -79.645 -178.075 ;
        RECT -79.355 -178.245 -79.185 -178.075 ;
        RECT -72.195 -178.245 -72.025 -178.075 ;
        RECT -71.735 -178.245 -71.565 -178.075 ;
        RECT -71.275 -178.245 -71.105 -178.075 ;
        RECT -70.815 -178.245 -70.645 -178.075 ;
        RECT -70.355 -178.245 -70.185 -178.075 ;
        RECT -69.895 -178.245 -69.725 -178.075 ;
        RECT -69.435 -178.245 -69.265 -178.075 ;
        RECT -62.275 -178.245 -62.105 -178.075 ;
        RECT -61.815 -178.245 -61.645 -178.075 ;
        RECT -61.355 -178.245 -61.185 -178.075 ;
        RECT -60.895 -178.245 -60.725 -178.075 ;
        RECT -60.435 -178.245 -60.265 -178.075 ;
        RECT -59.975 -178.245 -59.805 -178.075 ;
        RECT -59.515 -178.245 -59.345 -178.075 ;
        RECT -52.355 -178.245 -52.185 -178.075 ;
        RECT -51.895 -178.245 -51.725 -178.075 ;
        RECT -51.435 -178.245 -51.265 -178.075 ;
        RECT -50.975 -178.245 -50.805 -178.075 ;
        RECT -50.515 -178.245 -50.345 -178.075 ;
        RECT -50.055 -178.245 -49.885 -178.075 ;
        RECT -49.595 -178.245 -49.425 -178.075 ;
        RECT -42.435 -178.245 -42.265 -178.075 ;
        RECT -41.975 -178.245 -41.805 -178.075 ;
        RECT -41.515 -178.245 -41.345 -178.075 ;
        RECT -41.055 -178.245 -40.885 -178.075 ;
        RECT -40.595 -178.245 -40.425 -178.075 ;
        RECT -40.135 -178.245 -39.965 -178.075 ;
        RECT -39.675 -178.245 -39.505 -178.075 ;
        RECT -32.515 -178.245 -32.345 -178.075 ;
        RECT -32.055 -178.245 -31.885 -178.075 ;
        RECT -31.595 -178.245 -31.425 -178.075 ;
        RECT -31.135 -178.245 -30.965 -178.075 ;
        RECT -30.675 -178.245 -30.505 -178.075 ;
        RECT -30.215 -178.245 -30.045 -178.075 ;
        RECT -29.755 -178.245 -29.585 -178.075 ;
        RECT -22.595 -178.245 -22.425 -178.075 ;
        RECT -22.135 -178.245 -21.965 -178.075 ;
        RECT -21.675 -178.245 -21.505 -178.075 ;
        RECT -21.215 -178.245 -21.045 -178.075 ;
        RECT -20.755 -178.245 -20.585 -178.075 ;
        RECT -20.295 -178.245 -20.125 -178.075 ;
        RECT -19.835 -178.245 -19.665 -178.075 ;
        RECT -12.675 -178.245 -12.505 -178.075 ;
        RECT -12.215 -178.245 -12.045 -178.075 ;
        RECT -11.755 -178.245 -11.585 -178.075 ;
        RECT -11.295 -178.245 -11.125 -178.075 ;
        RECT -10.835 -178.245 -10.665 -178.075 ;
        RECT -10.375 -178.245 -10.205 -178.075 ;
        RECT -9.915 -178.245 -9.745 -178.075 ;
        RECT -2.755 -178.245 -2.585 -178.075 ;
        RECT -2.295 -178.245 -2.125 -178.075 ;
        RECT -1.835 -178.245 -1.665 -178.075 ;
        RECT -1.375 -178.245 -1.205 -178.075 ;
        RECT -0.915 -178.245 -0.745 -178.075 ;
        RECT -0.455 -178.245 -0.285 -178.075 ;
        RECT 0.005 -178.245 0.175 -178.075 ;
        RECT 7.165 -178.245 7.335 -178.075 ;
        RECT 7.625 -178.245 7.795 -178.075 ;
        RECT 8.085 -178.245 8.255 -178.075 ;
        RECT 8.545 -178.245 8.715 -178.075 ;
        RECT 9.005 -178.245 9.175 -178.075 ;
        RECT 9.465 -178.245 9.635 -178.075 ;
        RECT 9.925 -178.245 10.095 -178.075 ;
        RECT 17.085 -178.245 17.255 -178.075 ;
        RECT 17.545 -178.245 17.715 -178.075 ;
        RECT 18.005 -178.245 18.175 -178.075 ;
        RECT 18.465 -178.245 18.635 -178.075 ;
        RECT 18.925 -178.245 19.095 -178.075 ;
        RECT 19.385 -178.245 19.555 -178.075 ;
        RECT 19.845 -178.245 20.015 -178.075 ;
        RECT 27.005 -178.245 27.175 -178.075 ;
        RECT 27.465 -178.245 27.635 -178.075 ;
        RECT 27.925 -178.245 28.095 -178.075 ;
        RECT 28.385 -178.245 28.555 -178.075 ;
        RECT -284.565 -178.905 -284.395 -178.735 ;
        RECT -284.095 -178.830 -283.925 -178.660 ;
        RECT -284.565 -179.365 -284.395 -179.195 ;
        RECT -284.565 -179.825 -284.395 -179.655 ;
        RECT -283.625 -178.905 -283.455 -178.735 ;
        RECT -274.645 -178.905 -274.475 -178.735 ;
        RECT -274.175 -178.830 -274.005 -178.660 ;
        RECT -283.625 -179.365 -283.455 -179.195 ;
        RECT -274.645 -179.365 -274.475 -179.195 ;
        RECT -283.625 -179.825 -283.455 -179.655 ;
        RECT -274.645 -179.825 -274.475 -179.655 ;
        RECT -273.705 -178.905 -273.535 -178.735 ;
        RECT -264.725 -178.905 -264.555 -178.735 ;
        RECT -264.255 -178.830 -264.085 -178.660 ;
        RECT -273.705 -179.365 -273.535 -179.195 ;
        RECT -264.725 -179.365 -264.555 -179.195 ;
        RECT -273.705 -179.825 -273.535 -179.655 ;
        RECT -264.725 -179.825 -264.555 -179.655 ;
        RECT -263.785 -178.905 -263.615 -178.735 ;
        RECT -254.805 -178.905 -254.635 -178.735 ;
        RECT -254.335 -178.830 -254.165 -178.660 ;
        RECT -263.785 -179.365 -263.615 -179.195 ;
        RECT -254.805 -179.365 -254.635 -179.195 ;
        RECT -263.785 -179.825 -263.615 -179.655 ;
        RECT -254.805 -179.825 -254.635 -179.655 ;
        RECT -253.865 -178.905 -253.695 -178.735 ;
        RECT -244.885 -178.905 -244.715 -178.735 ;
        RECT -244.415 -178.830 -244.245 -178.660 ;
        RECT -253.865 -179.365 -253.695 -179.195 ;
        RECT -244.885 -179.365 -244.715 -179.195 ;
        RECT -253.865 -179.825 -253.695 -179.655 ;
        RECT -244.885 -179.825 -244.715 -179.655 ;
        RECT -243.945 -178.905 -243.775 -178.735 ;
        RECT -234.965 -178.905 -234.795 -178.735 ;
        RECT -234.495 -178.830 -234.325 -178.660 ;
        RECT -243.945 -179.365 -243.775 -179.195 ;
        RECT -234.965 -179.365 -234.795 -179.195 ;
        RECT -243.945 -179.825 -243.775 -179.655 ;
        RECT -234.965 -179.825 -234.795 -179.655 ;
        RECT -234.025 -178.905 -233.855 -178.735 ;
        RECT -225.045 -178.905 -224.875 -178.735 ;
        RECT -224.575 -178.830 -224.405 -178.660 ;
        RECT -234.025 -179.365 -233.855 -179.195 ;
        RECT -225.045 -179.365 -224.875 -179.195 ;
        RECT -234.025 -179.825 -233.855 -179.655 ;
        RECT -225.045 -179.825 -224.875 -179.655 ;
        RECT -224.105 -178.905 -223.935 -178.735 ;
        RECT -215.125 -178.905 -214.955 -178.735 ;
        RECT -214.655 -178.830 -214.485 -178.660 ;
        RECT -224.105 -179.365 -223.935 -179.195 ;
        RECT -215.125 -179.365 -214.955 -179.195 ;
        RECT -224.105 -179.825 -223.935 -179.655 ;
        RECT -215.125 -179.825 -214.955 -179.655 ;
        RECT -214.185 -178.905 -214.015 -178.735 ;
        RECT -205.205 -178.905 -205.035 -178.735 ;
        RECT -204.735 -178.830 -204.565 -178.660 ;
        RECT -214.185 -179.365 -214.015 -179.195 ;
        RECT -205.205 -179.365 -205.035 -179.195 ;
        RECT -214.185 -179.825 -214.015 -179.655 ;
        RECT -205.205 -179.825 -205.035 -179.655 ;
        RECT -204.265 -178.905 -204.095 -178.735 ;
        RECT -195.285 -178.905 -195.115 -178.735 ;
        RECT -194.815 -178.830 -194.645 -178.660 ;
        RECT -204.265 -179.365 -204.095 -179.195 ;
        RECT -195.285 -179.365 -195.115 -179.195 ;
        RECT -204.265 -179.825 -204.095 -179.655 ;
        RECT -195.285 -179.825 -195.115 -179.655 ;
        RECT -194.345 -178.905 -194.175 -178.735 ;
        RECT -185.365 -178.905 -185.195 -178.735 ;
        RECT -184.895 -178.830 -184.725 -178.660 ;
        RECT -194.345 -179.365 -194.175 -179.195 ;
        RECT -185.365 -179.365 -185.195 -179.195 ;
        RECT -194.345 -179.825 -194.175 -179.655 ;
        RECT -185.365 -179.825 -185.195 -179.655 ;
        RECT -184.425 -178.905 -184.255 -178.735 ;
        RECT -175.445 -178.905 -175.275 -178.735 ;
        RECT -174.975 -178.830 -174.805 -178.660 ;
        RECT -184.425 -179.365 -184.255 -179.195 ;
        RECT -175.445 -179.365 -175.275 -179.195 ;
        RECT -184.425 -179.825 -184.255 -179.655 ;
        RECT -175.445 -179.825 -175.275 -179.655 ;
        RECT -174.505 -178.905 -174.335 -178.735 ;
        RECT -165.525 -178.905 -165.355 -178.735 ;
        RECT -165.055 -178.830 -164.885 -178.660 ;
        RECT -174.505 -179.365 -174.335 -179.195 ;
        RECT -165.525 -179.365 -165.355 -179.195 ;
        RECT -174.505 -179.825 -174.335 -179.655 ;
        RECT -165.525 -179.825 -165.355 -179.655 ;
        RECT -164.585 -178.905 -164.415 -178.735 ;
        RECT -155.605 -178.905 -155.435 -178.735 ;
        RECT -155.135 -178.830 -154.965 -178.660 ;
        RECT -164.585 -179.365 -164.415 -179.195 ;
        RECT -155.605 -179.365 -155.435 -179.195 ;
        RECT -164.585 -179.825 -164.415 -179.655 ;
        RECT -155.605 -179.825 -155.435 -179.655 ;
        RECT -154.665 -178.905 -154.495 -178.735 ;
        RECT -145.685 -178.905 -145.515 -178.735 ;
        RECT -145.215 -178.830 -145.045 -178.660 ;
        RECT -154.665 -179.365 -154.495 -179.195 ;
        RECT -145.685 -179.365 -145.515 -179.195 ;
        RECT -154.665 -179.825 -154.495 -179.655 ;
        RECT -145.685 -179.825 -145.515 -179.655 ;
        RECT -144.745 -178.905 -144.575 -178.735 ;
        RECT -135.765 -178.905 -135.595 -178.735 ;
        RECT -135.295 -178.830 -135.125 -178.660 ;
        RECT -144.745 -179.365 -144.575 -179.195 ;
        RECT -135.765 -179.365 -135.595 -179.195 ;
        RECT -144.745 -179.825 -144.575 -179.655 ;
        RECT -135.765 -179.825 -135.595 -179.655 ;
        RECT -134.825 -178.905 -134.655 -178.735 ;
        RECT -125.845 -178.905 -125.675 -178.735 ;
        RECT -125.375 -178.830 -125.205 -178.660 ;
        RECT -134.825 -179.365 -134.655 -179.195 ;
        RECT -125.845 -179.365 -125.675 -179.195 ;
        RECT -134.825 -179.825 -134.655 -179.655 ;
        RECT -125.845 -179.825 -125.675 -179.655 ;
        RECT -124.905 -178.905 -124.735 -178.735 ;
        RECT -115.925 -178.905 -115.755 -178.735 ;
        RECT -115.455 -178.830 -115.285 -178.660 ;
        RECT -124.905 -179.365 -124.735 -179.195 ;
        RECT -115.925 -179.365 -115.755 -179.195 ;
        RECT -124.905 -179.825 -124.735 -179.655 ;
        RECT -115.925 -179.825 -115.755 -179.655 ;
        RECT -114.985 -178.905 -114.815 -178.735 ;
        RECT -106.005 -178.905 -105.835 -178.735 ;
        RECT -105.535 -178.830 -105.365 -178.660 ;
        RECT -114.985 -179.365 -114.815 -179.195 ;
        RECT -106.005 -179.365 -105.835 -179.195 ;
        RECT -114.985 -179.825 -114.815 -179.655 ;
        RECT -106.005 -179.825 -105.835 -179.655 ;
        RECT -105.065 -178.905 -104.895 -178.735 ;
        RECT -96.085 -178.905 -95.915 -178.735 ;
        RECT -95.615 -178.830 -95.445 -178.660 ;
        RECT -105.065 -179.365 -104.895 -179.195 ;
        RECT -96.085 -179.365 -95.915 -179.195 ;
        RECT -105.065 -179.825 -104.895 -179.655 ;
        RECT -96.085 -179.825 -95.915 -179.655 ;
        RECT -95.145 -178.905 -94.975 -178.735 ;
        RECT -86.165 -178.905 -85.995 -178.735 ;
        RECT -85.695 -178.830 -85.525 -178.660 ;
        RECT -95.145 -179.365 -94.975 -179.195 ;
        RECT -86.165 -179.365 -85.995 -179.195 ;
        RECT -95.145 -179.825 -94.975 -179.655 ;
        RECT -86.165 -179.825 -85.995 -179.655 ;
        RECT -85.225 -178.905 -85.055 -178.735 ;
        RECT -76.245 -178.905 -76.075 -178.735 ;
        RECT -75.775 -178.830 -75.605 -178.660 ;
        RECT -85.225 -179.365 -85.055 -179.195 ;
        RECT -76.245 -179.365 -76.075 -179.195 ;
        RECT -85.225 -179.825 -85.055 -179.655 ;
        RECT -76.245 -179.825 -76.075 -179.655 ;
        RECT -75.305 -178.905 -75.135 -178.735 ;
        RECT -66.325 -178.905 -66.155 -178.735 ;
        RECT -65.855 -178.830 -65.685 -178.660 ;
        RECT -75.305 -179.365 -75.135 -179.195 ;
        RECT -66.325 -179.365 -66.155 -179.195 ;
        RECT -75.305 -179.825 -75.135 -179.655 ;
        RECT -66.325 -179.825 -66.155 -179.655 ;
        RECT -65.385 -178.905 -65.215 -178.735 ;
        RECT -56.405 -178.905 -56.235 -178.735 ;
        RECT -55.935 -178.830 -55.765 -178.660 ;
        RECT -65.385 -179.365 -65.215 -179.195 ;
        RECT -56.405 -179.365 -56.235 -179.195 ;
        RECT -65.385 -179.825 -65.215 -179.655 ;
        RECT -56.405 -179.825 -56.235 -179.655 ;
        RECT -55.465 -178.905 -55.295 -178.735 ;
        RECT -46.485 -178.905 -46.315 -178.735 ;
        RECT -46.015 -178.830 -45.845 -178.660 ;
        RECT -55.465 -179.365 -55.295 -179.195 ;
        RECT -46.485 -179.365 -46.315 -179.195 ;
        RECT -55.465 -179.825 -55.295 -179.655 ;
        RECT -46.485 -179.825 -46.315 -179.655 ;
        RECT -45.545 -178.905 -45.375 -178.735 ;
        RECT -36.565 -178.905 -36.395 -178.735 ;
        RECT -36.095 -178.830 -35.925 -178.660 ;
        RECT -45.545 -179.365 -45.375 -179.195 ;
        RECT -36.565 -179.365 -36.395 -179.195 ;
        RECT -45.545 -179.825 -45.375 -179.655 ;
        RECT -36.565 -179.825 -36.395 -179.655 ;
        RECT -35.625 -178.905 -35.455 -178.735 ;
        RECT -26.645 -178.905 -26.475 -178.735 ;
        RECT -26.175 -178.830 -26.005 -178.660 ;
        RECT -35.625 -179.365 -35.455 -179.195 ;
        RECT -26.645 -179.365 -26.475 -179.195 ;
        RECT -35.625 -179.825 -35.455 -179.655 ;
        RECT -26.645 -179.825 -26.475 -179.655 ;
        RECT -25.705 -178.905 -25.535 -178.735 ;
        RECT -16.725 -178.905 -16.555 -178.735 ;
        RECT -16.255 -178.830 -16.085 -178.660 ;
        RECT -25.705 -179.365 -25.535 -179.195 ;
        RECT -16.725 -179.365 -16.555 -179.195 ;
        RECT -25.705 -179.825 -25.535 -179.655 ;
        RECT -16.725 -179.825 -16.555 -179.655 ;
        RECT -15.785 -178.905 -15.615 -178.735 ;
        RECT -6.805 -178.905 -6.635 -178.735 ;
        RECT -6.335 -178.830 -6.165 -178.660 ;
        RECT -15.785 -179.365 -15.615 -179.195 ;
        RECT -6.805 -179.365 -6.635 -179.195 ;
        RECT -15.785 -179.825 -15.615 -179.655 ;
        RECT -6.805 -179.825 -6.635 -179.655 ;
        RECT -5.865 -178.905 -5.695 -178.735 ;
        RECT 3.115 -178.905 3.285 -178.735 ;
        RECT 3.585 -178.830 3.755 -178.660 ;
        RECT -5.865 -179.365 -5.695 -179.195 ;
        RECT 3.115 -179.365 3.285 -179.195 ;
        RECT -5.865 -179.825 -5.695 -179.655 ;
        RECT 3.115 -179.825 3.285 -179.655 ;
        RECT 4.055 -178.905 4.225 -178.735 ;
        RECT 13.035 -178.905 13.205 -178.735 ;
        RECT 13.505 -178.830 13.675 -178.660 ;
        RECT 4.055 -179.365 4.225 -179.195 ;
        RECT 13.035 -179.365 13.205 -179.195 ;
        RECT 4.055 -179.825 4.225 -179.655 ;
        RECT 13.035 -179.825 13.205 -179.655 ;
        RECT 13.975 -178.905 14.145 -178.735 ;
        RECT 22.955 -178.905 23.125 -178.735 ;
        RECT 23.425 -178.830 23.595 -178.660 ;
        RECT 13.975 -179.365 14.145 -179.195 ;
        RECT 22.955 -179.365 23.125 -179.195 ;
        RECT 13.975 -179.825 14.145 -179.655 ;
        RECT 22.955 -179.825 23.125 -179.655 ;
        RECT 23.895 -178.905 24.065 -178.735 ;
        RECT 23.895 -179.365 24.065 -179.195 ;
        RECT 23.895 -179.825 24.065 -179.655 ;
      LAYER met1 ;
        RECT -281.540 95.140 -281.080 95.145 ;
        RECT -271.620 95.140 -271.160 95.145 ;
        RECT -261.700 95.140 -261.240 95.145 ;
        RECT -251.780 95.140 -251.320 95.145 ;
        RECT -241.860 95.140 -241.400 95.145 ;
        RECT -231.940 95.140 -231.480 95.145 ;
        RECT -222.020 95.140 -221.560 95.145 ;
        RECT -212.100 95.140 -211.640 95.145 ;
        RECT -202.180 95.140 -201.720 95.145 ;
        RECT -192.260 95.140 -191.800 95.145 ;
        RECT -182.340 95.140 -181.880 95.145 ;
        RECT -172.420 95.140 -171.960 95.145 ;
        RECT -162.500 95.140 -162.040 95.145 ;
        RECT -152.580 95.140 -152.120 95.145 ;
        RECT -142.660 95.140 -142.200 95.145 ;
        RECT -132.740 95.140 -132.280 95.145 ;
        RECT -122.820 95.140 -122.360 95.145 ;
        RECT -112.900 95.140 -112.440 95.145 ;
        RECT -102.980 95.140 -102.520 95.145 ;
        RECT -93.060 95.140 -92.600 95.145 ;
        RECT -83.140 95.140 -82.680 95.145 ;
        RECT -73.220 95.140 -72.760 95.145 ;
        RECT -63.300 95.140 -62.840 95.145 ;
        RECT -53.380 95.140 -52.920 95.145 ;
        RECT -43.460 95.140 -43.000 95.145 ;
        RECT -33.540 95.140 -33.080 95.145 ;
        RECT -23.620 95.140 -23.160 95.145 ;
        RECT -13.700 95.140 -13.240 95.145 ;
        RECT -3.780 95.140 -3.320 95.145 ;
        RECT 6.140 95.140 6.600 95.145 ;
        RECT 16.060 95.140 16.520 95.145 ;
        RECT 25.980 95.140 26.440 95.145 ;
        RECT -282.020 93.760 -280.600 95.140 ;
        RECT -272.100 93.760 -270.680 95.140 ;
        RECT -262.180 93.760 -260.760 95.140 ;
        RECT -252.260 93.760 -250.840 95.140 ;
        RECT -242.340 93.760 -240.920 95.140 ;
        RECT -232.420 93.760 -231.000 95.140 ;
        RECT -222.500 93.760 -221.080 95.140 ;
        RECT -212.580 93.760 -211.160 95.140 ;
        RECT -202.660 93.760 -201.240 95.140 ;
        RECT -192.740 93.760 -191.320 95.140 ;
        RECT -182.820 93.760 -181.400 95.140 ;
        RECT -172.900 93.760 -171.480 95.140 ;
        RECT -162.980 93.760 -161.560 95.140 ;
        RECT -153.060 93.760 -151.640 95.140 ;
        RECT -143.140 93.760 -141.720 95.140 ;
        RECT -133.220 93.760 -131.800 95.140 ;
        RECT -123.300 93.760 -121.880 95.140 ;
        RECT -113.380 93.760 -111.960 95.140 ;
        RECT -103.460 93.760 -102.040 95.140 ;
        RECT -93.540 93.760 -92.120 95.140 ;
        RECT -83.620 93.760 -82.200 95.140 ;
        RECT -73.700 93.760 -72.280 95.140 ;
        RECT -63.780 93.760 -62.360 95.140 ;
        RECT -53.860 93.760 -52.440 95.140 ;
        RECT -43.940 93.760 -42.520 95.140 ;
        RECT -34.020 93.760 -32.600 95.140 ;
        RECT -24.100 93.760 -22.680 95.140 ;
        RECT -14.180 93.760 -12.760 95.140 ;
        RECT -4.260 93.760 -2.840 95.140 ;
        RECT 5.660 93.760 7.080 95.140 ;
        RECT 15.580 93.760 17.000 95.140 ;
        RECT 25.500 93.760 26.440 95.140 ;
        RECT -287.880 93.090 -284.660 93.570 ;
        RECT -277.960 93.090 -274.740 93.570 ;
        RECT -268.040 93.090 -264.820 93.570 ;
        RECT -258.120 93.090 -254.900 93.570 ;
        RECT -248.200 93.090 -244.980 93.570 ;
        RECT -238.280 93.090 -235.060 93.570 ;
        RECT -228.360 93.090 -225.140 93.570 ;
        RECT -218.440 93.090 -215.220 93.570 ;
        RECT -208.520 93.090 -205.300 93.570 ;
        RECT -198.600 93.090 -195.380 93.570 ;
        RECT -188.680 93.090 -185.460 93.570 ;
        RECT -178.760 93.090 -175.540 93.570 ;
        RECT -168.840 93.090 -165.620 93.570 ;
        RECT -158.920 93.090 -155.700 93.570 ;
        RECT -149.000 93.090 -145.780 93.570 ;
        RECT -139.080 93.090 -135.860 93.570 ;
        RECT -129.160 93.090 -125.940 93.570 ;
        RECT -119.240 93.090 -116.020 93.570 ;
        RECT -109.320 93.090 -106.100 93.570 ;
        RECT -99.400 93.090 -96.180 93.570 ;
        RECT -89.480 93.090 -86.260 93.570 ;
        RECT -79.560 93.090 -76.340 93.570 ;
        RECT -69.640 93.090 -66.420 93.570 ;
        RECT -59.720 93.090 -56.500 93.570 ;
        RECT -49.800 93.090 -46.580 93.570 ;
        RECT -39.880 93.090 -36.660 93.570 ;
        RECT -29.960 93.090 -26.740 93.570 ;
        RECT -20.040 93.090 -16.820 93.570 ;
        RECT -10.120 93.090 -6.900 93.570 ;
        RECT -0.200 93.090 3.020 93.570 ;
        RECT 9.720 93.090 12.940 93.570 ;
        RECT 19.640 93.090 22.860 93.570 ;
        RECT -282.920 90.370 -279.700 90.850 ;
        RECT -273.000 90.370 -269.780 90.850 ;
        RECT -263.080 90.370 -259.860 90.850 ;
        RECT -253.160 90.370 -249.940 90.850 ;
        RECT -243.240 90.370 -240.020 90.850 ;
        RECT -233.320 90.370 -230.100 90.850 ;
        RECT -223.400 90.370 -220.180 90.850 ;
        RECT -213.480 90.370 -210.260 90.850 ;
        RECT -203.560 90.370 -200.340 90.850 ;
        RECT -193.640 90.370 -190.420 90.850 ;
        RECT -183.720 90.370 -180.500 90.850 ;
        RECT -173.800 90.370 -170.580 90.850 ;
        RECT -163.880 90.370 -160.660 90.850 ;
        RECT -153.960 90.370 -150.740 90.850 ;
        RECT -144.040 90.370 -140.820 90.850 ;
        RECT -134.120 90.370 -130.900 90.850 ;
        RECT -124.200 90.370 -120.980 90.850 ;
        RECT -114.280 90.370 -111.060 90.850 ;
        RECT -104.360 90.370 -101.140 90.850 ;
        RECT -94.440 90.370 -91.220 90.850 ;
        RECT -84.520 90.370 -81.300 90.850 ;
        RECT -74.600 90.370 -71.380 90.850 ;
        RECT -64.680 90.370 -61.460 90.850 ;
        RECT -54.760 90.370 -51.540 90.850 ;
        RECT -44.840 90.370 -41.620 90.850 ;
        RECT -34.920 90.370 -31.700 90.850 ;
        RECT -25.000 90.370 -21.780 90.850 ;
        RECT -15.080 90.370 -11.860 90.850 ;
        RECT -5.160 90.370 -1.940 90.850 ;
        RECT 4.760 90.370 7.980 90.850 ;
        RECT 14.680 90.370 17.900 90.850 ;
        RECT 24.600 90.370 26.440 90.850 ;
        RECT -222.030 90.360 -220.180 90.370 ;
        RECT -142.670 90.360 -140.820 90.370 ;
        RECT -63.310 90.360 -61.460 90.370 ;
        RECT 16.050 90.360 17.900 90.370 ;
        RECT -286.980 88.800 -285.560 90.180 ;
        RECT -277.060 88.800 -275.640 90.180 ;
        RECT -267.140 88.800 -265.720 90.180 ;
        RECT -257.220 88.800 -255.800 90.180 ;
        RECT -247.300 88.800 -245.880 90.180 ;
        RECT -237.380 88.800 -235.960 90.180 ;
        RECT -227.460 88.800 -226.040 90.180 ;
        RECT -217.540 88.800 -216.120 90.180 ;
        RECT -207.620 88.800 -206.200 90.180 ;
        RECT -197.700 88.800 -196.280 90.180 ;
        RECT -187.780 88.800 -186.360 90.180 ;
        RECT -177.860 88.800 -176.440 90.180 ;
        RECT -167.940 88.800 -166.520 90.180 ;
        RECT -158.020 88.800 -156.600 90.180 ;
        RECT -148.100 88.800 -146.680 90.180 ;
        RECT -138.180 88.800 -136.760 90.180 ;
        RECT -128.260 88.800 -126.840 90.180 ;
        RECT -118.340 88.800 -116.920 90.180 ;
        RECT -108.420 88.800 -107.000 90.180 ;
        RECT -98.500 88.800 -97.080 90.180 ;
        RECT -88.580 88.800 -87.160 90.180 ;
        RECT -78.660 88.800 -77.240 90.180 ;
        RECT -68.740 88.800 -67.320 90.180 ;
        RECT -58.820 88.800 -57.400 90.180 ;
        RECT -48.900 88.800 -47.480 90.180 ;
        RECT -38.980 88.800 -37.560 90.180 ;
        RECT -29.060 88.800 -27.640 90.180 ;
        RECT -19.140 88.800 -17.720 90.180 ;
        RECT -9.220 88.800 -7.800 90.180 ;
        RECT 0.700 88.800 2.120 90.180 ;
        RECT 10.620 88.800 12.040 90.180 ;
        RECT 20.540 88.800 21.960 90.180 ;
        RECT -281.290 7.430 -280.830 7.435 ;
        RECT -271.370 7.430 -270.910 7.435 ;
        RECT -261.450 7.430 -260.990 7.435 ;
        RECT -251.530 7.430 -251.070 7.435 ;
        RECT -241.610 7.430 -241.150 7.435 ;
        RECT -231.690 7.430 -231.230 7.435 ;
        RECT -221.770 7.430 -221.310 7.435 ;
        RECT -211.850 7.430 -211.390 7.435 ;
        RECT -201.930 7.430 -201.470 7.435 ;
        RECT -192.010 7.430 -191.550 7.435 ;
        RECT -182.090 7.430 -181.630 7.435 ;
        RECT -172.170 7.430 -171.710 7.435 ;
        RECT -162.250 7.430 -161.790 7.435 ;
        RECT -152.330 7.430 -151.870 7.435 ;
        RECT -142.410 7.430 -141.950 7.435 ;
        RECT -132.490 7.430 -132.030 7.435 ;
        RECT -122.570 7.430 -122.110 7.435 ;
        RECT -112.650 7.430 -112.190 7.435 ;
        RECT -102.730 7.430 -102.270 7.435 ;
        RECT -92.810 7.430 -92.350 7.435 ;
        RECT -82.890 7.430 -82.430 7.435 ;
        RECT -72.970 7.430 -72.510 7.435 ;
        RECT -63.050 7.430 -62.590 7.435 ;
        RECT -53.130 7.430 -52.670 7.435 ;
        RECT -43.210 7.430 -42.750 7.435 ;
        RECT -33.290 7.430 -32.830 7.435 ;
        RECT -23.370 7.430 -22.910 7.435 ;
        RECT -13.450 7.430 -12.990 7.435 ;
        RECT -3.530 7.430 -3.070 7.435 ;
        RECT 6.390 7.430 6.850 7.435 ;
        RECT 16.310 7.430 16.770 7.435 ;
        RECT 26.230 7.430 26.690 7.435 ;
        RECT -281.770 6.050 -280.350 7.430 ;
        RECT -271.850 6.050 -270.430 7.430 ;
        RECT -261.930 6.050 -260.510 7.430 ;
        RECT -252.010 6.050 -250.590 7.430 ;
        RECT -242.090 6.050 -240.670 7.430 ;
        RECT -232.170 6.050 -230.750 7.430 ;
        RECT -222.250 6.050 -220.830 7.430 ;
        RECT -212.330 6.050 -210.910 7.430 ;
        RECT -202.410 6.050 -200.990 7.430 ;
        RECT -192.490 6.050 -191.070 7.430 ;
        RECT -182.570 6.050 -181.150 7.430 ;
        RECT -172.650 6.050 -171.230 7.430 ;
        RECT -162.730 6.050 -161.310 7.430 ;
        RECT -152.810 6.050 -151.390 7.430 ;
        RECT -142.890 6.050 -141.470 7.430 ;
        RECT -132.970 6.050 -131.550 7.430 ;
        RECT -123.050 6.050 -121.630 7.430 ;
        RECT -113.130 6.050 -111.710 7.430 ;
        RECT -103.210 6.050 -101.790 7.430 ;
        RECT -93.290 6.050 -91.870 7.430 ;
        RECT -83.370 6.050 -81.950 7.430 ;
        RECT -73.450 6.050 -72.030 7.430 ;
        RECT -63.530 6.050 -62.110 7.430 ;
        RECT -53.610 6.050 -52.190 7.430 ;
        RECT -43.690 6.050 -42.270 7.430 ;
        RECT -33.770 6.050 -32.350 7.430 ;
        RECT -23.850 6.050 -22.430 7.430 ;
        RECT -13.930 6.050 -12.510 7.430 ;
        RECT -4.010 6.050 -2.590 7.430 ;
        RECT 5.910 6.050 7.330 7.430 ;
        RECT 15.830 6.050 17.250 7.430 ;
        RECT 25.750 6.050 26.690 7.430 ;
        RECT -287.630 5.380 -284.410 5.860 ;
        RECT -277.710 5.380 -274.490 5.860 ;
        RECT -267.790 5.380 -264.570 5.860 ;
        RECT -257.870 5.380 -254.650 5.860 ;
        RECT -247.950 5.380 -244.730 5.860 ;
        RECT -238.030 5.380 -234.810 5.860 ;
        RECT -228.110 5.380 -224.890 5.860 ;
        RECT -218.190 5.380 -214.970 5.860 ;
        RECT -208.270 5.380 -205.050 5.860 ;
        RECT -198.350 5.380 -195.130 5.860 ;
        RECT -188.430 5.380 -185.210 5.860 ;
        RECT -178.510 5.380 -175.290 5.860 ;
        RECT -168.590 5.380 -165.370 5.860 ;
        RECT -158.670 5.380 -155.450 5.860 ;
        RECT -148.750 5.380 -145.530 5.860 ;
        RECT -138.830 5.380 -135.610 5.860 ;
        RECT -128.910 5.380 -125.690 5.860 ;
        RECT -118.990 5.380 -115.770 5.860 ;
        RECT -109.070 5.380 -105.850 5.860 ;
        RECT -99.150 5.380 -95.930 5.860 ;
        RECT -89.230 5.380 -86.010 5.860 ;
        RECT -79.310 5.380 -76.090 5.860 ;
        RECT -69.390 5.380 -66.170 5.860 ;
        RECT -59.470 5.380 -56.250 5.860 ;
        RECT -49.550 5.380 -46.330 5.860 ;
        RECT -39.630 5.380 -36.410 5.860 ;
        RECT -29.710 5.380 -26.490 5.860 ;
        RECT -19.790 5.380 -16.570 5.860 ;
        RECT -9.870 5.380 -6.650 5.860 ;
        RECT 0.050 5.380 3.270 5.860 ;
        RECT 9.970 5.380 13.190 5.860 ;
        RECT 19.890 5.380 23.110 5.860 ;
        RECT -282.670 2.660 -279.450 3.140 ;
        RECT -272.750 2.660 -269.530 3.140 ;
        RECT -262.830 2.660 -259.610 3.140 ;
        RECT -252.910 2.660 -249.690 3.140 ;
        RECT -242.990 2.660 -239.770 3.140 ;
        RECT -233.070 2.660 -229.850 3.140 ;
        RECT -223.150 2.660 -219.930 3.140 ;
        RECT -213.230 2.660 -210.010 3.140 ;
        RECT -203.310 2.660 -200.090 3.140 ;
        RECT -193.390 2.660 -190.170 3.140 ;
        RECT -183.470 2.660 -180.250 3.140 ;
        RECT -173.550 2.660 -170.330 3.140 ;
        RECT -163.630 2.660 -160.410 3.140 ;
        RECT -153.710 2.660 -150.490 3.140 ;
        RECT -143.790 2.660 -140.570 3.140 ;
        RECT -133.870 2.660 -130.650 3.140 ;
        RECT -123.950 2.660 -120.730 3.140 ;
        RECT -114.030 2.660 -110.810 3.140 ;
        RECT -104.110 2.660 -100.890 3.140 ;
        RECT -94.190 2.660 -90.970 3.140 ;
        RECT -84.270 2.660 -81.050 3.140 ;
        RECT -74.350 2.660 -71.130 3.140 ;
        RECT -64.430 2.660 -61.210 3.140 ;
        RECT -54.510 2.660 -51.290 3.140 ;
        RECT -44.590 2.660 -41.370 3.140 ;
        RECT -34.670 2.660 -31.450 3.140 ;
        RECT -24.750 2.660 -21.530 3.140 ;
        RECT -14.830 2.660 -11.610 3.140 ;
        RECT -4.910 2.660 -1.690 3.140 ;
        RECT 5.010 2.660 8.230 3.140 ;
        RECT 14.930 2.660 18.150 3.140 ;
        RECT 24.850 2.660 26.690 3.140 ;
        RECT -221.780 2.650 -219.930 2.660 ;
        RECT -142.420 2.650 -140.570 2.660 ;
        RECT -63.060 2.650 -61.210 2.660 ;
        RECT 16.300 2.650 18.150 2.660 ;
        RECT -286.730 1.090 -285.310 2.470 ;
        RECT -276.810 1.090 -275.390 2.470 ;
        RECT -266.890 1.090 -265.470 2.470 ;
        RECT -256.970 1.090 -255.550 2.470 ;
        RECT -247.050 1.090 -245.630 2.470 ;
        RECT -237.130 1.090 -235.710 2.470 ;
        RECT -227.210 1.090 -225.790 2.470 ;
        RECT -217.290 1.090 -215.870 2.470 ;
        RECT -207.370 1.090 -205.950 2.470 ;
        RECT -197.450 1.090 -196.030 2.470 ;
        RECT -187.530 1.090 -186.110 2.470 ;
        RECT -177.610 1.090 -176.190 2.470 ;
        RECT -167.690 1.090 -166.270 2.470 ;
        RECT -157.770 1.090 -156.350 2.470 ;
        RECT -147.850 1.090 -146.430 2.470 ;
        RECT -137.930 1.090 -136.510 2.470 ;
        RECT -128.010 1.090 -126.590 2.470 ;
        RECT -118.090 1.090 -116.670 2.470 ;
        RECT -108.170 1.090 -106.750 2.470 ;
        RECT -98.250 1.090 -96.830 2.470 ;
        RECT -88.330 1.090 -86.910 2.470 ;
        RECT -78.410 1.090 -76.990 2.470 ;
        RECT -68.490 1.090 -67.070 2.470 ;
        RECT -58.570 1.090 -57.150 2.470 ;
        RECT -48.650 1.090 -47.230 2.470 ;
        RECT -38.730 1.090 -37.310 2.470 ;
        RECT -28.810 1.090 -27.390 2.470 ;
        RECT -18.890 1.090 -17.470 2.470 ;
        RECT -8.970 1.090 -7.550 2.470 ;
        RECT 0.950 1.090 2.370 2.470 ;
        RECT 10.870 1.090 12.290 2.470 ;
        RECT 20.790 1.090 22.210 2.470 ;
        RECT -279.530 -85.920 -279.070 -85.915 ;
        RECT -269.610 -85.920 -269.150 -85.915 ;
        RECT -259.690 -85.920 -259.230 -85.915 ;
        RECT -249.770 -85.920 -249.310 -85.915 ;
        RECT -239.850 -85.920 -239.390 -85.915 ;
        RECT -229.930 -85.920 -229.470 -85.915 ;
        RECT -220.010 -85.920 -219.550 -85.915 ;
        RECT -210.090 -85.920 -209.630 -85.915 ;
        RECT -200.170 -85.920 -199.710 -85.915 ;
        RECT -190.250 -85.920 -189.790 -85.915 ;
        RECT -180.330 -85.920 -179.870 -85.915 ;
        RECT -170.410 -85.920 -169.950 -85.915 ;
        RECT -160.490 -85.920 -160.030 -85.915 ;
        RECT -150.570 -85.920 -150.110 -85.915 ;
        RECT -140.650 -85.920 -140.190 -85.915 ;
        RECT -130.730 -85.920 -130.270 -85.915 ;
        RECT -120.810 -85.920 -120.350 -85.915 ;
        RECT -110.890 -85.920 -110.430 -85.915 ;
        RECT -100.970 -85.920 -100.510 -85.915 ;
        RECT -91.050 -85.920 -90.590 -85.915 ;
        RECT -81.130 -85.920 -80.670 -85.915 ;
        RECT -71.210 -85.920 -70.750 -85.915 ;
        RECT -61.290 -85.920 -60.830 -85.915 ;
        RECT -51.370 -85.920 -50.910 -85.915 ;
        RECT -41.450 -85.920 -40.990 -85.915 ;
        RECT -31.530 -85.920 -31.070 -85.915 ;
        RECT -21.610 -85.920 -21.150 -85.915 ;
        RECT -11.690 -85.920 -11.230 -85.915 ;
        RECT -1.770 -85.920 -1.310 -85.915 ;
        RECT 8.150 -85.920 8.610 -85.915 ;
        RECT 18.070 -85.920 18.530 -85.915 ;
        RECT 27.990 -85.920 28.450 -85.915 ;
        RECT -280.010 -87.300 -278.590 -85.920 ;
        RECT -270.090 -87.300 -268.670 -85.920 ;
        RECT -260.170 -87.300 -258.750 -85.920 ;
        RECT -250.250 -87.300 -248.830 -85.920 ;
        RECT -240.330 -87.300 -238.910 -85.920 ;
        RECT -230.410 -87.300 -228.990 -85.920 ;
        RECT -220.490 -87.300 -219.070 -85.920 ;
        RECT -210.570 -87.300 -209.150 -85.920 ;
        RECT -200.650 -87.300 -199.230 -85.920 ;
        RECT -190.730 -87.300 -189.310 -85.920 ;
        RECT -180.810 -87.300 -179.390 -85.920 ;
        RECT -170.890 -87.300 -169.470 -85.920 ;
        RECT -160.970 -87.300 -159.550 -85.920 ;
        RECT -151.050 -87.300 -149.630 -85.920 ;
        RECT -141.130 -87.300 -139.710 -85.920 ;
        RECT -131.210 -87.300 -129.790 -85.920 ;
        RECT -121.290 -87.300 -119.870 -85.920 ;
        RECT -111.370 -87.300 -109.950 -85.920 ;
        RECT -101.450 -87.300 -100.030 -85.920 ;
        RECT -91.530 -87.300 -90.110 -85.920 ;
        RECT -81.610 -87.300 -80.190 -85.920 ;
        RECT -71.690 -87.300 -70.270 -85.920 ;
        RECT -61.770 -87.300 -60.350 -85.920 ;
        RECT -51.850 -87.300 -50.430 -85.920 ;
        RECT -41.930 -87.300 -40.510 -85.920 ;
        RECT -32.010 -87.300 -30.590 -85.920 ;
        RECT -22.090 -87.300 -20.670 -85.920 ;
        RECT -12.170 -87.300 -10.750 -85.920 ;
        RECT -2.250 -87.300 -0.830 -85.920 ;
        RECT 7.670 -87.300 9.090 -85.920 ;
        RECT 17.590 -87.300 19.010 -85.920 ;
        RECT 27.510 -87.300 28.450 -85.920 ;
        RECT -285.870 -87.970 -282.650 -87.490 ;
        RECT -275.950 -87.970 -272.730 -87.490 ;
        RECT -266.030 -87.970 -262.810 -87.490 ;
        RECT -256.110 -87.970 -252.890 -87.490 ;
        RECT -246.190 -87.970 -242.970 -87.490 ;
        RECT -236.270 -87.970 -233.050 -87.490 ;
        RECT -226.350 -87.970 -223.130 -87.490 ;
        RECT -216.430 -87.970 -213.210 -87.490 ;
        RECT -206.510 -87.970 -203.290 -87.490 ;
        RECT -196.590 -87.970 -193.370 -87.490 ;
        RECT -186.670 -87.970 -183.450 -87.490 ;
        RECT -176.750 -87.970 -173.530 -87.490 ;
        RECT -166.830 -87.970 -163.610 -87.490 ;
        RECT -156.910 -87.970 -153.690 -87.490 ;
        RECT -146.990 -87.970 -143.770 -87.490 ;
        RECT -137.070 -87.970 -133.850 -87.490 ;
        RECT -127.150 -87.970 -123.930 -87.490 ;
        RECT -117.230 -87.970 -114.010 -87.490 ;
        RECT -107.310 -87.970 -104.090 -87.490 ;
        RECT -97.390 -87.970 -94.170 -87.490 ;
        RECT -87.470 -87.970 -84.250 -87.490 ;
        RECT -77.550 -87.970 -74.330 -87.490 ;
        RECT -67.630 -87.970 -64.410 -87.490 ;
        RECT -57.710 -87.970 -54.490 -87.490 ;
        RECT -47.790 -87.970 -44.570 -87.490 ;
        RECT -37.870 -87.970 -34.650 -87.490 ;
        RECT -27.950 -87.970 -24.730 -87.490 ;
        RECT -18.030 -87.970 -14.810 -87.490 ;
        RECT -8.110 -87.970 -4.890 -87.490 ;
        RECT 1.810 -87.970 5.030 -87.490 ;
        RECT 11.730 -87.970 14.950 -87.490 ;
        RECT 21.650 -87.970 24.870 -87.490 ;
        RECT -280.910 -90.690 -277.690 -90.210 ;
        RECT -270.990 -90.690 -267.770 -90.210 ;
        RECT -261.070 -90.690 -257.850 -90.210 ;
        RECT -251.150 -90.690 -247.930 -90.210 ;
        RECT -241.230 -90.690 -238.010 -90.210 ;
        RECT -231.310 -90.690 -228.090 -90.210 ;
        RECT -221.390 -90.690 -218.170 -90.210 ;
        RECT -211.470 -90.690 -208.250 -90.210 ;
        RECT -201.550 -90.690 -198.330 -90.210 ;
        RECT -191.630 -90.690 -188.410 -90.210 ;
        RECT -181.710 -90.690 -178.490 -90.210 ;
        RECT -171.790 -90.690 -168.570 -90.210 ;
        RECT -161.870 -90.690 -158.650 -90.210 ;
        RECT -151.950 -90.690 -148.730 -90.210 ;
        RECT -142.030 -90.690 -138.810 -90.210 ;
        RECT -132.110 -90.690 -128.890 -90.210 ;
        RECT -122.190 -90.690 -118.970 -90.210 ;
        RECT -112.270 -90.690 -109.050 -90.210 ;
        RECT -102.350 -90.690 -99.130 -90.210 ;
        RECT -92.430 -90.690 -89.210 -90.210 ;
        RECT -82.510 -90.690 -79.290 -90.210 ;
        RECT -72.590 -90.690 -69.370 -90.210 ;
        RECT -62.670 -90.690 -59.450 -90.210 ;
        RECT -52.750 -90.690 -49.530 -90.210 ;
        RECT -42.830 -90.690 -39.610 -90.210 ;
        RECT -32.910 -90.690 -29.690 -90.210 ;
        RECT -22.990 -90.690 -19.770 -90.210 ;
        RECT -13.070 -90.690 -9.850 -90.210 ;
        RECT -3.150 -90.690 0.070 -90.210 ;
        RECT 6.770 -90.690 9.990 -90.210 ;
        RECT 16.690 -90.690 19.910 -90.210 ;
        RECT 26.610 -90.690 28.450 -90.210 ;
        RECT -220.020 -90.700 -218.170 -90.690 ;
        RECT -140.660 -90.700 -138.810 -90.690 ;
        RECT -61.300 -90.700 -59.450 -90.690 ;
        RECT 18.060 -90.700 19.910 -90.690 ;
        RECT -284.970 -92.260 -283.550 -90.880 ;
        RECT -275.050 -92.260 -273.630 -90.880 ;
        RECT -265.130 -92.260 -263.710 -90.880 ;
        RECT -255.210 -92.260 -253.790 -90.880 ;
        RECT -245.290 -92.260 -243.870 -90.880 ;
        RECT -235.370 -92.260 -233.950 -90.880 ;
        RECT -225.450 -92.260 -224.030 -90.880 ;
        RECT -215.530 -92.260 -214.110 -90.880 ;
        RECT -205.610 -92.260 -204.190 -90.880 ;
        RECT -195.690 -92.260 -194.270 -90.880 ;
        RECT -185.770 -92.260 -184.350 -90.880 ;
        RECT -175.850 -92.260 -174.430 -90.880 ;
        RECT -165.930 -92.260 -164.510 -90.880 ;
        RECT -156.010 -92.260 -154.590 -90.880 ;
        RECT -146.090 -92.260 -144.670 -90.880 ;
        RECT -136.170 -92.260 -134.750 -90.880 ;
        RECT -126.250 -92.260 -124.830 -90.880 ;
        RECT -116.330 -92.260 -114.910 -90.880 ;
        RECT -106.410 -92.260 -104.990 -90.880 ;
        RECT -96.490 -92.260 -95.070 -90.880 ;
        RECT -86.570 -92.260 -85.150 -90.880 ;
        RECT -76.650 -92.260 -75.230 -90.880 ;
        RECT -66.730 -92.260 -65.310 -90.880 ;
        RECT -56.810 -92.260 -55.390 -90.880 ;
        RECT -46.890 -92.260 -45.470 -90.880 ;
        RECT -36.970 -92.260 -35.550 -90.880 ;
        RECT -27.050 -92.260 -25.630 -90.880 ;
        RECT -17.130 -92.260 -15.710 -90.880 ;
        RECT -7.210 -92.260 -5.790 -90.880 ;
        RECT 2.710 -92.260 4.130 -90.880 ;
        RECT 12.630 -92.260 14.050 -90.880 ;
        RECT 22.550 -92.260 23.970 -90.880 ;
        RECT -279.280 -173.630 -278.820 -173.625 ;
        RECT -269.360 -173.630 -268.900 -173.625 ;
        RECT -259.440 -173.630 -258.980 -173.625 ;
        RECT -249.520 -173.630 -249.060 -173.625 ;
        RECT -239.600 -173.630 -239.140 -173.625 ;
        RECT -229.680 -173.630 -229.220 -173.625 ;
        RECT -219.760 -173.630 -219.300 -173.625 ;
        RECT -209.840 -173.630 -209.380 -173.625 ;
        RECT -199.920 -173.630 -199.460 -173.625 ;
        RECT -190.000 -173.630 -189.540 -173.625 ;
        RECT -180.080 -173.630 -179.620 -173.625 ;
        RECT -170.160 -173.630 -169.700 -173.625 ;
        RECT -160.240 -173.630 -159.780 -173.625 ;
        RECT -150.320 -173.630 -149.860 -173.625 ;
        RECT -140.400 -173.630 -139.940 -173.625 ;
        RECT -130.480 -173.630 -130.020 -173.625 ;
        RECT -120.560 -173.630 -120.100 -173.625 ;
        RECT -110.640 -173.630 -110.180 -173.625 ;
        RECT -100.720 -173.630 -100.260 -173.625 ;
        RECT -90.800 -173.630 -90.340 -173.625 ;
        RECT -80.880 -173.630 -80.420 -173.625 ;
        RECT -70.960 -173.630 -70.500 -173.625 ;
        RECT -61.040 -173.630 -60.580 -173.625 ;
        RECT -51.120 -173.630 -50.660 -173.625 ;
        RECT -41.200 -173.630 -40.740 -173.625 ;
        RECT -31.280 -173.630 -30.820 -173.625 ;
        RECT -21.360 -173.630 -20.900 -173.625 ;
        RECT -11.440 -173.630 -10.980 -173.625 ;
        RECT -1.520 -173.630 -1.060 -173.625 ;
        RECT 8.400 -173.630 8.860 -173.625 ;
        RECT 18.320 -173.630 18.780 -173.625 ;
        RECT 28.240 -173.630 28.700 -173.625 ;
        RECT -279.760 -175.010 -278.340 -173.630 ;
        RECT -269.840 -175.010 -268.420 -173.630 ;
        RECT -259.920 -175.010 -258.500 -173.630 ;
        RECT -250.000 -175.010 -248.580 -173.630 ;
        RECT -240.080 -175.010 -238.660 -173.630 ;
        RECT -230.160 -175.010 -228.740 -173.630 ;
        RECT -220.240 -175.010 -218.820 -173.630 ;
        RECT -210.320 -175.010 -208.900 -173.630 ;
        RECT -200.400 -175.010 -198.980 -173.630 ;
        RECT -190.480 -175.010 -189.060 -173.630 ;
        RECT -180.560 -175.010 -179.140 -173.630 ;
        RECT -170.640 -175.010 -169.220 -173.630 ;
        RECT -160.720 -175.010 -159.300 -173.630 ;
        RECT -150.800 -175.010 -149.380 -173.630 ;
        RECT -140.880 -175.010 -139.460 -173.630 ;
        RECT -130.960 -175.010 -129.540 -173.630 ;
        RECT -121.040 -175.010 -119.620 -173.630 ;
        RECT -111.120 -175.010 -109.700 -173.630 ;
        RECT -101.200 -175.010 -99.780 -173.630 ;
        RECT -91.280 -175.010 -89.860 -173.630 ;
        RECT -81.360 -175.010 -79.940 -173.630 ;
        RECT -71.440 -175.010 -70.020 -173.630 ;
        RECT -61.520 -175.010 -60.100 -173.630 ;
        RECT -51.600 -175.010 -50.180 -173.630 ;
        RECT -41.680 -175.010 -40.260 -173.630 ;
        RECT -31.760 -175.010 -30.340 -173.630 ;
        RECT -21.840 -175.010 -20.420 -173.630 ;
        RECT -11.920 -175.010 -10.500 -173.630 ;
        RECT -2.000 -175.010 -0.580 -173.630 ;
        RECT 7.920 -175.010 9.340 -173.630 ;
        RECT 17.840 -175.010 19.260 -173.630 ;
        RECT 27.760 -175.010 28.700 -173.630 ;
        RECT -285.620 -175.680 -282.400 -175.200 ;
        RECT -275.700 -175.680 -272.480 -175.200 ;
        RECT -265.780 -175.680 -262.560 -175.200 ;
        RECT -255.860 -175.680 -252.640 -175.200 ;
        RECT -245.940 -175.680 -242.720 -175.200 ;
        RECT -236.020 -175.680 -232.800 -175.200 ;
        RECT -226.100 -175.680 -222.880 -175.200 ;
        RECT -216.180 -175.680 -212.960 -175.200 ;
        RECT -206.260 -175.680 -203.040 -175.200 ;
        RECT -196.340 -175.680 -193.120 -175.200 ;
        RECT -186.420 -175.680 -183.200 -175.200 ;
        RECT -176.500 -175.680 -173.280 -175.200 ;
        RECT -166.580 -175.680 -163.360 -175.200 ;
        RECT -156.660 -175.680 -153.440 -175.200 ;
        RECT -146.740 -175.680 -143.520 -175.200 ;
        RECT -136.820 -175.680 -133.600 -175.200 ;
        RECT -126.900 -175.680 -123.680 -175.200 ;
        RECT -116.980 -175.680 -113.760 -175.200 ;
        RECT -107.060 -175.680 -103.840 -175.200 ;
        RECT -97.140 -175.680 -93.920 -175.200 ;
        RECT -87.220 -175.680 -84.000 -175.200 ;
        RECT -77.300 -175.680 -74.080 -175.200 ;
        RECT -67.380 -175.680 -64.160 -175.200 ;
        RECT -57.460 -175.680 -54.240 -175.200 ;
        RECT -47.540 -175.680 -44.320 -175.200 ;
        RECT -37.620 -175.680 -34.400 -175.200 ;
        RECT -27.700 -175.680 -24.480 -175.200 ;
        RECT -17.780 -175.680 -14.560 -175.200 ;
        RECT -7.860 -175.680 -4.640 -175.200 ;
        RECT 2.060 -175.680 5.280 -175.200 ;
        RECT 11.980 -175.680 15.200 -175.200 ;
        RECT 21.900 -175.680 25.120 -175.200 ;
        RECT -280.660 -178.400 -277.440 -177.920 ;
        RECT -270.740 -178.400 -267.520 -177.920 ;
        RECT -260.820 -178.400 -257.600 -177.920 ;
        RECT -250.900 -178.400 -247.680 -177.920 ;
        RECT -240.980 -178.400 -237.760 -177.920 ;
        RECT -231.060 -178.400 -227.840 -177.920 ;
        RECT -221.140 -178.400 -217.920 -177.920 ;
        RECT -211.220 -178.400 -208.000 -177.920 ;
        RECT -201.300 -178.400 -198.080 -177.920 ;
        RECT -191.380 -178.400 -188.160 -177.920 ;
        RECT -181.460 -178.400 -178.240 -177.920 ;
        RECT -171.540 -178.400 -168.320 -177.920 ;
        RECT -161.620 -178.400 -158.400 -177.920 ;
        RECT -151.700 -178.400 -148.480 -177.920 ;
        RECT -141.780 -178.400 -138.560 -177.920 ;
        RECT -131.860 -178.400 -128.640 -177.920 ;
        RECT -121.940 -178.400 -118.720 -177.920 ;
        RECT -112.020 -178.400 -108.800 -177.920 ;
        RECT -102.100 -178.400 -98.880 -177.920 ;
        RECT -92.180 -178.400 -88.960 -177.920 ;
        RECT -82.260 -178.400 -79.040 -177.920 ;
        RECT -72.340 -178.400 -69.120 -177.920 ;
        RECT -62.420 -178.400 -59.200 -177.920 ;
        RECT -52.500 -178.400 -49.280 -177.920 ;
        RECT -42.580 -178.400 -39.360 -177.920 ;
        RECT -32.660 -178.400 -29.440 -177.920 ;
        RECT -22.740 -178.400 -19.520 -177.920 ;
        RECT -12.820 -178.400 -9.600 -177.920 ;
        RECT -2.900 -178.400 0.320 -177.920 ;
        RECT 7.020 -178.400 10.240 -177.920 ;
        RECT 16.940 -178.400 20.160 -177.920 ;
        RECT 26.860 -178.400 28.700 -177.920 ;
        RECT -219.770 -178.410 -217.920 -178.400 ;
        RECT -140.410 -178.410 -138.560 -178.400 ;
        RECT -61.050 -178.410 -59.200 -178.400 ;
        RECT 18.310 -178.410 20.160 -178.400 ;
        RECT -284.720 -179.970 -283.300 -178.590 ;
        RECT -274.800 -179.970 -273.380 -178.590 ;
        RECT -264.880 -179.970 -263.460 -178.590 ;
        RECT -254.960 -179.970 -253.540 -178.590 ;
        RECT -245.040 -179.970 -243.620 -178.590 ;
        RECT -235.120 -179.970 -233.700 -178.590 ;
        RECT -225.200 -179.970 -223.780 -178.590 ;
        RECT -215.280 -179.970 -213.860 -178.590 ;
        RECT -205.360 -179.970 -203.940 -178.590 ;
        RECT -195.440 -179.970 -194.020 -178.590 ;
        RECT -185.520 -179.970 -184.100 -178.590 ;
        RECT -175.600 -179.970 -174.180 -178.590 ;
        RECT -165.680 -179.970 -164.260 -178.590 ;
        RECT -155.760 -179.970 -154.340 -178.590 ;
        RECT -145.840 -179.970 -144.420 -178.590 ;
        RECT -135.920 -179.970 -134.500 -178.590 ;
        RECT -126.000 -179.970 -124.580 -178.590 ;
        RECT -116.080 -179.970 -114.660 -178.590 ;
        RECT -106.160 -179.970 -104.740 -178.590 ;
        RECT -96.240 -179.970 -94.820 -178.590 ;
        RECT -86.320 -179.970 -84.900 -178.590 ;
        RECT -76.400 -179.970 -74.980 -178.590 ;
        RECT -66.480 -179.970 -65.060 -178.590 ;
        RECT -56.560 -179.970 -55.140 -178.590 ;
        RECT -46.640 -179.970 -45.220 -178.590 ;
        RECT -36.720 -179.970 -35.300 -178.590 ;
        RECT -26.800 -179.970 -25.380 -178.590 ;
        RECT -16.880 -179.970 -15.460 -178.590 ;
        RECT -6.960 -179.970 -5.540 -178.590 ;
        RECT 2.960 -179.970 4.380 -178.590 ;
        RECT 12.880 -179.970 14.300 -178.590 ;
        RECT 22.800 -179.970 24.220 -178.590 ;
      LAYER via ;
        RECT -281.915 94.780 -281.655 95.040 ;
        RECT -280.975 94.770 -280.715 95.030 ;
        RECT -271.285 94.775 -271.025 95.035 ;
        RECT -262.075 94.780 -261.815 95.040 ;
        RECT -261.135 94.770 -260.875 95.030 ;
        RECT -252.155 94.780 -251.895 95.040 ;
        RECT -251.215 94.770 -250.955 95.030 ;
        RECT -242.235 94.780 -241.975 95.040 ;
        RECT -241.295 94.770 -241.035 95.030 ;
        RECT -232.315 94.780 -232.055 95.040 ;
        RECT -231.375 94.770 -231.115 95.030 ;
        RECT -222.395 94.780 -222.135 95.040 ;
        RECT -221.455 94.770 -221.195 95.030 ;
        RECT -212.475 94.780 -212.215 95.040 ;
        RECT -211.535 94.770 -211.275 95.030 ;
        RECT -202.555 94.780 -202.295 95.040 ;
        RECT -201.615 94.770 -201.355 95.030 ;
        RECT -192.635 94.780 -192.375 95.040 ;
        RECT -191.695 94.770 -191.435 95.030 ;
        RECT -182.715 94.780 -182.455 95.040 ;
        RECT -181.775 94.770 -181.515 95.030 ;
        RECT -172.795 94.780 -172.535 95.040 ;
        RECT -171.855 94.770 -171.595 95.030 ;
        RECT -162.875 94.780 -162.615 95.040 ;
        RECT -161.935 94.770 -161.675 95.030 ;
        RECT -152.955 94.780 -152.695 95.040 ;
        RECT -152.015 94.770 -151.755 95.030 ;
        RECT -143.035 94.780 -142.775 95.040 ;
        RECT -142.095 94.770 -141.835 95.030 ;
        RECT -133.115 94.780 -132.855 95.040 ;
        RECT -132.175 94.770 -131.915 95.030 ;
        RECT -123.195 94.780 -122.935 95.040 ;
        RECT -122.255 94.770 -121.995 95.030 ;
        RECT -113.275 94.780 -113.015 95.040 ;
        RECT -112.335 94.770 -112.075 95.030 ;
        RECT -103.355 94.780 -103.095 95.040 ;
        RECT -102.415 94.770 -102.155 95.030 ;
        RECT -93.435 94.780 -93.175 95.040 ;
        RECT -92.495 94.770 -92.235 95.030 ;
        RECT -83.515 94.780 -83.255 95.040 ;
        RECT -82.575 94.770 -82.315 95.030 ;
        RECT -73.595 94.780 -73.335 95.040 ;
        RECT -72.655 94.770 -72.395 95.030 ;
        RECT -63.675 94.780 -63.415 95.040 ;
        RECT -62.735 94.770 -62.475 95.030 ;
        RECT -53.755 94.780 -53.495 95.040 ;
        RECT -52.815 94.770 -52.555 95.030 ;
        RECT -43.835 94.780 -43.575 95.040 ;
        RECT -42.895 94.770 -42.635 95.030 ;
        RECT -33.915 94.780 -33.655 95.040 ;
        RECT -32.975 94.770 -32.715 95.030 ;
        RECT -23.995 94.780 -23.735 95.040 ;
        RECT -23.055 94.770 -22.795 95.030 ;
        RECT -14.075 94.780 -13.815 95.040 ;
        RECT -13.135 94.770 -12.875 95.030 ;
        RECT -4.155 94.780 -3.895 95.040 ;
        RECT -3.215 94.770 -2.955 95.030 ;
        RECT 5.765 94.780 6.025 95.040 ;
        RECT 6.705 94.770 6.965 95.030 ;
        RECT 15.685 94.780 15.945 95.040 ;
        RECT 16.625 94.770 16.885 95.030 ;
        RECT 25.605 94.780 25.865 95.040 ;
        RECT -286.635 93.190 -286.375 93.450 ;
        RECT -286.175 93.190 -285.915 93.450 ;
        RECT -276.715 93.190 -276.455 93.450 ;
        RECT -276.255 93.190 -275.995 93.450 ;
        RECT -266.795 93.190 -266.535 93.450 ;
        RECT -266.335 93.190 -266.075 93.450 ;
        RECT -256.875 93.190 -256.615 93.450 ;
        RECT -256.415 93.190 -256.155 93.450 ;
        RECT -246.955 93.190 -246.695 93.450 ;
        RECT -246.495 93.190 -246.235 93.450 ;
        RECT -237.035 93.190 -236.775 93.450 ;
        RECT -236.575 93.190 -236.315 93.450 ;
        RECT -227.115 93.190 -226.855 93.450 ;
        RECT -226.655 93.190 -226.395 93.450 ;
        RECT -217.195 93.190 -216.935 93.450 ;
        RECT -216.735 93.190 -216.475 93.450 ;
        RECT -207.275 93.190 -207.015 93.450 ;
        RECT -206.815 93.190 -206.555 93.450 ;
        RECT -197.355 93.190 -197.095 93.450 ;
        RECT -196.895 93.190 -196.635 93.450 ;
        RECT -187.435 93.190 -187.175 93.450 ;
        RECT -186.975 93.190 -186.715 93.450 ;
        RECT -177.515 93.190 -177.255 93.450 ;
        RECT -177.055 93.190 -176.795 93.450 ;
        RECT -167.595 93.190 -167.335 93.450 ;
        RECT -167.135 93.190 -166.875 93.450 ;
        RECT -157.675 93.190 -157.415 93.450 ;
        RECT -157.215 93.190 -156.955 93.450 ;
        RECT -147.755 93.190 -147.495 93.450 ;
        RECT -147.295 93.190 -147.035 93.450 ;
        RECT -137.835 93.190 -137.575 93.450 ;
        RECT -137.375 93.190 -137.115 93.450 ;
        RECT -127.915 93.190 -127.655 93.450 ;
        RECT -127.455 93.190 -127.195 93.450 ;
        RECT -117.995 93.190 -117.735 93.450 ;
        RECT -117.535 93.190 -117.275 93.450 ;
        RECT -108.075 93.190 -107.815 93.450 ;
        RECT -107.615 93.190 -107.355 93.450 ;
        RECT -98.155 93.190 -97.895 93.450 ;
        RECT -97.695 93.190 -97.435 93.450 ;
        RECT -88.235 93.190 -87.975 93.450 ;
        RECT -87.775 93.190 -87.515 93.450 ;
        RECT -78.315 93.190 -78.055 93.450 ;
        RECT -77.855 93.190 -77.595 93.450 ;
        RECT -68.395 93.190 -68.135 93.450 ;
        RECT -67.935 93.190 -67.675 93.450 ;
        RECT -58.475 93.190 -58.215 93.450 ;
        RECT -58.015 93.190 -57.755 93.450 ;
        RECT -48.555 93.190 -48.295 93.450 ;
        RECT -48.095 93.190 -47.835 93.450 ;
        RECT -38.635 93.190 -38.375 93.450 ;
        RECT -38.175 93.190 -37.915 93.450 ;
        RECT -28.715 93.190 -28.455 93.450 ;
        RECT -28.255 93.190 -27.995 93.450 ;
        RECT -18.795 93.190 -18.535 93.450 ;
        RECT -18.335 93.190 -18.075 93.450 ;
        RECT -8.875 93.190 -8.615 93.450 ;
        RECT -8.415 93.190 -8.155 93.450 ;
        RECT 1.045 93.190 1.305 93.450 ;
        RECT 1.505 93.190 1.765 93.450 ;
        RECT 10.965 93.190 11.225 93.450 ;
        RECT 11.425 93.190 11.685 93.450 ;
        RECT 20.885 93.190 21.145 93.450 ;
        RECT 21.345 93.190 21.605 93.450 ;
        RECT -281.675 90.480 -281.415 90.740 ;
        RECT -281.215 90.480 -280.955 90.740 ;
        RECT -271.755 90.480 -271.495 90.740 ;
        RECT -271.295 90.480 -271.035 90.740 ;
        RECT -261.835 90.480 -261.575 90.740 ;
        RECT -261.375 90.480 -261.115 90.740 ;
        RECT -251.915 90.480 -251.655 90.740 ;
        RECT -251.455 90.480 -251.195 90.740 ;
        RECT -241.995 90.480 -241.735 90.740 ;
        RECT -241.535 90.480 -241.275 90.740 ;
        RECT -232.075 90.480 -231.815 90.740 ;
        RECT -231.615 90.480 -231.355 90.740 ;
        RECT -222.155 90.480 -221.895 90.740 ;
        RECT -221.695 90.480 -221.435 90.740 ;
        RECT -212.235 90.480 -211.975 90.740 ;
        RECT -211.775 90.480 -211.515 90.740 ;
        RECT -202.315 90.480 -202.055 90.740 ;
        RECT -201.855 90.480 -201.595 90.740 ;
        RECT -192.395 90.480 -192.135 90.740 ;
        RECT -191.935 90.480 -191.675 90.740 ;
        RECT -182.475 90.480 -182.215 90.740 ;
        RECT -182.015 90.480 -181.755 90.740 ;
        RECT -172.555 90.480 -172.295 90.740 ;
        RECT -172.095 90.480 -171.835 90.740 ;
        RECT -162.635 90.480 -162.375 90.740 ;
        RECT -162.175 90.480 -161.915 90.740 ;
        RECT -152.715 90.480 -152.455 90.740 ;
        RECT -152.255 90.480 -151.995 90.740 ;
        RECT -142.795 90.480 -142.535 90.740 ;
        RECT -142.335 90.480 -142.075 90.740 ;
        RECT -132.875 90.480 -132.615 90.740 ;
        RECT -132.415 90.480 -132.155 90.740 ;
        RECT -122.955 90.480 -122.695 90.740 ;
        RECT -122.495 90.480 -122.235 90.740 ;
        RECT -113.035 90.480 -112.775 90.740 ;
        RECT -112.575 90.480 -112.315 90.740 ;
        RECT -103.115 90.480 -102.855 90.740 ;
        RECT -102.655 90.480 -102.395 90.740 ;
        RECT -93.195 90.480 -92.935 90.740 ;
        RECT -92.735 90.480 -92.475 90.740 ;
        RECT -83.275 90.480 -83.015 90.740 ;
        RECT -82.815 90.480 -82.555 90.740 ;
        RECT -73.355 90.480 -73.095 90.740 ;
        RECT -72.895 90.480 -72.635 90.740 ;
        RECT -63.435 90.480 -63.175 90.740 ;
        RECT -62.975 90.480 -62.715 90.740 ;
        RECT -53.515 90.480 -53.255 90.740 ;
        RECT -53.055 90.480 -52.795 90.740 ;
        RECT -43.595 90.480 -43.335 90.740 ;
        RECT -43.135 90.480 -42.875 90.740 ;
        RECT -33.675 90.480 -33.415 90.740 ;
        RECT -33.215 90.480 -32.955 90.740 ;
        RECT -23.755 90.480 -23.495 90.740 ;
        RECT -23.295 90.480 -23.035 90.740 ;
        RECT -13.835 90.480 -13.575 90.740 ;
        RECT -13.375 90.480 -13.115 90.740 ;
        RECT -3.915 90.480 -3.655 90.740 ;
        RECT -3.455 90.480 -3.195 90.740 ;
        RECT 6.005 90.480 6.265 90.740 ;
        RECT 6.465 90.480 6.725 90.740 ;
        RECT 15.925 90.480 16.185 90.740 ;
        RECT 16.385 90.480 16.645 90.740 ;
        RECT 25.845 90.480 26.105 90.740 ;
        RECT -286.865 88.890 -286.605 89.150 ;
        RECT -285.935 88.890 -285.675 89.150 ;
        RECT -276.945 88.890 -276.685 89.150 ;
        RECT -276.015 88.890 -275.755 89.150 ;
        RECT -267.025 88.890 -266.765 89.150 ;
        RECT -266.095 88.890 -265.835 89.150 ;
        RECT -257.105 88.890 -256.845 89.150 ;
        RECT -256.175 88.890 -255.915 89.150 ;
        RECT -247.185 88.890 -246.925 89.150 ;
        RECT -246.255 88.890 -245.995 89.150 ;
        RECT -237.265 88.890 -237.005 89.150 ;
        RECT -236.335 88.890 -236.075 89.150 ;
        RECT -227.345 88.890 -227.085 89.150 ;
        RECT -226.415 88.890 -226.155 89.150 ;
        RECT -217.425 88.890 -217.165 89.150 ;
        RECT -216.495 88.890 -216.235 89.150 ;
        RECT -207.505 88.890 -207.245 89.150 ;
        RECT -206.575 88.890 -206.315 89.150 ;
        RECT -197.585 88.890 -197.325 89.150 ;
        RECT -196.655 88.890 -196.395 89.150 ;
        RECT -187.665 88.890 -187.405 89.150 ;
        RECT -186.735 88.890 -186.475 89.150 ;
        RECT -177.745 88.890 -177.485 89.150 ;
        RECT -176.815 88.890 -176.555 89.150 ;
        RECT -167.825 88.890 -167.565 89.150 ;
        RECT -166.895 88.890 -166.635 89.150 ;
        RECT -157.905 88.890 -157.645 89.150 ;
        RECT -156.975 88.890 -156.715 89.150 ;
        RECT -147.985 88.890 -147.725 89.150 ;
        RECT -147.055 88.890 -146.795 89.150 ;
        RECT -138.065 88.890 -137.805 89.150 ;
        RECT -137.135 88.890 -136.875 89.150 ;
        RECT -128.145 88.890 -127.885 89.150 ;
        RECT -127.215 88.890 -126.955 89.150 ;
        RECT -118.225 88.890 -117.965 89.150 ;
        RECT -117.295 88.890 -117.035 89.150 ;
        RECT -108.305 88.890 -108.045 89.150 ;
        RECT -107.375 88.890 -107.115 89.150 ;
        RECT -98.385 88.890 -98.125 89.150 ;
        RECT -97.455 88.890 -97.195 89.150 ;
        RECT -88.465 88.890 -88.205 89.150 ;
        RECT -87.535 88.890 -87.275 89.150 ;
        RECT -78.545 88.890 -78.285 89.150 ;
        RECT -77.615 88.890 -77.355 89.150 ;
        RECT -68.625 88.890 -68.365 89.150 ;
        RECT -67.695 88.890 -67.435 89.150 ;
        RECT -58.705 88.890 -58.445 89.150 ;
        RECT -57.775 88.890 -57.515 89.150 ;
        RECT -48.785 88.890 -48.525 89.150 ;
        RECT -47.855 88.890 -47.595 89.150 ;
        RECT -38.865 88.890 -38.605 89.150 ;
        RECT -37.935 88.890 -37.675 89.150 ;
        RECT -28.945 88.890 -28.685 89.150 ;
        RECT -28.015 88.890 -27.755 89.150 ;
        RECT -19.025 88.890 -18.765 89.150 ;
        RECT -18.095 88.890 -17.835 89.150 ;
        RECT -9.105 88.890 -8.845 89.150 ;
        RECT -8.175 88.890 -7.915 89.150 ;
        RECT 0.815 88.890 1.075 89.150 ;
        RECT 1.745 88.890 2.005 89.150 ;
        RECT 10.735 88.890 10.995 89.150 ;
        RECT 11.665 88.890 11.925 89.150 ;
        RECT 20.655 88.890 20.915 89.150 ;
        RECT 21.585 88.890 21.845 89.150 ;
        RECT -281.665 7.070 -281.405 7.330 ;
        RECT -280.725 7.060 -280.465 7.320 ;
        RECT -271.035 7.065 -270.775 7.325 ;
        RECT -261.825 7.070 -261.565 7.330 ;
        RECT -260.885 7.060 -260.625 7.320 ;
        RECT -251.905 7.070 -251.645 7.330 ;
        RECT -250.965 7.060 -250.705 7.320 ;
        RECT -241.985 7.070 -241.725 7.330 ;
        RECT -241.045 7.060 -240.785 7.320 ;
        RECT -232.065 7.070 -231.805 7.330 ;
        RECT -231.125 7.060 -230.865 7.320 ;
        RECT -222.145 7.070 -221.885 7.330 ;
        RECT -221.205 7.060 -220.945 7.320 ;
        RECT -212.225 7.070 -211.965 7.330 ;
        RECT -211.285 7.060 -211.025 7.320 ;
        RECT -202.305 7.070 -202.045 7.330 ;
        RECT -201.365 7.060 -201.105 7.320 ;
        RECT -192.385 7.070 -192.125 7.330 ;
        RECT -191.445 7.060 -191.185 7.320 ;
        RECT -182.465 7.070 -182.205 7.330 ;
        RECT -181.525 7.060 -181.265 7.320 ;
        RECT -172.545 7.070 -172.285 7.330 ;
        RECT -171.605 7.060 -171.345 7.320 ;
        RECT -162.625 7.070 -162.365 7.330 ;
        RECT -161.685 7.060 -161.425 7.320 ;
        RECT -152.705 7.070 -152.445 7.330 ;
        RECT -151.765 7.060 -151.505 7.320 ;
        RECT -142.785 7.070 -142.525 7.330 ;
        RECT -141.845 7.060 -141.585 7.320 ;
        RECT -132.865 7.070 -132.605 7.330 ;
        RECT -131.925 7.060 -131.665 7.320 ;
        RECT -122.945 7.070 -122.685 7.330 ;
        RECT -122.005 7.060 -121.745 7.320 ;
        RECT -113.025 7.070 -112.765 7.330 ;
        RECT -112.085 7.060 -111.825 7.320 ;
        RECT -103.105 7.070 -102.845 7.330 ;
        RECT -102.165 7.060 -101.905 7.320 ;
        RECT -93.185 7.070 -92.925 7.330 ;
        RECT -92.245 7.060 -91.985 7.320 ;
        RECT -83.265 7.070 -83.005 7.330 ;
        RECT -82.325 7.060 -82.065 7.320 ;
        RECT -73.345 7.070 -73.085 7.330 ;
        RECT -72.405 7.060 -72.145 7.320 ;
        RECT -63.425 7.070 -63.165 7.330 ;
        RECT -62.485 7.060 -62.225 7.320 ;
        RECT -53.505 7.070 -53.245 7.330 ;
        RECT -52.565 7.060 -52.305 7.320 ;
        RECT -43.585 7.070 -43.325 7.330 ;
        RECT -42.645 7.060 -42.385 7.320 ;
        RECT -33.665 7.070 -33.405 7.330 ;
        RECT -32.725 7.060 -32.465 7.320 ;
        RECT -23.745 7.070 -23.485 7.330 ;
        RECT -22.805 7.060 -22.545 7.320 ;
        RECT -13.825 7.070 -13.565 7.330 ;
        RECT -12.885 7.060 -12.625 7.320 ;
        RECT -3.905 7.070 -3.645 7.330 ;
        RECT -2.965 7.060 -2.705 7.320 ;
        RECT 6.015 7.070 6.275 7.330 ;
        RECT 6.955 7.060 7.215 7.320 ;
        RECT 15.935 7.070 16.195 7.330 ;
        RECT 16.875 7.060 17.135 7.320 ;
        RECT 25.855 7.070 26.115 7.330 ;
        RECT -286.385 5.480 -286.125 5.740 ;
        RECT -285.925 5.480 -285.665 5.740 ;
        RECT -276.465 5.480 -276.205 5.740 ;
        RECT -276.005 5.480 -275.745 5.740 ;
        RECT -266.545 5.480 -266.285 5.740 ;
        RECT -266.085 5.480 -265.825 5.740 ;
        RECT -256.625 5.480 -256.365 5.740 ;
        RECT -256.165 5.480 -255.905 5.740 ;
        RECT -246.705 5.480 -246.445 5.740 ;
        RECT -246.245 5.480 -245.985 5.740 ;
        RECT -236.785 5.480 -236.525 5.740 ;
        RECT -236.325 5.480 -236.065 5.740 ;
        RECT -226.865 5.480 -226.605 5.740 ;
        RECT -226.405 5.480 -226.145 5.740 ;
        RECT -216.945 5.480 -216.685 5.740 ;
        RECT -216.485 5.480 -216.225 5.740 ;
        RECT -207.025 5.480 -206.765 5.740 ;
        RECT -206.565 5.480 -206.305 5.740 ;
        RECT -197.105 5.480 -196.845 5.740 ;
        RECT -196.645 5.480 -196.385 5.740 ;
        RECT -187.185 5.480 -186.925 5.740 ;
        RECT -186.725 5.480 -186.465 5.740 ;
        RECT -177.265 5.480 -177.005 5.740 ;
        RECT -176.805 5.480 -176.545 5.740 ;
        RECT -167.345 5.480 -167.085 5.740 ;
        RECT -166.885 5.480 -166.625 5.740 ;
        RECT -157.425 5.480 -157.165 5.740 ;
        RECT -156.965 5.480 -156.705 5.740 ;
        RECT -147.505 5.480 -147.245 5.740 ;
        RECT -147.045 5.480 -146.785 5.740 ;
        RECT -137.585 5.480 -137.325 5.740 ;
        RECT -137.125 5.480 -136.865 5.740 ;
        RECT -127.665 5.480 -127.405 5.740 ;
        RECT -127.205 5.480 -126.945 5.740 ;
        RECT -117.745 5.480 -117.485 5.740 ;
        RECT -117.285 5.480 -117.025 5.740 ;
        RECT -107.825 5.480 -107.565 5.740 ;
        RECT -107.365 5.480 -107.105 5.740 ;
        RECT -97.905 5.480 -97.645 5.740 ;
        RECT -97.445 5.480 -97.185 5.740 ;
        RECT -87.985 5.480 -87.725 5.740 ;
        RECT -87.525 5.480 -87.265 5.740 ;
        RECT -78.065 5.480 -77.805 5.740 ;
        RECT -77.605 5.480 -77.345 5.740 ;
        RECT -68.145 5.480 -67.885 5.740 ;
        RECT -67.685 5.480 -67.425 5.740 ;
        RECT -58.225 5.480 -57.965 5.740 ;
        RECT -57.765 5.480 -57.505 5.740 ;
        RECT -48.305 5.480 -48.045 5.740 ;
        RECT -47.845 5.480 -47.585 5.740 ;
        RECT -38.385 5.480 -38.125 5.740 ;
        RECT -37.925 5.480 -37.665 5.740 ;
        RECT -28.465 5.480 -28.205 5.740 ;
        RECT -28.005 5.480 -27.745 5.740 ;
        RECT -18.545 5.480 -18.285 5.740 ;
        RECT -18.085 5.480 -17.825 5.740 ;
        RECT -8.625 5.480 -8.365 5.740 ;
        RECT -8.165 5.480 -7.905 5.740 ;
        RECT 1.295 5.480 1.555 5.740 ;
        RECT 1.755 5.480 2.015 5.740 ;
        RECT 11.215 5.480 11.475 5.740 ;
        RECT 11.675 5.480 11.935 5.740 ;
        RECT 21.135 5.480 21.395 5.740 ;
        RECT 21.595 5.480 21.855 5.740 ;
        RECT -281.425 2.770 -281.165 3.030 ;
        RECT -280.965 2.770 -280.705 3.030 ;
        RECT -271.505 2.770 -271.245 3.030 ;
        RECT -271.045 2.770 -270.785 3.030 ;
        RECT -261.585 2.770 -261.325 3.030 ;
        RECT -261.125 2.770 -260.865 3.030 ;
        RECT -251.665 2.770 -251.405 3.030 ;
        RECT -251.205 2.770 -250.945 3.030 ;
        RECT -241.745 2.770 -241.485 3.030 ;
        RECT -241.285 2.770 -241.025 3.030 ;
        RECT -231.825 2.770 -231.565 3.030 ;
        RECT -231.365 2.770 -231.105 3.030 ;
        RECT -221.905 2.770 -221.645 3.030 ;
        RECT -221.445 2.770 -221.185 3.030 ;
        RECT -211.985 2.770 -211.725 3.030 ;
        RECT -211.525 2.770 -211.265 3.030 ;
        RECT -202.065 2.770 -201.805 3.030 ;
        RECT -201.605 2.770 -201.345 3.030 ;
        RECT -192.145 2.770 -191.885 3.030 ;
        RECT -191.685 2.770 -191.425 3.030 ;
        RECT -182.225 2.770 -181.965 3.030 ;
        RECT -181.765 2.770 -181.505 3.030 ;
        RECT -172.305 2.770 -172.045 3.030 ;
        RECT -171.845 2.770 -171.585 3.030 ;
        RECT -162.385 2.770 -162.125 3.030 ;
        RECT -161.925 2.770 -161.665 3.030 ;
        RECT -152.465 2.770 -152.205 3.030 ;
        RECT -152.005 2.770 -151.745 3.030 ;
        RECT -142.545 2.770 -142.285 3.030 ;
        RECT -142.085 2.770 -141.825 3.030 ;
        RECT -132.625 2.770 -132.365 3.030 ;
        RECT -132.165 2.770 -131.905 3.030 ;
        RECT -122.705 2.770 -122.445 3.030 ;
        RECT -122.245 2.770 -121.985 3.030 ;
        RECT -112.785 2.770 -112.525 3.030 ;
        RECT -112.325 2.770 -112.065 3.030 ;
        RECT -102.865 2.770 -102.605 3.030 ;
        RECT -102.405 2.770 -102.145 3.030 ;
        RECT -92.945 2.770 -92.685 3.030 ;
        RECT -92.485 2.770 -92.225 3.030 ;
        RECT -83.025 2.770 -82.765 3.030 ;
        RECT -82.565 2.770 -82.305 3.030 ;
        RECT -73.105 2.770 -72.845 3.030 ;
        RECT -72.645 2.770 -72.385 3.030 ;
        RECT -63.185 2.770 -62.925 3.030 ;
        RECT -62.725 2.770 -62.465 3.030 ;
        RECT -53.265 2.770 -53.005 3.030 ;
        RECT -52.805 2.770 -52.545 3.030 ;
        RECT -43.345 2.770 -43.085 3.030 ;
        RECT -42.885 2.770 -42.625 3.030 ;
        RECT -33.425 2.770 -33.165 3.030 ;
        RECT -32.965 2.770 -32.705 3.030 ;
        RECT -23.505 2.770 -23.245 3.030 ;
        RECT -23.045 2.770 -22.785 3.030 ;
        RECT -13.585 2.770 -13.325 3.030 ;
        RECT -13.125 2.770 -12.865 3.030 ;
        RECT -3.665 2.770 -3.405 3.030 ;
        RECT -3.205 2.770 -2.945 3.030 ;
        RECT 6.255 2.770 6.515 3.030 ;
        RECT 6.715 2.770 6.975 3.030 ;
        RECT 16.175 2.770 16.435 3.030 ;
        RECT 16.635 2.770 16.895 3.030 ;
        RECT 26.095 2.770 26.355 3.030 ;
        RECT -286.615 1.180 -286.355 1.440 ;
        RECT -285.685 1.180 -285.425 1.440 ;
        RECT -276.695 1.180 -276.435 1.440 ;
        RECT -275.765 1.180 -275.505 1.440 ;
        RECT -266.775 1.180 -266.515 1.440 ;
        RECT -265.845 1.180 -265.585 1.440 ;
        RECT -256.855 1.180 -256.595 1.440 ;
        RECT -255.925 1.180 -255.665 1.440 ;
        RECT -246.935 1.180 -246.675 1.440 ;
        RECT -246.005 1.180 -245.745 1.440 ;
        RECT -237.015 1.180 -236.755 1.440 ;
        RECT -236.085 1.180 -235.825 1.440 ;
        RECT -227.095 1.180 -226.835 1.440 ;
        RECT -226.165 1.180 -225.905 1.440 ;
        RECT -217.175 1.180 -216.915 1.440 ;
        RECT -216.245 1.180 -215.985 1.440 ;
        RECT -207.255 1.180 -206.995 1.440 ;
        RECT -206.325 1.180 -206.065 1.440 ;
        RECT -197.335 1.180 -197.075 1.440 ;
        RECT -196.405 1.180 -196.145 1.440 ;
        RECT -187.415 1.180 -187.155 1.440 ;
        RECT -186.485 1.180 -186.225 1.440 ;
        RECT -177.495 1.180 -177.235 1.440 ;
        RECT -176.565 1.180 -176.305 1.440 ;
        RECT -167.575 1.180 -167.315 1.440 ;
        RECT -166.645 1.180 -166.385 1.440 ;
        RECT -157.655 1.180 -157.395 1.440 ;
        RECT -156.725 1.180 -156.465 1.440 ;
        RECT -147.735 1.180 -147.475 1.440 ;
        RECT -146.805 1.180 -146.545 1.440 ;
        RECT -137.815 1.180 -137.555 1.440 ;
        RECT -136.885 1.180 -136.625 1.440 ;
        RECT -127.895 1.180 -127.635 1.440 ;
        RECT -126.965 1.180 -126.705 1.440 ;
        RECT -117.975 1.180 -117.715 1.440 ;
        RECT -117.045 1.180 -116.785 1.440 ;
        RECT -108.055 1.180 -107.795 1.440 ;
        RECT -107.125 1.180 -106.865 1.440 ;
        RECT -98.135 1.180 -97.875 1.440 ;
        RECT -97.205 1.180 -96.945 1.440 ;
        RECT -88.215 1.180 -87.955 1.440 ;
        RECT -87.285 1.180 -87.025 1.440 ;
        RECT -78.295 1.180 -78.035 1.440 ;
        RECT -77.365 1.180 -77.105 1.440 ;
        RECT -68.375 1.180 -68.115 1.440 ;
        RECT -67.445 1.180 -67.185 1.440 ;
        RECT -58.455 1.180 -58.195 1.440 ;
        RECT -57.525 1.180 -57.265 1.440 ;
        RECT -48.535 1.180 -48.275 1.440 ;
        RECT -47.605 1.180 -47.345 1.440 ;
        RECT -38.615 1.180 -38.355 1.440 ;
        RECT -37.685 1.180 -37.425 1.440 ;
        RECT -28.695 1.180 -28.435 1.440 ;
        RECT -27.765 1.180 -27.505 1.440 ;
        RECT -18.775 1.180 -18.515 1.440 ;
        RECT -17.845 1.180 -17.585 1.440 ;
        RECT -8.855 1.180 -8.595 1.440 ;
        RECT -7.925 1.180 -7.665 1.440 ;
        RECT 1.065 1.180 1.325 1.440 ;
        RECT 1.995 1.180 2.255 1.440 ;
        RECT 10.985 1.180 11.245 1.440 ;
        RECT 11.915 1.180 12.175 1.440 ;
        RECT 20.905 1.180 21.165 1.440 ;
        RECT 21.835 1.180 22.095 1.440 ;
        RECT -279.905 -86.280 -279.645 -86.020 ;
        RECT -278.965 -86.290 -278.705 -86.030 ;
        RECT -269.275 -86.285 -269.015 -86.025 ;
        RECT -260.065 -86.280 -259.805 -86.020 ;
        RECT -259.125 -86.290 -258.865 -86.030 ;
        RECT -250.145 -86.280 -249.885 -86.020 ;
        RECT -249.205 -86.290 -248.945 -86.030 ;
        RECT -240.225 -86.280 -239.965 -86.020 ;
        RECT -239.285 -86.290 -239.025 -86.030 ;
        RECT -230.305 -86.280 -230.045 -86.020 ;
        RECT -229.365 -86.290 -229.105 -86.030 ;
        RECT -220.385 -86.280 -220.125 -86.020 ;
        RECT -219.445 -86.290 -219.185 -86.030 ;
        RECT -210.465 -86.280 -210.205 -86.020 ;
        RECT -209.525 -86.290 -209.265 -86.030 ;
        RECT -200.545 -86.280 -200.285 -86.020 ;
        RECT -199.605 -86.290 -199.345 -86.030 ;
        RECT -190.625 -86.280 -190.365 -86.020 ;
        RECT -189.685 -86.290 -189.425 -86.030 ;
        RECT -180.705 -86.280 -180.445 -86.020 ;
        RECT -179.765 -86.290 -179.505 -86.030 ;
        RECT -170.785 -86.280 -170.525 -86.020 ;
        RECT -169.845 -86.290 -169.585 -86.030 ;
        RECT -160.865 -86.280 -160.605 -86.020 ;
        RECT -159.925 -86.290 -159.665 -86.030 ;
        RECT -150.945 -86.280 -150.685 -86.020 ;
        RECT -150.005 -86.290 -149.745 -86.030 ;
        RECT -141.025 -86.280 -140.765 -86.020 ;
        RECT -140.085 -86.290 -139.825 -86.030 ;
        RECT -131.105 -86.280 -130.845 -86.020 ;
        RECT -130.165 -86.290 -129.905 -86.030 ;
        RECT -121.185 -86.280 -120.925 -86.020 ;
        RECT -120.245 -86.290 -119.985 -86.030 ;
        RECT -111.265 -86.280 -111.005 -86.020 ;
        RECT -110.325 -86.290 -110.065 -86.030 ;
        RECT -101.345 -86.280 -101.085 -86.020 ;
        RECT -100.405 -86.290 -100.145 -86.030 ;
        RECT -91.425 -86.280 -91.165 -86.020 ;
        RECT -90.485 -86.290 -90.225 -86.030 ;
        RECT -81.505 -86.280 -81.245 -86.020 ;
        RECT -80.565 -86.290 -80.305 -86.030 ;
        RECT -71.585 -86.280 -71.325 -86.020 ;
        RECT -70.645 -86.290 -70.385 -86.030 ;
        RECT -61.665 -86.280 -61.405 -86.020 ;
        RECT -60.725 -86.290 -60.465 -86.030 ;
        RECT -51.745 -86.280 -51.485 -86.020 ;
        RECT -50.805 -86.290 -50.545 -86.030 ;
        RECT -41.825 -86.280 -41.565 -86.020 ;
        RECT -40.885 -86.290 -40.625 -86.030 ;
        RECT -31.905 -86.280 -31.645 -86.020 ;
        RECT -30.965 -86.290 -30.705 -86.030 ;
        RECT -21.985 -86.280 -21.725 -86.020 ;
        RECT -21.045 -86.290 -20.785 -86.030 ;
        RECT -12.065 -86.280 -11.805 -86.020 ;
        RECT -11.125 -86.290 -10.865 -86.030 ;
        RECT -2.145 -86.280 -1.885 -86.020 ;
        RECT -1.205 -86.290 -0.945 -86.030 ;
        RECT 7.775 -86.280 8.035 -86.020 ;
        RECT 8.715 -86.290 8.975 -86.030 ;
        RECT 17.695 -86.280 17.955 -86.020 ;
        RECT 18.635 -86.290 18.895 -86.030 ;
        RECT 27.615 -86.280 27.875 -86.020 ;
        RECT -284.625 -87.870 -284.365 -87.610 ;
        RECT -284.165 -87.870 -283.905 -87.610 ;
        RECT -274.705 -87.870 -274.445 -87.610 ;
        RECT -274.245 -87.870 -273.985 -87.610 ;
        RECT -264.785 -87.870 -264.525 -87.610 ;
        RECT -264.325 -87.870 -264.065 -87.610 ;
        RECT -254.865 -87.870 -254.605 -87.610 ;
        RECT -254.405 -87.870 -254.145 -87.610 ;
        RECT -244.945 -87.870 -244.685 -87.610 ;
        RECT -244.485 -87.870 -244.225 -87.610 ;
        RECT -235.025 -87.870 -234.765 -87.610 ;
        RECT -234.565 -87.870 -234.305 -87.610 ;
        RECT -225.105 -87.870 -224.845 -87.610 ;
        RECT -224.645 -87.870 -224.385 -87.610 ;
        RECT -215.185 -87.870 -214.925 -87.610 ;
        RECT -214.725 -87.870 -214.465 -87.610 ;
        RECT -205.265 -87.870 -205.005 -87.610 ;
        RECT -204.805 -87.870 -204.545 -87.610 ;
        RECT -195.345 -87.870 -195.085 -87.610 ;
        RECT -194.885 -87.870 -194.625 -87.610 ;
        RECT -185.425 -87.870 -185.165 -87.610 ;
        RECT -184.965 -87.870 -184.705 -87.610 ;
        RECT -175.505 -87.870 -175.245 -87.610 ;
        RECT -175.045 -87.870 -174.785 -87.610 ;
        RECT -165.585 -87.870 -165.325 -87.610 ;
        RECT -165.125 -87.870 -164.865 -87.610 ;
        RECT -155.665 -87.870 -155.405 -87.610 ;
        RECT -155.205 -87.870 -154.945 -87.610 ;
        RECT -145.745 -87.870 -145.485 -87.610 ;
        RECT -145.285 -87.870 -145.025 -87.610 ;
        RECT -135.825 -87.870 -135.565 -87.610 ;
        RECT -135.365 -87.870 -135.105 -87.610 ;
        RECT -125.905 -87.870 -125.645 -87.610 ;
        RECT -125.445 -87.870 -125.185 -87.610 ;
        RECT -115.985 -87.870 -115.725 -87.610 ;
        RECT -115.525 -87.870 -115.265 -87.610 ;
        RECT -106.065 -87.870 -105.805 -87.610 ;
        RECT -105.605 -87.870 -105.345 -87.610 ;
        RECT -96.145 -87.870 -95.885 -87.610 ;
        RECT -95.685 -87.870 -95.425 -87.610 ;
        RECT -86.225 -87.870 -85.965 -87.610 ;
        RECT -85.765 -87.870 -85.505 -87.610 ;
        RECT -76.305 -87.870 -76.045 -87.610 ;
        RECT -75.845 -87.870 -75.585 -87.610 ;
        RECT -66.385 -87.870 -66.125 -87.610 ;
        RECT -65.925 -87.870 -65.665 -87.610 ;
        RECT -56.465 -87.870 -56.205 -87.610 ;
        RECT -56.005 -87.870 -55.745 -87.610 ;
        RECT -46.545 -87.870 -46.285 -87.610 ;
        RECT -46.085 -87.870 -45.825 -87.610 ;
        RECT -36.625 -87.870 -36.365 -87.610 ;
        RECT -36.165 -87.870 -35.905 -87.610 ;
        RECT -26.705 -87.870 -26.445 -87.610 ;
        RECT -26.245 -87.870 -25.985 -87.610 ;
        RECT -16.785 -87.870 -16.525 -87.610 ;
        RECT -16.325 -87.870 -16.065 -87.610 ;
        RECT -6.865 -87.870 -6.605 -87.610 ;
        RECT -6.405 -87.870 -6.145 -87.610 ;
        RECT 3.055 -87.870 3.315 -87.610 ;
        RECT 3.515 -87.870 3.775 -87.610 ;
        RECT 12.975 -87.870 13.235 -87.610 ;
        RECT 13.435 -87.870 13.695 -87.610 ;
        RECT 22.895 -87.870 23.155 -87.610 ;
        RECT 23.355 -87.870 23.615 -87.610 ;
        RECT -279.665 -90.580 -279.405 -90.320 ;
        RECT -279.205 -90.580 -278.945 -90.320 ;
        RECT -269.745 -90.580 -269.485 -90.320 ;
        RECT -269.285 -90.580 -269.025 -90.320 ;
        RECT -259.825 -90.580 -259.565 -90.320 ;
        RECT -259.365 -90.580 -259.105 -90.320 ;
        RECT -249.905 -90.580 -249.645 -90.320 ;
        RECT -249.445 -90.580 -249.185 -90.320 ;
        RECT -239.985 -90.580 -239.725 -90.320 ;
        RECT -239.525 -90.580 -239.265 -90.320 ;
        RECT -230.065 -90.580 -229.805 -90.320 ;
        RECT -229.605 -90.580 -229.345 -90.320 ;
        RECT -220.145 -90.580 -219.885 -90.320 ;
        RECT -219.685 -90.580 -219.425 -90.320 ;
        RECT -210.225 -90.580 -209.965 -90.320 ;
        RECT -209.765 -90.580 -209.505 -90.320 ;
        RECT -200.305 -90.580 -200.045 -90.320 ;
        RECT -199.845 -90.580 -199.585 -90.320 ;
        RECT -190.385 -90.580 -190.125 -90.320 ;
        RECT -189.925 -90.580 -189.665 -90.320 ;
        RECT -180.465 -90.580 -180.205 -90.320 ;
        RECT -180.005 -90.580 -179.745 -90.320 ;
        RECT -170.545 -90.580 -170.285 -90.320 ;
        RECT -170.085 -90.580 -169.825 -90.320 ;
        RECT -160.625 -90.580 -160.365 -90.320 ;
        RECT -160.165 -90.580 -159.905 -90.320 ;
        RECT -150.705 -90.580 -150.445 -90.320 ;
        RECT -150.245 -90.580 -149.985 -90.320 ;
        RECT -140.785 -90.580 -140.525 -90.320 ;
        RECT -140.325 -90.580 -140.065 -90.320 ;
        RECT -130.865 -90.580 -130.605 -90.320 ;
        RECT -130.405 -90.580 -130.145 -90.320 ;
        RECT -120.945 -90.580 -120.685 -90.320 ;
        RECT -120.485 -90.580 -120.225 -90.320 ;
        RECT -111.025 -90.580 -110.765 -90.320 ;
        RECT -110.565 -90.580 -110.305 -90.320 ;
        RECT -101.105 -90.580 -100.845 -90.320 ;
        RECT -100.645 -90.580 -100.385 -90.320 ;
        RECT -91.185 -90.580 -90.925 -90.320 ;
        RECT -90.725 -90.580 -90.465 -90.320 ;
        RECT -81.265 -90.580 -81.005 -90.320 ;
        RECT -80.805 -90.580 -80.545 -90.320 ;
        RECT -71.345 -90.580 -71.085 -90.320 ;
        RECT -70.885 -90.580 -70.625 -90.320 ;
        RECT -61.425 -90.580 -61.165 -90.320 ;
        RECT -60.965 -90.580 -60.705 -90.320 ;
        RECT -51.505 -90.580 -51.245 -90.320 ;
        RECT -51.045 -90.580 -50.785 -90.320 ;
        RECT -41.585 -90.580 -41.325 -90.320 ;
        RECT -41.125 -90.580 -40.865 -90.320 ;
        RECT -31.665 -90.580 -31.405 -90.320 ;
        RECT -31.205 -90.580 -30.945 -90.320 ;
        RECT -21.745 -90.580 -21.485 -90.320 ;
        RECT -21.285 -90.580 -21.025 -90.320 ;
        RECT -11.825 -90.580 -11.565 -90.320 ;
        RECT -11.365 -90.580 -11.105 -90.320 ;
        RECT -1.905 -90.580 -1.645 -90.320 ;
        RECT -1.445 -90.580 -1.185 -90.320 ;
        RECT 8.015 -90.580 8.275 -90.320 ;
        RECT 8.475 -90.580 8.735 -90.320 ;
        RECT 17.935 -90.580 18.195 -90.320 ;
        RECT 18.395 -90.580 18.655 -90.320 ;
        RECT 27.855 -90.580 28.115 -90.320 ;
        RECT -284.855 -92.170 -284.595 -91.910 ;
        RECT -283.925 -92.170 -283.665 -91.910 ;
        RECT -274.935 -92.170 -274.675 -91.910 ;
        RECT -274.005 -92.170 -273.745 -91.910 ;
        RECT -265.015 -92.170 -264.755 -91.910 ;
        RECT -264.085 -92.170 -263.825 -91.910 ;
        RECT -255.095 -92.170 -254.835 -91.910 ;
        RECT -254.165 -92.170 -253.905 -91.910 ;
        RECT -245.175 -92.170 -244.915 -91.910 ;
        RECT -244.245 -92.170 -243.985 -91.910 ;
        RECT -235.255 -92.170 -234.995 -91.910 ;
        RECT -234.325 -92.170 -234.065 -91.910 ;
        RECT -225.335 -92.170 -225.075 -91.910 ;
        RECT -224.405 -92.170 -224.145 -91.910 ;
        RECT -215.415 -92.170 -215.155 -91.910 ;
        RECT -214.485 -92.170 -214.225 -91.910 ;
        RECT -205.495 -92.170 -205.235 -91.910 ;
        RECT -204.565 -92.170 -204.305 -91.910 ;
        RECT -195.575 -92.170 -195.315 -91.910 ;
        RECT -194.645 -92.170 -194.385 -91.910 ;
        RECT -185.655 -92.170 -185.395 -91.910 ;
        RECT -184.725 -92.170 -184.465 -91.910 ;
        RECT -175.735 -92.170 -175.475 -91.910 ;
        RECT -174.805 -92.170 -174.545 -91.910 ;
        RECT -165.815 -92.170 -165.555 -91.910 ;
        RECT -164.885 -92.170 -164.625 -91.910 ;
        RECT -155.895 -92.170 -155.635 -91.910 ;
        RECT -154.965 -92.170 -154.705 -91.910 ;
        RECT -145.975 -92.170 -145.715 -91.910 ;
        RECT -145.045 -92.170 -144.785 -91.910 ;
        RECT -136.055 -92.170 -135.795 -91.910 ;
        RECT -135.125 -92.170 -134.865 -91.910 ;
        RECT -126.135 -92.170 -125.875 -91.910 ;
        RECT -125.205 -92.170 -124.945 -91.910 ;
        RECT -116.215 -92.170 -115.955 -91.910 ;
        RECT -115.285 -92.170 -115.025 -91.910 ;
        RECT -106.295 -92.170 -106.035 -91.910 ;
        RECT -105.365 -92.170 -105.105 -91.910 ;
        RECT -96.375 -92.170 -96.115 -91.910 ;
        RECT -95.445 -92.170 -95.185 -91.910 ;
        RECT -86.455 -92.170 -86.195 -91.910 ;
        RECT -85.525 -92.170 -85.265 -91.910 ;
        RECT -76.535 -92.170 -76.275 -91.910 ;
        RECT -75.605 -92.170 -75.345 -91.910 ;
        RECT -66.615 -92.170 -66.355 -91.910 ;
        RECT -65.685 -92.170 -65.425 -91.910 ;
        RECT -56.695 -92.170 -56.435 -91.910 ;
        RECT -55.765 -92.170 -55.505 -91.910 ;
        RECT -46.775 -92.170 -46.515 -91.910 ;
        RECT -45.845 -92.170 -45.585 -91.910 ;
        RECT -36.855 -92.170 -36.595 -91.910 ;
        RECT -35.925 -92.170 -35.665 -91.910 ;
        RECT -26.935 -92.170 -26.675 -91.910 ;
        RECT -26.005 -92.170 -25.745 -91.910 ;
        RECT -17.015 -92.170 -16.755 -91.910 ;
        RECT -16.085 -92.170 -15.825 -91.910 ;
        RECT -7.095 -92.170 -6.835 -91.910 ;
        RECT -6.165 -92.170 -5.905 -91.910 ;
        RECT 2.825 -92.170 3.085 -91.910 ;
        RECT 3.755 -92.170 4.015 -91.910 ;
        RECT 12.745 -92.170 13.005 -91.910 ;
        RECT 13.675 -92.170 13.935 -91.910 ;
        RECT 22.665 -92.170 22.925 -91.910 ;
        RECT 23.595 -92.170 23.855 -91.910 ;
        RECT -279.655 -173.990 -279.395 -173.730 ;
        RECT -278.715 -174.000 -278.455 -173.740 ;
        RECT -269.025 -173.995 -268.765 -173.735 ;
        RECT -259.815 -173.990 -259.555 -173.730 ;
        RECT -258.875 -174.000 -258.615 -173.740 ;
        RECT -249.895 -173.990 -249.635 -173.730 ;
        RECT -248.955 -174.000 -248.695 -173.740 ;
        RECT -239.975 -173.990 -239.715 -173.730 ;
        RECT -239.035 -174.000 -238.775 -173.740 ;
        RECT -230.055 -173.990 -229.795 -173.730 ;
        RECT -229.115 -174.000 -228.855 -173.740 ;
        RECT -220.135 -173.990 -219.875 -173.730 ;
        RECT -219.195 -174.000 -218.935 -173.740 ;
        RECT -210.215 -173.990 -209.955 -173.730 ;
        RECT -209.275 -174.000 -209.015 -173.740 ;
        RECT -200.295 -173.990 -200.035 -173.730 ;
        RECT -199.355 -174.000 -199.095 -173.740 ;
        RECT -190.375 -173.990 -190.115 -173.730 ;
        RECT -189.435 -174.000 -189.175 -173.740 ;
        RECT -180.455 -173.990 -180.195 -173.730 ;
        RECT -179.515 -174.000 -179.255 -173.740 ;
        RECT -170.535 -173.990 -170.275 -173.730 ;
        RECT -169.595 -174.000 -169.335 -173.740 ;
        RECT -160.615 -173.990 -160.355 -173.730 ;
        RECT -159.675 -174.000 -159.415 -173.740 ;
        RECT -150.695 -173.990 -150.435 -173.730 ;
        RECT -149.755 -174.000 -149.495 -173.740 ;
        RECT -140.775 -173.990 -140.515 -173.730 ;
        RECT -139.835 -174.000 -139.575 -173.740 ;
        RECT -130.855 -173.990 -130.595 -173.730 ;
        RECT -129.915 -174.000 -129.655 -173.740 ;
        RECT -120.935 -173.990 -120.675 -173.730 ;
        RECT -119.995 -174.000 -119.735 -173.740 ;
        RECT -111.015 -173.990 -110.755 -173.730 ;
        RECT -110.075 -174.000 -109.815 -173.740 ;
        RECT -101.095 -173.990 -100.835 -173.730 ;
        RECT -100.155 -174.000 -99.895 -173.740 ;
        RECT -91.175 -173.990 -90.915 -173.730 ;
        RECT -90.235 -174.000 -89.975 -173.740 ;
        RECT -81.255 -173.990 -80.995 -173.730 ;
        RECT -80.315 -174.000 -80.055 -173.740 ;
        RECT -71.335 -173.990 -71.075 -173.730 ;
        RECT -70.395 -174.000 -70.135 -173.740 ;
        RECT -61.415 -173.990 -61.155 -173.730 ;
        RECT -60.475 -174.000 -60.215 -173.740 ;
        RECT -51.495 -173.990 -51.235 -173.730 ;
        RECT -50.555 -174.000 -50.295 -173.740 ;
        RECT -41.575 -173.990 -41.315 -173.730 ;
        RECT -40.635 -174.000 -40.375 -173.740 ;
        RECT -31.655 -173.990 -31.395 -173.730 ;
        RECT -30.715 -174.000 -30.455 -173.740 ;
        RECT -21.735 -173.990 -21.475 -173.730 ;
        RECT -20.795 -174.000 -20.535 -173.740 ;
        RECT -11.815 -173.990 -11.555 -173.730 ;
        RECT -10.875 -174.000 -10.615 -173.740 ;
        RECT -1.895 -173.990 -1.635 -173.730 ;
        RECT -0.955 -174.000 -0.695 -173.740 ;
        RECT 8.025 -173.990 8.285 -173.730 ;
        RECT 8.965 -174.000 9.225 -173.740 ;
        RECT 17.945 -173.990 18.205 -173.730 ;
        RECT 18.885 -174.000 19.145 -173.740 ;
        RECT 27.865 -173.990 28.125 -173.730 ;
        RECT -284.375 -175.580 -284.115 -175.320 ;
        RECT -283.915 -175.580 -283.655 -175.320 ;
        RECT -274.455 -175.580 -274.195 -175.320 ;
        RECT -273.995 -175.580 -273.735 -175.320 ;
        RECT -264.535 -175.580 -264.275 -175.320 ;
        RECT -264.075 -175.580 -263.815 -175.320 ;
        RECT -254.615 -175.580 -254.355 -175.320 ;
        RECT -254.155 -175.580 -253.895 -175.320 ;
        RECT -244.695 -175.580 -244.435 -175.320 ;
        RECT -244.235 -175.580 -243.975 -175.320 ;
        RECT -234.775 -175.580 -234.515 -175.320 ;
        RECT -234.315 -175.580 -234.055 -175.320 ;
        RECT -224.855 -175.580 -224.595 -175.320 ;
        RECT -224.395 -175.580 -224.135 -175.320 ;
        RECT -214.935 -175.580 -214.675 -175.320 ;
        RECT -214.475 -175.580 -214.215 -175.320 ;
        RECT -205.015 -175.580 -204.755 -175.320 ;
        RECT -204.555 -175.580 -204.295 -175.320 ;
        RECT -195.095 -175.580 -194.835 -175.320 ;
        RECT -194.635 -175.580 -194.375 -175.320 ;
        RECT -185.175 -175.580 -184.915 -175.320 ;
        RECT -184.715 -175.580 -184.455 -175.320 ;
        RECT -175.255 -175.580 -174.995 -175.320 ;
        RECT -174.795 -175.580 -174.535 -175.320 ;
        RECT -165.335 -175.580 -165.075 -175.320 ;
        RECT -164.875 -175.580 -164.615 -175.320 ;
        RECT -155.415 -175.580 -155.155 -175.320 ;
        RECT -154.955 -175.580 -154.695 -175.320 ;
        RECT -145.495 -175.580 -145.235 -175.320 ;
        RECT -145.035 -175.580 -144.775 -175.320 ;
        RECT -135.575 -175.580 -135.315 -175.320 ;
        RECT -135.115 -175.580 -134.855 -175.320 ;
        RECT -125.655 -175.580 -125.395 -175.320 ;
        RECT -125.195 -175.580 -124.935 -175.320 ;
        RECT -115.735 -175.580 -115.475 -175.320 ;
        RECT -115.275 -175.580 -115.015 -175.320 ;
        RECT -105.815 -175.580 -105.555 -175.320 ;
        RECT -105.355 -175.580 -105.095 -175.320 ;
        RECT -95.895 -175.580 -95.635 -175.320 ;
        RECT -95.435 -175.580 -95.175 -175.320 ;
        RECT -85.975 -175.580 -85.715 -175.320 ;
        RECT -85.515 -175.580 -85.255 -175.320 ;
        RECT -76.055 -175.580 -75.795 -175.320 ;
        RECT -75.595 -175.580 -75.335 -175.320 ;
        RECT -66.135 -175.580 -65.875 -175.320 ;
        RECT -65.675 -175.580 -65.415 -175.320 ;
        RECT -56.215 -175.580 -55.955 -175.320 ;
        RECT -55.755 -175.580 -55.495 -175.320 ;
        RECT -46.295 -175.580 -46.035 -175.320 ;
        RECT -45.835 -175.580 -45.575 -175.320 ;
        RECT -36.375 -175.580 -36.115 -175.320 ;
        RECT -35.915 -175.580 -35.655 -175.320 ;
        RECT -26.455 -175.580 -26.195 -175.320 ;
        RECT -25.995 -175.580 -25.735 -175.320 ;
        RECT -16.535 -175.580 -16.275 -175.320 ;
        RECT -16.075 -175.580 -15.815 -175.320 ;
        RECT -6.615 -175.580 -6.355 -175.320 ;
        RECT -6.155 -175.580 -5.895 -175.320 ;
        RECT 3.305 -175.580 3.565 -175.320 ;
        RECT 3.765 -175.580 4.025 -175.320 ;
        RECT 13.225 -175.580 13.485 -175.320 ;
        RECT 13.685 -175.580 13.945 -175.320 ;
        RECT 23.145 -175.580 23.405 -175.320 ;
        RECT 23.605 -175.580 23.865 -175.320 ;
        RECT -279.415 -178.290 -279.155 -178.030 ;
        RECT -278.955 -178.290 -278.695 -178.030 ;
        RECT -269.495 -178.290 -269.235 -178.030 ;
        RECT -269.035 -178.290 -268.775 -178.030 ;
        RECT -259.575 -178.290 -259.315 -178.030 ;
        RECT -259.115 -178.290 -258.855 -178.030 ;
        RECT -249.655 -178.290 -249.395 -178.030 ;
        RECT -249.195 -178.290 -248.935 -178.030 ;
        RECT -239.735 -178.290 -239.475 -178.030 ;
        RECT -239.275 -178.290 -239.015 -178.030 ;
        RECT -229.815 -178.290 -229.555 -178.030 ;
        RECT -229.355 -178.290 -229.095 -178.030 ;
        RECT -219.895 -178.290 -219.635 -178.030 ;
        RECT -219.435 -178.290 -219.175 -178.030 ;
        RECT -209.975 -178.290 -209.715 -178.030 ;
        RECT -209.515 -178.290 -209.255 -178.030 ;
        RECT -200.055 -178.290 -199.795 -178.030 ;
        RECT -199.595 -178.290 -199.335 -178.030 ;
        RECT -190.135 -178.290 -189.875 -178.030 ;
        RECT -189.675 -178.290 -189.415 -178.030 ;
        RECT -180.215 -178.290 -179.955 -178.030 ;
        RECT -179.755 -178.290 -179.495 -178.030 ;
        RECT -170.295 -178.290 -170.035 -178.030 ;
        RECT -169.835 -178.290 -169.575 -178.030 ;
        RECT -160.375 -178.290 -160.115 -178.030 ;
        RECT -159.915 -178.290 -159.655 -178.030 ;
        RECT -150.455 -178.290 -150.195 -178.030 ;
        RECT -149.995 -178.290 -149.735 -178.030 ;
        RECT -140.535 -178.290 -140.275 -178.030 ;
        RECT -140.075 -178.290 -139.815 -178.030 ;
        RECT -130.615 -178.290 -130.355 -178.030 ;
        RECT -130.155 -178.290 -129.895 -178.030 ;
        RECT -120.695 -178.290 -120.435 -178.030 ;
        RECT -120.235 -178.290 -119.975 -178.030 ;
        RECT -110.775 -178.290 -110.515 -178.030 ;
        RECT -110.315 -178.290 -110.055 -178.030 ;
        RECT -100.855 -178.290 -100.595 -178.030 ;
        RECT -100.395 -178.290 -100.135 -178.030 ;
        RECT -90.935 -178.290 -90.675 -178.030 ;
        RECT -90.475 -178.290 -90.215 -178.030 ;
        RECT -81.015 -178.290 -80.755 -178.030 ;
        RECT -80.555 -178.290 -80.295 -178.030 ;
        RECT -71.095 -178.290 -70.835 -178.030 ;
        RECT -70.635 -178.290 -70.375 -178.030 ;
        RECT -61.175 -178.290 -60.915 -178.030 ;
        RECT -60.715 -178.290 -60.455 -178.030 ;
        RECT -51.255 -178.290 -50.995 -178.030 ;
        RECT -50.795 -178.290 -50.535 -178.030 ;
        RECT -41.335 -178.290 -41.075 -178.030 ;
        RECT -40.875 -178.290 -40.615 -178.030 ;
        RECT -31.415 -178.290 -31.155 -178.030 ;
        RECT -30.955 -178.290 -30.695 -178.030 ;
        RECT -21.495 -178.290 -21.235 -178.030 ;
        RECT -21.035 -178.290 -20.775 -178.030 ;
        RECT -11.575 -178.290 -11.315 -178.030 ;
        RECT -11.115 -178.290 -10.855 -178.030 ;
        RECT -1.655 -178.290 -1.395 -178.030 ;
        RECT -1.195 -178.290 -0.935 -178.030 ;
        RECT 8.265 -178.290 8.525 -178.030 ;
        RECT 8.725 -178.290 8.985 -178.030 ;
        RECT 18.185 -178.290 18.445 -178.030 ;
        RECT 18.645 -178.290 18.905 -178.030 ;
        RECT 28.105 -178.290 28.365 -178.030 ;
        RECT -284.605 -179.880 -284.345 -179.620 ;
        RECT -283.675 -179.880 -283.415 -179.620 ;
        RECT -274.685 -179.880 -274.425 -179.620 ;
        RECT -273.755 -179.880 -273.495 -179.620 ;
        RECT -264.765 -179.880 -264.505 -179.620 ;
        RECT -263.835 -179.880 -263.575 -179.620 ;
        RECT -254.845 -179.880 -254.585 -179.620 ;
        RECT -253.915 -179.880 -253.655 -179.620 ;
        RECT -244.925 -179.880 -244.665 -179.620 ;
        RECT -243.995 -179.880 -243.735 -179.620 ;
        RECT -235.005 -179.880 -234.745 -179.620 ;
        RECT -234.075 -179.880 -233.815 -179.620 ;
        RECT -225.085 -179.880 -224.825 -179.620 ;
        RECT -224.155 -179.880 -223.895 -179.620 ;
        RECT -215.165 -179.880 -214.905 -179.620 ;
        RECT -214.235 -179.880 -213.975 -179.620 ;
        RECT -205.245 -179.880 -204.985 -179.620 ;
        RECT -204.315 -179.880 -204.055 -179.620 ;
        RECT -195.325 -179.880 -195.065 -179.620 ;
        RECT -194.395 -179.880 -194.135 -179.620 ;
        RECT -185.405 -179.880 -185.145 -179.620 ;
        RECT -184.475 -179.880 -184.215 -179.620 ;
        RECT -175.485 -179.880 -175.225 -179.620 ;
        RECT -174.555 -179.880 -174.295 -179.620 ;
        RECT -165.565 -179.880 -165.305 -179.620 ;
        RECT -164.635 -179.880 -164.375 -179.620 ;
        RECT -155.645 -179.880 -155.385 -179.620 ;
        RECT -154.715 -179.880 -154.455 -179.620 ;
        RECT -145.725 -179.880 -145.465 -179.620 ;
        RECT -144.795 -179.880 -144.535 -179.620 ;
        RECT -135.805 -179.880 -135.545 -179.620 ;
        RECT -134.875 -179.880 -134.615 -179.620 ;
        RECT -125.885 -179.880 -125.625 -179.620 ;
        RECT -124.955 -179.880 -124.695 -179.620 ;
        RECT -115.965 -179.880 -115.705 -179.620 ;
        RECT -115.035 -179.880 -114.775 -179.620 ;
        RECT -106.045 -179.880 -105.785 -179.620 ;
        RECT -105.115 -179.880 -104.855 -179.620 ;
        RECT -96.125 -179.880 -95.865 -179.620 ;
        RECT -95.195 -179.880 -94.935 -179.620 ;
        RECT -86.205 -179.880 -85.945 -179.620 ;
        RECT -85.275 -179.880 -85.015 -179.620 ;
        RECT -76.285 -179.880 -76.025 -179.620 ;
        RECT -75.355 -179.880 -75.095 -179.620 ;
        RECT -66.365 -179.880 -66.105 -179.620 ;
        RECT -65.435 -179.880 -65.175 -179.620 ;
        RECT -56.445 -179.880 -56.185 -179.620 ;
        RECT -55.515 -179.880 -55.255 -179.620 ;
        RECT -46.525 -179.880 -46.265 -179.620 ;
        RECT -45.595 -179.880 -45.335 -179.620 ;
        RECT -36.605 -179.880 -36.345 -179.620 ;
        RECT -35.675 -179.880 -35.415 -179.620 ;
        RECT -26.685 -179.880 -26.425 -179.620 ;
        RECT -25.755 -179.880 -25.495 -179.620 ;
        RECT -16.765 -179.880 -16.505 -179.620 ;
        RECT -15.835 -179.880 -15.575 -179.620 ;
        RECT -6.845 -179.880 -6.585 -179.620 ;
        RECT -5.915 -179.880 -5.655 -179.620 ;
        RECT 3.075 -179.880 3.335 -179.620 ;
        RECT 4.005 -179.880 4.265 -179.620 ;
        RECT 12.995 -179.880 13.255 -179.620 ;
        RECT 13.925 -179.880 14.185 -179.620 ;
        RECT 22.915 -179.880 23.175 -179.620 ;
        RECT 23.845 -179.880 24.105 -179.620 ;
      LAYER met2 ;
        RECT -282.020 94.730 -280.600 95.140 ;
        RECT -272.100 94.730 -270.680 95.140 ;
        RECT -262.180 94.730 -260.760 95.140 ;
        RECT -252.260 94.730 -250.840 95.140 ;
        RECT -242.340 94.730 -240.920 95.140 ;
        RECT -232.420 94.730 -231.000 95.140 ;
        RECT -222.500 94.730 -221.080 95.140 ;
        RECT -212.580 94.730 -211.160 95.140 ;
        RECT -202.660 94.730 -201.240 95.140 ;
        RECT -192.740 94.730 -191.320 95.140 ;
        RECT -182.820 94.730 -181.400 95.140 ;
        RECT -172.900 94.730 -171.480 95.140 ;
        RECT -162.980 94.730 -161.560 95.140 ;
        RECT -153.060 94.730 -151.640 95.140 ;
        RECT -143.140 94.730 -141.720 95.140 ;
        RECT -133.220 94.730 -131.800 95.140 ;
        RECT -123.300 94.730 -121.880 95.140 ;
        RECT -113.380 94.730 -111.960 95.140 ;
        RECT -103.460 94.730 -102.040 95.140 ;
        RECT -93.540 94.730 -92.120 95.140 ;
        RECT -83.620 94.730 -82.200 95.140 ;
        RECT -73.700 94.730 -72.280 95.140 ;
        RECT -63.780 94.730 -62.360 95.140 ;
        RECT -53.860 94.730 -52.440 95.140 ;
        RECT -43.940 94.730 -42.520 95.140 ;
        RECT -34.020 94.730 -32.600 95.140 ;
        RECT -24.100 94.730 -22.680 95.140 ;
        RECT -14.180 94.730 -12.760 95.140 ;
        RECT -4.260 94.730 -2.840 95.140 ;
        RECT 5.660 94.730 7.080 95.140 ;
        RECT 15.580 94.730 17.000 95.140 ;
        RECT 25.500 94.730 26.440 95.140 ;
        RECT -272.100 94.360 -270.690 94.730 ;
        RECT -286.870 93.090 -285.670 93.570 ;
        RECT -276.950 93.090 -275.750 93.570 ;
        RECT -267.030 93.090 -265.830 93.570 ;
        RECT -257.110 93.090 -255.910 93.570 ;
        RECT -247.190 93.090 -245.990 93.570 ;
        RECT -237.270 93.090 -236.070 93.570 ;
        RECT -227.350 93.090 -226.150 93.570 ;
        RECT -217.430 93.090 -216.230 93.570 ;
        RECT -207.510 93.090 -206.310 93.570 ;
        RECT -197.590 93.090 -196.390 93.570 ;
        RECT -187.670 93.090 -186.470 93.570 ;
        RECT -177.750 93.090 -176.550 93.570 ;
        RECT -167.830 93.090 -166.630 93.570 ;
        RECT -157.910 93.090 -156.710 93.570 ;
        RECT -147.990 93.090 -146.790 93.570 ;
        RECT -138.070 93.090 -136.870 93.570 ;
        RECT -128.150 93.090 -126.950 93.570 ;
        RECT -118.230 93.090 -117.030 93.570 ;
        RECT -108.310 93.090 -107.110 93.570 ;
        RECT -98.390 93.090 -97.190 93.570 ;
        RECT -88.470 93.090 -87.270 93.570 ;
        RECT -78.550 93.090 -77.350 93.570 ;
        RECT -68.630 93.090 -67.430 93.570 ;
        RECT -58.710 93.090 -57.510 93.570 ;
        RECT -48.790 93.090 -47.590 93.570 ;
        RECT -38.870 93.090 -37.670 93.570 ;
        RECT -28.950 93.090 -27.750 93.570 ;
        RECT -19.030 93.090 -17.830 93.570 ;
        RECT -9.110 93.090 -7.910 93.570 ;
        RECT 0.810 93.090 2.010 93.570 ;
        RECT 10.730 93.090 11.930 93.570 ;
        RECT 20.650 93.090 21.850 93.570 ;
        RECT -281.910 90.370 -280.710 90.850 ;
        RECT -271.990 90.370 -270.790 90.850 ;
        RECT -262.070 90.370 -260.870 90.850 ;
        RECT -252.150 90.370 -250.950 90.850 ;
        RECT -242.230 90.370 -241.030 90.850 ;
        RECT -232.310 90.370 -231.110 90.850 ;
        RECT -222.390 90.370 -221.190 90.850 ;
        RECT -212.470 90.370 -211.270 90.850 ;
        RECT -202.550 90.370 -201.350 90.850 ;
        RECT -192.630 90.370 -191.430 90.850 ;
        RECT -182.710 90.370 -181.510 90.850 ;
        RECT -172.790 90.370 -171.590 90.850 ;
        RECT -162.870 90.370 -161.670 90.850 ;
        RECT -152.950 90.370 -151.750 90.850 ;
        RECT -143.030 90.370 -141.830 90.850 ;
        RECT -133.110 90.370 -131.910 90.850 ;
        RECT -123.190 90.370 -121.990 90.850 ;
        RECT -113.270 90.370 -112.070 90.850 ;
        RECT -103.350 90.370 -102.150 90.850 ;
        RECT -93.430 90.370 -92.230 90.850 ;
        RECT -83.510 90.370 -82.310 90.850 ;
        RECT -73.590 90.370 -72.390 90.850 ;
        RECT -63.670 90.370 -62.470 90.850 ;
        RECT -53.750 90.370 -52.550 90.850 ;
        RECT -43.830 90.370 -42.630 90.850 ;
        RECT -33.910 90.370 -32.710 90.850 ;
        RECT -23.990 90.370 -22.790 90.850 ;
        RECT -14.070 90.370 -12.870 90.850 ;
        RECT -4.150 90.370 -2.950 90.850 ;
        RECT 5.770 90.370 6.970 90.850 ;
        RECT 15.690 90.370 16.890 90.850 ;
        RECT 25.610 90.370 26.440 90.850 ;
        RECT -286.980 88.800 -285.560 89.210 ;
        RECT -277.060 88.800 -275.640 89.210 ;
        RECT -267.140 88.800 -265.720 89.210 ;
        RECT -257.220 88.800 -255.800 89.210 ;
        RECT -247.300 88.800 -245.880 89.210 ;
        RECT -237.380 88.800 -235.960 89.210 ;
        RECT -227.460 88.800 -226.040 89.210 ;
        RECT -217.540 88.800 -216.120 89.210 ;
        RECT -207.620 88.800 -206.200 89.210 ;
        RECT -197.700 88.800 -196.280 89.210 ;
        RECT -187.780 88.800 -186.360 89.210 ;
        RECT -177.860 88.800 -176.440 89.210 ;
        RECT -167.940 88.800 -166.520 89.210 ;
        RECT -158.020 88.800 -156.600 89.210 ;
        RECT -148.100 88.800 -146.680 89.210 ;
        RECT -138.180 88.800 -136.760 89.210 ;
        RECT -128.260 88.800 -126.840 89.210 ;
        RECT -118.340 88.800 -116.920 89.210 ;
        RECT -108.420 88.800 -107.000 89.210 ;
        RECT -98.500 88.800 -97.080 89.210 ;
        RECT -88.580 88.800 -87.160 89.210 ;
        RECT -78.660 88.800 -77.240 89.210 ;
        RECT -68.740 88.800 -67.320 89.210 ;
        RECT -58.820 88.800 -57.400 89.210 ;
        RECT -48.900 88.800 -47.480 89.210 ;
        RECT -38.980 88.800 -37.560 89.210 ;
        RECT -29.060 88.800 -27.640 89.210 ;
        RECT -19.140 88.800 -17.720 89.210 ;
        RECT -9.220 88.800 -7.800 89.210 ;
        RECT 0.700 88.800 2.120 89.210 ;
        RECT 10.620 88.800 12.040 89.210 ;
        RECT 20.540 88.800 21.960 89.210 ;
        RECT -281.770 7.020 -280.350 7.430 ;
        RECT -271.850 7.020 -270.430 7.430 ;
        RECT -261.930 7.020 -260.510 7.430 ;
        RECT -252.010 7.020 -250.590 7.430 ;
        RECT -242.090 7.020 -240.670 7.430 ;
        RECT -232.170 7.020 -230.750 7.430 ;
        RECT -222.250 7.020 -220.830 7.430 ;
        RECT -212.330 7.020 -210.910 7.430 ;
        RECT -202.410 7.020 -200.990 7.430 ;
        RECT -192.490 7.020 -191.070 7.430 ;
        RECT -182.570 7.020 -181.150 7.430 ;
        RECT -172.650 7.020 -171.230 7.430 ;
        RECT -162.730 7.020 -161.310 7.430 ;
        RECT -152.810 7.020 -151.390 7.430 ;
        RECT -142.890 7.020 -141.470 7.430 ;
        RECT -132.970 7.020 -131.550 7.430 ;
        RECT -123.050 7.020 -121.630 7.430 ;
        RECT -113.130 7.020 -111.710 7.430 ;
        RECT -103.210 7.020 -101.790 7.430 ;
        RECT -93.290 7.020 -91.870 7.430 ;
        RECT -83.370 7.020 -81.950 7.430 ;
        RECT -73.450 7.020 -72.030 7.430 ;
        RECT -63.530 7.020 -62.110 7.430 ;
        RECT -53.610 7.020 -52.190 7.430 ;
        RECT -43.690 7.020 -42.270 7.430 ;
        RECT -33.770 7.020 -32.350 7.430 ;
        RECT -23.850 7.020 -22.430 7.430 ;
        RECT -13.930 7.020 -12.510 7.430 ;
        RECT -4.010 7.020 -2.590 7.430 ;
        RECT 5.910 7.020 7.330 7.430 ;
        RECT 15.830 7.020 17.250 7.430 ;
        RECT 25.750 7.020 26.690 7.430 ;
        RECT -271.850 6.650 -270.440 7.020 ;
        RECT -286.620 5.380 -285.420 5.860 ;
        RECT -276.700 5.380 -275.500 5.860 ;
        RECT -266.780 5.380 -265.580 5.860 ;
        RECT -256.860 5.380 -255.660 5.860 ;
        RECT -246.940 5.380 -245.740 5.860 ;
        RECT -237.020 5.380 -235.820 5.860 ;
        RECT -227.100 5.380 -225.900 5.860 ;
        RECT -217.180 5.380 -215.980 5.860 ;
        RECT -207.260 5.380 -206.060 5.860 ;
        RECT -197.340 5.380 -196.140 5.860 ;
        RECT -187.420 5.380 -186.220 5.860 ;
        RECT -177.500 5.380 -176.300 5.860 ;
        RECT -167.580 5.380 -166.380 5.860 ;
        RECT -157.660 5.380 -156.460 5.860 ;
        RECT -147.740 5.380 -146.540 5.860 ;
        RECT -137.820 5.380 -136.620 5.860 ;
        RECT -127.900 5.380 -126.700 5.860 ;
        RECT -117.980 5.380 -116.780 5.860 ;
        RECT -108.060 5.380 -106.860 5.860 ;
        RECT -98.140 5.380 -96.940 5.860 ;
        RECT -88.220 5.380 -87.020 5.860 ;
        RECT -78.300 5.380 -77.100 5.860 ;
        RECT -68.380 5.380 -67.180 5.860 ;
        RECT -58.460 5.380 -57.260 5.860 ;
        RECT -48.540 5.380 -47.340 5.860 ;
        RECT -38.620 5.380 -37.420 5.860 ;
        RECT -28.700 5.380 -27.500 5.860 ;
        RECT -18.780 5.380 -17.580 5.860 ;
        RECT -8.860 5.380 -7.660 5.860 ;
        RECT 1.060 5.380 2.260 5.860 ;
        RECT 10.980 5.380 12.180 5.860 ;
        RECT 20.900 5.380 22.100 5.860 ;
        RECT -281.660 2.660 -280.460 3.140 ;
        RECT -271.740 2.660 -270.540 3.140 ;
        RECT -261.820 2.660 -260.620 3.140 ;
        RECT -251.900 2.660 -250.700 3.140 ;
        RECT -241.980 2.660 -240.780 3.140 ;
        RECT -232.060 2.660 -230.860 3.140 ;
        RECT -222.140 2.660 -220.940 3.140 ;
        RECT -212.220 2.660 -211.020 3.140 ;
        RECT -202.300 2.660 -201.100 3.140 ;
        RECT -192.380 2.660 -191.180 3.140 ;
        RECT -182.460 2.660 -181.260 3.140 ;
        RECT -172.540 2.660 -171.340 3.140 ;
        RECT -162.620 2.660 -161.420 3.140 ;
        RECT -152.700 2.660 -151.500 3.140 ;
        RECT -142.780 2.660 -141.580 3.140 ;
        RECT -132.860 2.660 -131.660 3.140 ;
        RECT -122.940 2.660 -121.740 3.140 ;
        RECT -113.020 2.660 -111.820 3.140 ;
        RECT -103.100 2.660 -101.900 3.140 ;
        RECT -93.180 2.660 -91.980 3.140 ;
        RECT -83.260 2.660 -82.060 3.140 ;
        RECT -73.340 2.660 -72.140 3.140 ;
        RECT -63.420 2.660 -62.220 3.140 ;
        RECT -53.500 2.660 -52.300 3.140 ;
        RECT -43.580 2.660 -42.380 3.140 ;
        RECT -33.660 2.660 -32.460 3.140 ;
        RECT -23.740 2.660 -22.540 3.140 ;
        RECT -13.820 2.660 -12.620 3.140 ;
        RECT -3.900 2.660 -2.700 3.140 ;
        RECT 6.020 2.660 7.220 3.140 ;
        RECT 15.940 2.660 17.140 3.140 ;
        RECT 25.860 2.660 26.690 3.140 ;
        RECT -286.730 1.090 -285.310 1.500 ;
        RECT -276.810 1.090 -275.390 1.500 ;
        RECT -266.890 1.090 -265.470 1.500 ;
        RECT -256.970 1.090 -255.550 1.500 ;
        RECT -247.050 1.090 -245.630 1.500 ;
        RECT -237.130 1.090 -235.710 1.500 ;
        RECT -227.210 1.090 -225.790 1.500 ;
        RECT -217.290 1.090 -215.870 1.500 ;
        RECT -207.370 1.090 -205.950 1.500 ;
        RECT -197.450 1.090 -196.030 1.500 ;
        RECT -187.530 1.090 -186.110 1.500 ;
        RECT -177.610 1.090 -176.190 1.500 ;
        RECT -167.690 1.090 -166.270 1.500 ;
        RECT -157.770 1.090 -156.350 1.500 ;
        RECT -147.850 1.090 -146.430 1.500 ;
        RECT -137.930 1.090 -136.510 1.500 ;
        RECT -128.010 1.090 -126.590 1.500 ;
        RECT -118.090 1.090 -116.670 1.500 ;
        RECT -108.170 1.090 -106.750 1.500 ;
        RECT -98.250 1.090 -96.830 1.500 ;
        RECT -88.330 1.090 -86.910 1.500 ;
        RECT -78.410 1.090 -76.990 1.500 ;
        RECT -68.490 1.090 -67.070 1.500 ;
        RECT -58.570 1.090 -57.150 1.500 ;
        RECT -48.650 1.090 -47.230 1.500 ;
        RECT -38.730 1.090 -37.310 1.500 ;
        RECT -28.810 1.090 -27.390 1.500 ;
        RECT -18.890 1.090 -17.470 1.500 ;
        RECT -8.970 1.090 -7.550 1.500 ;
        RECT 0.950 1.090 2.370 1.500 ;
        RECT 10.870 1.090 12.290 1.500 ;
        RECT 20.790 1.090 22.210 1.500 ;
        RECT -280.010 -86.330 -278.590 -85.920 ;
        RECT -270.090 -86.330 -268.670 -85.920 ;
        RECT -260.170 -86.330 -258.750 -85.920 ;
        RECT -250.250 -86.330 -248.830 -85.920 ;
        RECT -240.330 -86.330 -238.910 -85.920 ;
        RECT -230.410 -86.330 -228.990 -85.920 ;
        RECT -220.490 -86.330 -219.070 -85.920 ;
        RECT -210.570 -86.330 -209.150 -85.920 ;
        RECT -200.650 -86.330 -199.230 -85.920 ;
        RECT -190.730 -86.330 -189.310 -85.920 ;
        RECT -180.810 -86.330 -179.390 -85.920 ;
        RECT -170.890 -86.330 -169.470 -85.920 ;
        RECT -160.970 -86.330 -159.550 -85.920 ;
        RECT -151.050 -86.330 -149.630 -85.920 ;
        RECT -141.130 -86.330 -139.710 -85.920 ;
        RECT -131.210 -86.330 -129.790 -85.920 ;
        RECT -121.290 -86.330 -119.870 -85.920 ;
        RECT -111.370 -86.330 -109.950 -85.920 ;
        RECT -101.450 -86.330 -100.030 -85.920 ;
        RECT -91.530 -86.330 -90.110 -85.920 ;
        RECT -81.610 -86.330 -80.190 -85.920 ;
        RECT -71.690 -86.330 -70.270 -85.920 ;
        RECT -61.770 -86.330 -60.350 -85.920 ;
        RECT -51.850 -86.330 -50.430 -85.920 ;
        RECT -41.930 -86.330 -40.510 -85.920 ;
        RECT -32.010 -86.330 -30.590 -85.920 ;
        RECT -22.090 -86.330 -20.670 -85.920 ;
        RECT -12.170 -86.330 -10.750 -85.920 ;
        RECT -2.250 -86.330 -0.830 -85.920 ;
        RECT 7.670 -86.330 9.090 -85.920 ;
        RECT 17.590 -86.330 19.010 -85.920 ;
        RECT 27.510 -86.330 28.450 -85.920 ;
        RECT -270.090 -86.700 -268.680 -86.330 ;
        RECT -284.860 -87.970 -283.660 -87.490 ;
        RECT -274.940 -87.970 -273.740 -87.490 ;
        RECT -265.020 -87.970 -263.820 -87.490 ;
        RECT -255.100 -87.970 -253.900 -87.490 ;
        RECT -245.180 -87.970 -243.980 -87.490 ;
        RECT -235.260 -87.970 -234.060 -87.490 ;
        RECT -225.340 -87.970 -224.140 -87.490 ;
        RECT -215.420 -87.970 -214.220 -87.490 ;
        RECT -205.500 -87.970 -204.300 -87.490 ;
        RECT -195.580 -87.970 -194.380 -87.490 ;
        RECT -185.660 -87.970 -184.460 -87.490 ;
        RECT -175.740 -87.970 -174.540 -87.490 ;
        RECT -165.820 -87.970 -164.620 -87.490 ;
        RECT -155.900 -87.970 -154.700 -87.490 ;
        RECT -145.980 -87.970 -144.780 -87.490 ;
        RECT -136.060 -87.970 -134.860 -87.490 ;
        RECT -126.140 -87.970 -124.940 -87.490 ;
        RECT -116.220 -87.970 -115.020 -87.490 ;
        RECT -106.300 -87.970 -105.100 -87.490 ;
        RECT -96.380 -87.970 -95.180 -87.490 ;
        RECT -86.460 -87.970 -85.260 -87.490 ;
        RECT -76.540 -87.970 -75.340 -87.490 ;
        RECT -66.620 -87.970 -65.420 -87.490 ;
        RECT -56.700 -87.970 -55.500 -87.490 ;
        RECT -46.780 -87.970 -45.580 -87.490 ;
        RECT -36.860 -87.970 -35.660 -87.490 ;
        RECT -26.940 -87.970 -25.740 -87.490 ;
        RECT -17.020 -87.970 -15.820 -87.490 ;
        RECT -7.100 -87.970 -5.900 -87.490 ;
        RECT 2.820 -87.970 4.020 -87.490 ;
        RECT 12.740 -87.970 13.940 -87.490 ;
        RECT 22.660 -87.970 23.860 -87.490 ;
        RECT -279.900 -90.690 -278.700 -90.210 ;
        RECT -269.980 -90.690 -268.780 -90.210 ;
        RECT -260.060 -90.690 -258.860 -90.210 ;
        RECT -250.140 -90.690 -248.940 -90.210 ;
        RECT -240.220 -90.690 -239.020 -90.210 ;
        RECT -230.300 -90.690 -229.100 -90.210 ;
        RECT -220.380 -90.690 -219.180 -90.210 ;
        RECT -210.460 -90.690 -209.260 -90.210 ;
        RECT -200.540 -90.690 -199.340 -90.210 ;
        RECT -190.620 -90.690 -189.420 -90.210 ;
        RECT -180.700 -90.690 -179.500 -90.210 ;
        RECT -170.780 -90.690 -169.580 -90.210 ;
        RECT -160.860 -90.690 -159.660 -90.210 ;
        RECT -150.940 -90.690 -149.740 -90.210 ;
        RECT -141.020 -90.690 -139.820 -90.210 ;
        RECT -131.100 -90.690 -129.900 -90.210 ;
        RECT -121.180 -90.690 -119.980 -90.210 ;
        RECT -111.260 -90.690 -110.060 -90.210 ;
        RECT -101.340 -90.690 -100.140 -90.210 ;
        RECT -91.420 -90.690 -90.220 -90.210 ;
        RECT -81.500 -90.690 -80.300 -90.210 ;
        RECT -71.580 -90.690 -70.380 -90.210 ;
        RECT -61.660 -90.690 -60.460 -90.210 ;
        RECT -51.740 -90.690 -50.540 -90.210 ;
        RECT -41.820 -90.690 -40.620 -90.210 ;
        RECT -31.900 -90.690 -30.700 -90.210 ;
        RECT -21.980 -90.690 -20.780 -90.210 ;
        RECT -12.060 -90.690 -10.860 -90.210 ;
        RECT -2.140 -90.690 -0.940 -90.210 ;
        RECT 7.780 -90.690 8.980 -90.210 ;
        RECT 17.700 -90.690 18.900 -90.210 ;
        RECT 27.620 -90.690 28.450 -90.210 ;
        RECT -284.970 -92.260 -283.550 -91.850 ;
        RECT -275.050 -92.260 -273.630 -91.850 ;
        RECT -265.130 -92.260 -263.710 -91.850 ;
        RECT -255.210 -92.260 -253.790 -91.850 ;
        RECT -245.290 -92.260 -243.870 -91.850 ;
        RECT -235.370 -92.260 -233.950 -91.850 ;
        RECT -225.450 -92.260 -224.030 -91.850 ;
        RECT -215.530 -92.260 -214.110 -91.850 ;
        RECT -205.610 -92.260 -204.190 -91.850 ;
        RECT -195.690 -92.260 -194.270 -91.850 ;
        RECT -185.770 -92.260 -184.350 -91.850 ;
        RECT -175.850 -92.260 -174.430 -91.850 ;
        RECT -165.930 -92.260 -164.510 -91.850 ;
        RECT -156.010 -92.260 -154.590 -91.850 ;
        RECT -146.090 -92.260 -144.670 -91.850 ;
        RECT -136.170 -92.260 -134.750 -91.850 ;
        RECT -126.250 -92.260 -124.830 -91.850 ;
        RECT -116.330 -92.260 -114.910 -91.850 ;
        RECT -106.410 -92.260 -104.990 -91.850 ;
        RECT -96.490 -92.260 -95.070 -91.850 ;
        RECT -86.570 -92.260 -85.150 -91.850 ;
        RECT -76.650 -92.260 -75.230 -91.850 ;
        RECT -66.730 -92.260 -65.310 -91.850 ;
        RECT -56.810 -92.260 -55.390 -91.850 ;
        RECT -46.890 -92.260 -45.470 -91.850 ;
        RECT -36.970 -92.260 -35.550 -91.850 ;
        RECT -27.050 -92.260 -25.630 -91.850 ;
        RECT -17.130 -92.260 -15.710 -91.850 ;
        RECT -7.210 -92.260 -5.790 -91.850 ;
        RECT 2.710 -92.260 4.130 -91.850 ;
        RECT 12.630 -92.260 14.050 -91.850 ;
        RECT 22.550 -92.260 23.970 -91.850 ;
        RECT -279.760 -174.040 -278.340 -173.630 ;
        RECT -269.840 -174.040 -268.420 -173.630 ;
        RECT -259.920 -174.040 -258.500 -173.630 ;
        RECT -250.000 -174.040 -248.580 -173.630 ;
        RECT -240.080 -174.040 -238.660 -173.630 ;
        RECT -230.160 -174.040 -228.740 -173.630 ;
        RECT -220.240 -174.040 -218.820 -173.630 ;
        RECT -210.320 -174.040 -208.900 -173.630 ;
        RECT -200.400 -174.040 -198.980 -173.630 ;
        RECT -190.480 -174.040 -189.060 -173.630 ;
        RECT -180.560 -174.040 -179.140 -173.630 ;
        RECT -170.640 -174.040 -169.220 -173.630 ;
        RECT -160.720 -174.040 -159.300 -173.630 ;
        RECT -150.800 -174.040 -149.380 -173.630 ;
        RECT -140.880 -174.040 -139.460 -173.630 ;
        RECT -130.960 -174.040 -129.540 -173.630 ;
        RECT -121.040 -174.040 -119.620 -173.630 ;
        RECT -111.120 -174.040 -109.700 -173.630 ;
        RECT -101.200 -174.040 -99.780 -173.630 ;
        RECT -91.280 -174.040 -89.860 -173.630 ;
        RECT -81.360 -174.040 -79.940 -173.630 ;
        RECT -71.440 -174.040 -70.020 -173.630 ;
        RECT -61.520 -174.040 -60.100 -173.630 ;
        RECT -51.600 -174.040 -50.180 -173.630 ;
        RECT -41.680 -174.040 -40.260 -173.630 ;
        RECT -31.760 -174.040 -30.340 -173.630 ;
        RECT -21.840 -174.040 -20.420 -173.630 ;
        RECT -11.920 -174.040 -10.500 -173.630 ;
        RECT -2.000 -174.040 -0.580 -173.630 ;
        RECT 7.920 -174.040 9.340 -173.630 ;
        RECT 17.840 -174.040 19.260 -173.630 ;
        RECT 27.760 -174.040 28.700 -173.630 ;
        RECT -269.840 -174.410 -268.430 -174.040 ;
        RECT -284.610 -175.680 -283.410 -175.200 ;
        RECT -274.690 -175.680 -273.490 -175.200 ;
        RECT -264.770 -175.680 -263.570 -175.200 ;
        RECT -254.850 -175.680 -253.650 -175.200 ;
        RECT -244.930 -175.680 -243.730 -175.200 ;
        RECT -235.010 -175.680 -233.810 -175.200 ;
        RECT -225.090 -175.680 -223.890 -175.200 ;
        RECT -215.170 -175.680 -213.970 -175.200 ;
        RECT -205.250 -175.680 -204.050 -175.200 ;
        RECT -195.330 -175.680 -194.130 -175.200 ;
        RECT -185.410 -175.680 -184.210 -175.200 ;
        RECT -175.490 -175.680 -174.290 -175.200 ;
        RECT -165.570 -175.680 -164.370 -175.200 ;
        RECT -155.650 -175.680 -154.450 -175.200 ;
        RECT -145.730 -175.680 -144.530 -175.200 ;
        RECT -135.810 -175.680 -134.610 -175.200 ;
        RECT -125.890 -175.680 -124.690 -175.200 ;
        RECT -115.970 -175.680 -114.770 -175.200 ;
        RECT -106.050 -175.680 -104.850 -175.200 ;
        RECT -96.130 -175.680 -94.930 -175.200 ;
        RECT -86.210 -175.680 -85.010 -175.200 ;
        RECT -76.290 -175.680 -75.090 -175.200 ;
        RECT -66.370 -175.680 -65.170 -175.200 ;
        RECT -56.450 -175.680 -55.250 -175.200 ;
        RECT -46.530 -175.680 -45.330 -175.200 ;
        RECT -36.610 -175.680 -35.410 -175.200 ;
        RECT -26.690 -175.680 -25.490 -175.200 ;
        RECT -16.770 -175.680 -15.570 -175.200 ;
        RECT -6.850 -175.680 -5.650 -175.200 ;
        RECT 3.070 -175.680 4.270 -175.200 ;
        RECT 12.990 -175.680 14.190 -175.200 ;
        RECT 22.910 -175.680 24.110 -175.200 ;
        RECT -279.650 -178.400 -278.450 -177.920 ;
        RECT -269.730 -178.400 -268.530 -177.920 ;
        RECT -259.810 -178.400 -258.610 -177.920 ;
        RECT -249.890 -178.400 -248.690 -177.920 ;
        RECT -239.970 -178.400 -238.770 -177.920 ;
        RECT -230.050 -178.400 -228.850 -177.920 ;
        RECT -220.130 -178.400 -218.930 -177.920 ;
        RECT -210.210 -178.400 -209.010 -177.920 ;
        RECT -200.290 -178.400 -199.090 -177.920 ;
        RECT -190.370 -178.400 -189.170 -177.920 ;
        RECT -180.450 -178.400 -179.250 -177.920 ;
        RECT -170.530 -178.400 -169.330 -177.920 ;
        RECT -160.610 -178.400 -159.410 -177.920 ;
        RECT -150.690 -178.400 -149.490 -177.920 ;
        RECT -140.770 -178.400 -139.570 -177.920 ;
        RECT -130.850 -178.400 -129.650 -177.920 ;
        RECT -120.930 -178.400 -119.730 -177.920 ;
        RECT -111.010 -178.400 -109.810 -177.920 ;
        RECT -101.090 -178.400 -99.890 -177.920 ;
        RECT -91.170 -178.400 -89.970 -177.920 ;
        RECT -81.250 -178.400 -80.050 -177.920 ;
        RECT -71.330 -178.400 -70.130 -177.920 ;
        RECT -61.410 -178.400 -60.210 -177.920 ;
        RECT -51.490 -178.400 -50.290 -177.920 ;
        RECT -41.570 -178.400 -40.370 -177.920 ;
        RECT -31.650 -178.400 -30.450 -177.920 ;
        RECT -21.730 -178.400 -20.530 -177.920 ;
        RECT -11.810 -178.400 -10.610 -177.920 ;
        RECT -1.890 -178.400 -0.690 -177.920 ;
        RECT 8.030 -178.400 9.230 -177.920 ;
        RECT 17.950 -178.400 19.150 -177.920 ;
        RECT 27.870 -178.400 28.700 -177.920 ;
        RECT -284.720 -179.970 -283.300 -179.560 ;
        RECT -274.800 -179.970 -273.380 -179.560 ;
        RECT -264.880 -179.970 -263.460 -179.560 ;
        RECT -254.960 -179.970 -253.540 -179.560 ;
        RECT -245.040 -179.970 -243.620 -179.560 ;
        RECT -235.120 -179.970 -233.700 -179.560 ;
        RECT -225.200 -179.970 -223.780 -179.560 ;
        RECT -215.280 -179.970 -213.860 -179.560 ;
        RECT -205.360 -179.970 -203.940 -179.560 ;
        RECT -195.440 -179.970 -194.020 -179.560 ;
        RECT -185.520 -179.970 -184.100 -179.560 ;
        RECT -175.600 -179.970 -174.180 -179.560 ;
        RECT -165.680 -179.970 -164.260 -179.560 ;
        RECT -155.760 -179.970 -154.340 -179.560 ;
        RECT -145.840 -179.970 -144.420 -179.560 ;
        RECT -135.920 -179.970 -134.500 -179.560 ;
        RECT -126.000 -179.970 -124.580 -179.560 ;
        RECT -116.080 -179.970 -114.660 -179.560 ;
        RECT -106.160 -179.970 -104.740 -179.560 ;
        RECT -96.240 -179.970 -94.820 -179.560 ;
        RECT -86.320 -179.970 -84.900 -179.560 ;
        RECT -76.400 -179.970 -74.980 -179.560 ;
        RECT -66.480 -179.970 -65.060 -179.560 ;
        RECT -56.560 -179.970 -55.140 -179.560 ;
        RECT -46.640 -179.970 -45.220 -179.560 ;
        RECT -36.720 -179.970 -35.300 -179.560 ;
        RECT -26.800 -179.970 -25.380 -179.560 ;
        RECT -16.880 -179.970 -15.460 -179.560 ;
        RECT -6.960 -179.970 -5.540 -179.560 ;
        RECT 2.960 -179.970 4.380 -179.560 ;
        RECT 12.880 -179.970 14.300 -179.560 ;
        RECT 22.800 -179.970 24.220 -179.560 ;
      LAYER via2 ;
        RECT -281.915 94.770 -281.635 95.050 ;
        RECT -280.985 94.760 -280.705 95.040 ;
        RECT -271.995 94.770 -271.715 95.050 ;
        RECT -271.065 94.760 -270.785 95.040 ;
        RECT -262.075 94.770 -261.795 95.050 ;
        RECT -261.145 94.760 -260.865 95.040 ;
        RECT -252.155 94.770 -251.875 95.050 ;
        RECT -251.225 94.760 -250.945 95.040 ;
        RECT -242.235 94.770 -241.955 95.050 ;
        RECT -241.305 94.760 -241.025 95.040 ;
        RECT -232.315 94.770 -232.035 95.050 ;
        RECT -231.385 94.760 -231.105 95.040 ;
        RECT -222.395 94.770 -222.115 95.050 ;
        RECT -221.465 94.760 -221.185 95.040 ;
        RECT -212.475 94.770 -212.195 95.050 ;
        RECT -211.545 94.760 -211.265 95.040 ;
        RECT -202.555 94.770 -202.275 95.050 ;
        RECT -201.625 94.760 -201.345 95.040 ;
        RECT -192.635 94.770 -192.355 95.050 ;
        RECT -191.705 94.760 -191.425 95.040 ;
        RECT -182.715 94.770 -182.435 95.050 ;
        RECT -181.785 94.760 -181.505 95.040 ;
        RECT -172.795 94.770 -172.515 95.050 ;
        RECT -171.865 94.760 -171.585 95.040 ;
        RECT -162.875 94.770 -162.595 95.050 ;
        RECT -161.945 94.760 -161.665 95.040 ;
        RECT -152.955 94.770 -152.675 95.050 ;
        RECT -152.025 94.760 -151.745 95.040 ;
        RECT -143.035 94.770 -142.755 95.050 ;
        RECT -142.105 94.760 -141.825 95.040 ;
        RECT -133.115 94.770 -132.835 95.050 ;
        RECT -132.185 94.760 -131.905 95.040 ;
        RECT -123.195 94.770 -122.915 95.050 ;
        RECT -122.265 94.760 -121.985 95.040 ;
        RECT -113.275 94.770 -112.995 95.050 ;
        RECT -112.345 94.760 -112.065 95.040 ;
        RECT -103.355 94.770 -103.075 95.050 ;
        RECT -102.425 94.760 -102.145 95.040 ;
        RECT -93.435 94.770 -93.155 95.050 ;
        RECT -92.505 94.760 -92.225 95.040 ;
        RECT -83.515 94.770 -83.235 95.050 ;
        RECT -82.585 94.760 -82.305 95.040 ;
        RECT -73.595 94.770 -73.315 95.050 ;
        RECT -72.665 94.760 -72.385 95.040 ;
        RECT -63.675 94.770 -63.395 95.050 ;
        RECT -62.745 94.760 -62.465 95.040 ;
        RECT -53.755 94.770 -53.475 95.050 ;
        RECT -52.825 94.760 -52.545 95.040 ;
        RECT -43.835 94.770 -43.555 95.050 ;
        RECT -42.905 94.760 -42.625 95.040 ;
        RECT -33.915 94.770 -33.635 95.050 ;
        RECT -32.985 94.760 -32.705 95.040 ;
        RECT -23.995 94.770 -23.715 95.050 ;
        RECT -23.065 94.760 -22.785 95.040 ;
        RECT -14.075 94.770 -13.795 95.050 ;
        RECT -13.145 94.760 -12.865 95.040 ;
        RECT -4.155 94.770 -3.875 95.050 ;
        RECT -3.225 94.760 -2.945 95.040 ;
        RECT 5.765 94.770 6.045 95.050 ;
        RECT 6.695 94.760 6.975 95.040 ;
        RECT 15.685 94.770 15.965 95.050 ;
        RECT 16.615 94.760 16.895 95.040 ;
        RECT 25.605 94.770 25.885 95.050 ;
        RECT -286.575 93.280 -286.295 93.560 ;
        RECT -276.655 93.280 -276.375 93.560 ;
        RECT -266.735 93.280 -266.455 93.560 ;
        RECT -256.815 93.280 -256.535 93.560 ;
        RECT -246.895 93.280 -246.615 93.560 ;
        RECT -236.975 93.280 -236.695 93.560 ;
        RECT -227.055 93.280 -226.775 93.560 ;
        RECT -217.135 93.280 -216.855 93.560 ;
        RECT -207.215 93.280 -206.935 93.560 ;
        RECT -197.295 93.280 -197.015 93.560 ;
        RECT -187.375 93.280 -187.095 93.560 ;
        RECT -177.455 93.280 -177.175 93.560 ;
        RECT -167.535 93.280 -167.255 93.560 ;
        RECT -157.615 93.280 -157.335 93.560 ;
        RECT -147.695 93.280 -147.415 93.560 ;
        RECT -137.775 93.280 -137.495 93.560 ;
        RECT -127.855 93.280 -127.575 93.560 ;
        RECT -117.935 93.280 -117.655 93.560 ;
        RECT -108.015 93.280 -107.735 93.560 ;
        RECT -98.095 93.280 -97.815 93.560 ;
        RECT -88.175 93.280 -87.895 93.560 ;
        RECT -78.255 93.280 -77.975 93.560 ;
        RECT -68.335 93.280 -68.055 93.560 ;
        RECT -58.415 93.280 -58.135 93.560 ;
        RECT -48.495 93.280 -48.215 93.560 ;
        RECT -38.575 93.280 -38.295 93.560 ;
        RECT -28.655 93.280 -28.375 93.560 ;
        RECT -18.735 93.280 -18.455 93.560 ;
        RECT -8.815 93.280 -8.535 93.560 ;
        RECT 1.105 93.280 1.385 93.560 ;
        RECT 11.025 93.280 11.305 93.560 ;
        RECT 20.945 93.280 21.225 93.560 ;
        RECT -281.535 90.420 -281.255 90.700 ;
        RECT -271.615 90.420 -271.335 90.700 ;
        RECT -261.695 90.420 -261.415 90.700 ;
        RECT -251.775 90.420 -251.495 90.700 ;
        RECT -241.855 90.420 -241.575 90.700 ;
        RECT -231.935 90.420 -231.655 90.700 ;
        RECT -222.015 90.420 -221.735 90.700 ;
        RECT -212.095 90.420 -211.815 90.700 ;
        RECT -202.175 90.420 -201.895 90.700 ;
        RECT -192.255 90.420 -191.975 90.700 ;
        RECT -182.335 90.420 -182.055 90.700 ;
        RECT -172.415 90.420 -172.135 90.700 ;
        RECT -162.495 90.420 -162.215 90.700 ;
        RECT -152.575 90.420 -152.295 90.700 ;
        RECT -142.655 90.420 -142.375 90.700 ;
        RECT -132.735 90.420 -132.455 90.700 ;
        RECT -122.815 90.420 -122.535 90.700 ;
        RECT -112.895 90.420 -112.615 90.700 ;
        RECT -102.975 90.420 -102.695 90.700 ;
        RECT -93.055 90.420 -92.775 90.700 ;
        RECT -83.135 90.420 -82.855 90.700 ;
        RECT -73.215 90.420 -72.935 90.700 ;
        RECT -63.295 90.420 -63.015 90.700 ;
        RECT -53.375 90.420 -53.095 90.700 ;
        RECT -43.455 90.420 -43.175 90.700 ;
        RECT -33.535 90.420 -33.255 90.700 ;
        RECT -23.615 90.420 -23.335 90.700 ;
        RECT -13.695 90.420 -13.415 90.700 ;
        RECT -3.775 90.420 -3.495 90.700 ;
        RECT 6.145 90.420 6.425 90.700 ;
        RECT 16.065 90.420 16.345 90.700 ;
        RECT 25.985 90.420 26.265 90.700 ;
        RECT -286.875 88.880 -286.595 89.160 ;
        RECT -285.945 88.880 -285.665 89.160 ;
        RECT -276.955 88.880 -276.675 89.160 ;
        RECT -276.025 88.880 -275.745 89.160 ;
        RECT -267.035 88.880 -266.755 89.160 ;
        RECT -266.105 88.880 -265.825 89.160 ;
        RECT -257.115 88.880 -256.835 89.160 ;
        RECT -256.185 88.880 -255.905 89.160 ;
        RECT -247.195 88.880 -246.915 89.160 ;
        RECT -246.265 88.880 -245.985 89.160 ;
        RECT -237.275 88.880 -236.995 89.160 ;
        RECT -236.345 88.880 -236.065 89.160 ;
        RECT -227.355 88.880 -227.075 89.160 ;
        RECT -226.425 88.880 -226.145 89.160 ;
        RECT -217.435 88.880 -217.155 89.160 ;
        RECT -216.505 88.880 -216.225 89.160 ;
        RECT -207.515 88.880 -207.235 89.160 ;
        RECT -206.585 88.880 -206.305 89.160 ;
        RECT -197.595 88.880 -197.315 89.160 ;
        RECT -196.665 88.880 -196.385 89.160 ;
        RECT -187.675 88.880 -187.395 89.160 ;
        RECT -186.745 88.880 -186.465 89.160 ;
        RECT -177.755 88.880 -177.475 89.160 ;
        RECT -176.825 88.880 -176.545 89.160 ;
        RECT -167.835 88.880 -167.555 89.160 ;
        RECT -166.905 88.880 -166.625 89.160 ;
        RECT -157.915 88.880 -157.635 89.160 ;
        RECT -156.985 88.880 -156.705 89.160 ;
        RECT -147.995 88.880 -147.715 89.160 ;
        RECT -147.065 88.880 -146.785 89.160 ;
        RECT -138.075 88.880 -137.795 89.160 ;
        RECT -137.145 88.880 -136.865 89.160 ;
        RECT -128.155 88.880 -127.875 89.160 ;
        RECT -127.225 88.880 -126.945 89.160 ;
        RECT -118.235 88.880 -117.955 89.160 ;
        RECT -117.305 88.880 -117.025 89.160 ;
        RECT -108.315 88.880 -108.035 89.160 ;
        RECT -107.385 88.880 -107.105 89.160 ;
        RECT -98.395 88.880 -98.115 89.160 ;
        RECT -97.465 88.880 -97.185 89.160 ;
        RECT -88.475 88.880 -88.195 89.160 ;
        RECT -87.545 88.880 -87.265 89.160 ;
        RECT -78.555 88.880 -78.275 89.160 ;
        RECT -77.625 88.880 -77.345 89.160 ;
        RECT -68.635 88.880 -68.355 89.160 ;
        RECT -67.705 88.880 -67.425 89.160 ;
        RECT -58.715 88.880 -58.435 89.160 ;
        RECT -57.785 88.880 -57.505 89.160 ;
        RECT -48.795 88.880 -48.515 89.160 ;
        RECT -47.865 88.880 -47.585 89.160 ;
        RECT -38.875 88.880 -38.595 89.160 ;
        RECT -37.945 88.880 -37.665 89.160 ;
        RECT -28.955 88.880 -28.675 89.160 ;
        RECT -28.025 88.880 -27.745 89.160 ;
        RECT -19.035 88.880 -18.755 89.160 ;
        RECT -18.105 88.880 -17.825 89.160 ;
        RECT -9.115 88.880 -8.835 89.160 ;
        RECT -8.185 88.880 -7.905 89.160 ;
        RECT 0.805 88.880 1.085 89.160 ;
        RECT 1.735 88.880 2.015 89.160 ;
        RECT 10.725 88.880 11.005 89.160 ;
        RECT 11.655 88.880 11.935 89.160 ;
        RECT 20.645 88.880 20.925 89.160 ;
        RECT 21.575 88.880 21.855 89.160 ;
        RECT -281.665 7.060 -281.385 7.340 ;
        RECT -280.735 7.050 -280.455 7.330 ;
        RECT -271.745 7.060 -271.465 7.340 ;
        RECT -270.815 7.050 -270.535 7.330 ;
        RECT -261.825 7.060 -261.545 7.340 ;
        RECT -260.895 7.050 -260.615 7.330 ;
        RECT -251.905 7.060 -251.625 7.340 ;
        RECT -250.975 7.050 -250.695 7.330 ;
        RECT -241.985 7.060 -241.705 7.340 ;
        RECT -241.055 7.050 -240.775 7.330 ;
        RECT -232.065 7.060 -231.785 7.340 ;
        RECT -231.135 7.050 -230.855 7.330 ;
        RECT -222.145 7.060 -221.865 7.340 ;
        RECT -221.215 7.050 -220.935 7.330 ;
        RECT -212.225 7.060 -211.945 7.340 ;
        RECT -211.295 7.050 -211.015 7.330 ;
        RECT -202.305 7.060 -202.025 7.340 ;
        RECT -201.375 7.050 -201.095 7.330 ;
        RECT -192.385 7.060 -192.105 7.340 ;
        RECT -191.455 7.050 -191.175 7.330 ;
        RECT -182.465 7.060 -182.185 7.340 ;
        RECT -181.535 7.050 -181.255 7.330 ;
        RECT -172.545 7.060 -172.265 7.340 ;
        RECT -171.615 7.050 -171.335 7.330 ;
        RECT -162.625 7.060 -162.345 7.340 ;
        RECT -161.695 7.050 -161.415 7.330 ;
        RECT -152.705 7.060 -152.425 7.340 ;
        RECT -151.775 7.050 -151.495 7.330 ;
        RECT -142.785 7.060 -142.505 7.340 ;
        RECT -141.855 7.050 -141.575 7.330 ;
        RECT -132.865 7.060 -132.585 7.340 ;
        RECT -131.935 7.050 -131.655 7.330 ;
        RECT -122.945 7.060 -122.665 7.340 ;
        RECT -122.015 7.050 -121.735 7.330 ;
        RECT -113.025 7.060 -112.745 7.340 ;
        RECT -112.095 7.050 -111.815 7.330 ;
        RECT -103.105 7.060 -102.825 7.340 ;
        RECT -102.175 7.050 -101.895 7.330 ;
        RECT -93.185 7.060 -92.905 7.340 ;
        RECT -92.255 7.050 -91.975 7.330 ;
        RECT -83.265 7.060 -82.985 7.340 ;
        RECT -82.335 7.050 -82.055 7.330 ;
        RECT -73.345 7.060 -73.065 7.340 ;
        RECT -72.415 7.050 -72.135 7.330 ;
        RECT -63.425 7.060 -63.145 7.340 ;
        RECT -62.495 7.050 -62.215 7.330 ;
        RECT -53.505 7.060 -53.225 7.340 ;
        RECT -52.575 7.050 -52.295 7.330 ;
        RECT -43.585 7.060 -43.305 7.340 ;
        RECT -42.655 7.050 -42.375 7.330 ;
        RECT -33.665 7.060 -33.385 7.340 ;
        RECT -32.735 7.050 -32.455 7.330 ;
        RECT -23.745 7.060 -23.465 7.340 ;
        RECT -22.815 7.050 -22.535 7.330 ;
        RECT -13.825 7.060 -13.545 7.340 ;
        RECT -12.895 7.050 -12.615 7.330 ;
        RECT -3.905 7.060 -3.625 7.340 ;
        RECT -2.975 7.050 -2.695 7.330 ;
        RECT 6.015 7.060 6.295 7.340 ;
        RECT 6.945 7.050 7.225 7.330 ;
        RECT 15.935 7.060 16.215 7.340 ;
        RECT 16.865 7.050 17.145 7.330 ;
        RECT 25.855 7.060 26.135 7.340 ;
        RECT -286.325 5.570 -286.045 5.850 ;
        RECT -276.405 5.570 -276.125 5.850 ;
        RECT -266.485 5.570 -266.205 5.850 ;
        RECT -256.565 5.570 -256.285 5.850 ;
        RECT -246.645 5.570 -246.365 5.850 ;
        RECT -236.725 5.570 -236.445 5.850 ;
        RECT -226.805 5.570 -226.525 5.850 ;
        RECT -216.885 5.570 -216.605 5.850 ;
        RECT -206.965 5.570 -206.685 5.850 ;
        RECT -197.045 5.570 -196.765 5.850 ;
        RECT -187.125 5.570 -186.845 5.850 ;
        RECT -177.205 5.570 -176.925 5.850 ;
        RECT -167.285 5.570 -167.005 5.850 ;
        RECT -157.365 5.570 -157.085 5.850 ;
        RECT -147.445 5.570 -147.165 5.850 ;
        RECT -137.525 5.570 -137.245 5.850 ;
        RECT -127.605 5.570 -127.325 5.850 ;
        RECT -117.685 5.570 -117.405 5.850 ;
        RECT -107.765 5.570 -107.485 5.850 ;
        RECT -97.845 5.570 -97.565 5.850 ;
        RECT -87.925 5.570 -87.645 5.850 ;
        RECT -78.005 5.570 -77.725 5.850 ;
        RECT -68.085 5.570 -67.805 5.850 ;
        RECT -58.165 5.570 -57.885 5.850 ;
        RECT -48.245 5.570 -47.965 5.850 ;
        RECT -38.325 5.570 -38.045 5.850 ;
        RECT -28.405 5.570 -28.125 5.850 ;
        RECT -18.485 5.570 -18.205 5.850 ;
        RECT -8.565 5.570 -8.285 5.850 ;
        RECT 1.355 5.570 1.635 5.850 ;
        RECT 11.275 5.570 11.555 5.850 ;
        RECT 21.195 5.570 21.475 5.850 ;
        RECT -281.285 2.710 -281.005 2.990 ;
        RECT -271.365 2.710 -271.085 2.990 ;
        RECT -261.445 2.710 -261.165 2.990 ;
        RECT -251.525 2.710 -251.245 2.990 ;
        RECT -241.605 2.710 -241.325 2.990 ;
        RECT -231.685 2.710 -231.405 2.990 ;
        RECT -221.765 2.710 -221.485 2.990 ;
        RECT -211.845 2.710 -211.565 2.990 ;
        RECT -201.925 2.710 -201.645 2.990 ;
        RECT -192.005 2.710 -191.725 2.990 ;
        RECT -182.085 2.710 -181.805 2.990 ;
        RECT -172.165 2.710 -171.885 2.990 ;
        RECT -162.245 2.710 -161.965 2.990 ;
        RECT -152.325 2.710 -152.045 2.990 ;
        RECT -142.405 2.710 -142.125 2.990 ;
        RECT -132.485 2.710 -132.205 2.990 ;
        RECT -122.565 2.710 -122.285 2.990 ;
        RECT -112.645 2.710 -112.365 2.990 ;
        RECT -102.725 2.710 -102.445 2.990 ;
        RECT -92.805 2.710 -92.525 2.990 ;
        RECT -82.885 2.710 -82.605 2.990 ;
        RECT -72.965 2.710 -72.685 2.990 ;
        RECT -63.045 2.710 -62.765 2.990 ;
        RECT -53.125 2.710 -52.845 2.990 ;
        RECT -43.205 2.710 -42.925 2.990 ;
        RECT -33.285 2.710 -33.005 2.990 ;
        RECT -23.365 2.710 -23.085 2.990 ;
        RECT -13.445 2.710 -13.165 2.990 ;
        RECT -3.525 2.710 -3.245 2.990 ;
        RECT 6.395 2.710 6.675 2.990 ;
        RECT 16.315 2.710 16.595 2.990 ;
        RECT 26.235 2.710 26.515 2.990 ;
        RECT -286.625 1.170 -286.345 1.450 ;
        RECT -285.695 1.170 -285.415 1.450 ;
        RECT -276.705 1.170 -276.425 1.450 ;
        RECT -275.775 1.170 -275.495 1.450 ;
        RECT -266.785 1.170 -266.505 1.450 ;
        RECT -265.855 1.170 -265.575 1.450 ;
        RECT -256.865 1.170 -256.585 1.450 ;
        RECT -255.935 1.170 -255.655 1.450 ;
        RECT -246.945 1.170 -246.665 1.450 ;
        RECT -246.015 1.170 -245.735 1.450 ;
        RECT -237.025 1.170 -236.745 1.450 ;
        RECT -236.095 1.170 -235.815 1.450 ;
        RECT -227.105 1.170 -226.825 1.450 ;
        RECT -226.175 1.170 -225.895 1.450 ;
        RECT -217.185 1.170 -216.905 1.450 ;
        RECT -216.255 1.170 -215.975 1.450 ;
        RECT -207.265 1.170 -206.985 1.450 ;
        RECT -206.335 1.170 -206.055 1.450 ;
        RECT -197.345 1.170 -197.065 1.450 ;
        RECT -196.415 1.170 -196.135 1.450 ;
        RECT -187.425 1.170 -187.145 1.450 ;
        RECT -186.495 1.170 -186.215 1.450 ;
        RECT -177.505 1.170 -177.225 1.450 ;
        RECT -176.575 1.170 -176.295 1.450 ;
        RECT -167.585 1.170 -167.305 1.450 ;
        RECT -166.655 1.170 -166.375 1.450 ;
        RECT -157.665 1.170 -157.385 1.450 ;
        RECT -156.735 1.170 -156.455 1.450 ;
        RECT -147.745 1.170 -147.465 1.450 ;
        RECT -146.815 1.170 -146.535 1.450 ;
        RECT -137.825 1.170 -137.545 1.450 ;
        RECT -136.895 1.170 -136.615 1.450 ;
        RECT -127.905 1.170 -127.625 1.450 ;
        RECT -126.975 1.170 -126.695 1.450 ;
        RECT -117.985 1.170 -117.705 1.450 ;
        RECT -117.055 1.170 -116.775 1.450 ;
        RECT -108.065 1.170 -107.785 1.450 ;
        RECT -107.135 1.170 -106.855 1.450 ;
        RECT -98.145 1.170 -97.865 1.450 ;
        RECT -97.215 1.170 -96.935 1.450 ;
        RECT -88.225 1.170 -87.945 1.450 ;
        RECT -87.295 1.170 -87.015 1.450 ;
        RECT -78.305 1.170 -78.025 1.450 ;
        RECT -77.375 1.170 -77.095 1.450 ;
        RECT -68.385 1.170 -68.105 1.450 ;
        RECT -67.455 1.170 -67.175 1.450 ;
        RECT -58.465 1.170 -58.185 1.450 ;
        RECT -57.535 1.170 -57.255 1.450 ;
        RECT -48.545 1.170 -48.265 1.450 ;
        RECT -47.615 1.170 -47.335 1.450 ;
        RECT -38.625 1.170 -38.345 1.450 ;
        RECT -37.695 1.170 -37.415 1.450 ;
        RECT -28.705 1.170 -28.425 1.450 ;
        RECT -27.775 1.170 -27.495 1.450 ;
        RECT -18.785 1.170 -18.505 1.450 ;
        RECT -17.855 1.170 -17.575 1.450 ;
        RECT -8.865 1.170 -8.585 1.450 ;
        RECT -7.935 1.170 -7.655 1.450 ;
        RECT 1.055 1.170 1.335 1.450 ;
        RECT 1.985 1.170 2.265 1.450 ;
        RECT 10.975 1.170 11.255 1.450 ;
        RECT 11.905 1.170 12.185 1.450 ;
        RECT 20.895 1.170 21.175 1.450 ;
        RECT 21.825 1.170 22.105 1.450 ;
        RECT -279.905 -86.290 -279.625 -86.010 ;
        RECT -278.975 -86.300 -278.695 -86.020 ;
        RECT -269.985 -86.290 -269.705 -86.010 ;
        RECT -269.055 -86.300 -268.775 -86.020 ;
        RECT -260.065 -86.290 -259.785 -86.010 ;
        RECT -259.135 -86.300 -258.855 -86.020 ;
        RECT -250.145 -86.290 -249.865 -86.010 ;
        RECT -249.215 -86.300 -248.935 -86.020 ;
        RECT -240.225 -86.290 -239.945 -86.010 ;
        RECT -239.295 -86.300 -239.015 -86.020 ;
        RECT -230.305 -86.290 -230.025 -86.010 ;
        RECT -229.375 -86.300 -229.095 -86.020 ;
        RECT -220.385 -86.290 -220.105 -86.010 ;
        RECT -219.455 -86.300 -219.175 -86.020 ;
        RECT -210.465 -86.290 -210.185 -86.010 ;
        RECT -209.535 -86.300 -209.255 -86.020 ;
        RECT -200.545 -86.290 -200.265 -86.010 ;
        RECT -199.615 -86.300 -199.335 -86.020 ;
        RECT -190.625 -86.290 -190.345 -86.010 ;
        RECT -189.695 -86.300 -189.415 -86.020 ;
        RECT -180.705 -86.290 -180.425 -86.010 ;
        RECT -179.775 -86.300 -179.495 -86.020 ;
        RECT -170.785 -86.290 -170.505 -86.010 ;
        RECT -169.855 -86.300 -169.575 -86.020 ;
        RECT -160.865 -86.290 -160.585 -86.010 ;
        RECT -159.935 -86.300 -159.655 -86.020 ;
        RECT -150.945 -86.290 -150.665 -86.010 ;
        RECT -150.015 -86.300 -149.735 -86.020 ;
        RECT -141.025 -86.290 -140.745 -86.010 ;
        RECT -140.095 -86.300 -139.815 -86.020 ;
        RECT -131.105 -86.290 -130.825 -86.010 ;
        RECT -130.175 -86.300 -129.895 -86.020 ;
        RECT -121.185 -86.290 -120.905 -86.010 ;
        RECT -120.255 -86.300 -119.975 -86.020 ;
        RECT -111.265 -86.290 -110.985 -86.010 ;
        RECT -110.335 -86.300 -110.055 -86.020 ;
        RECT -101.345 -86.290 -101.065 -86.010 ;
        RECT -100.415 -86.300 -100.135 -86.020 ;
        RECT -91.425 -86.290 -91.145 -86.010 ;
        RECT -90.495 -86.300 -90.215 -86.020 ;
        RECT -81.505 -86.290 -81.225 -86.010 ;
        RECT -80.575 -86.300 -80.295 -86.020 ;
        RECT -71.585 -86.290 -71.305 -86.010 ;
        RECT -70.655 -86.300 -70.375 -86.020 ;
        RECT -61.665 -86.290 -61.385 -86.010 ;
        RECT -60.735 -86.300 -60.455 -86.020 ;
        RECT -51.745 -86.290 -51.465 -86.010 ;
        RECT -50.815 -86.300 -50.535 -86.020 ;
        RECT -41.825 -86.290 -41.545 -86.010 ;
        RECT -40.895 -86.300 -40.615 -86.020 ;
        RECT -31.905 -86.290 -31.625 -86.010 ;
        RECT -30.975 -86.300 -30.695 -86.020 ;
        RECT -21.985 -86.290 -21.705 -86.010 ;
        RECT -21.055 -86.300 -20.775 -86.020 ;
        RECT -12.065 -86.290 -11.785 -86.010 ;
        RECT -11.135 -86.300 -10.855 -86.020 ;
        RECT -2.145 -86.290 -1.865 -86.010 ;
        RECT -1.215 -86.300 -0.935 -86.020 ;
        RECT 7.775 -86.290 8.055 -86.010 ;
        RECT 8.705 -86.300 8.985 -86.020 ;
        RECT 17.695 -86.290 17.975 -86.010 ;
        RECT 18.625 -86.300 18.905 -86.020 ;
        RECT 27.615 -86.290 27.895 -86.010 ;
        RECT -284.565 -87.780 -284.285 -87.500 ;
        RECT -274.645 -87.780 -274.365 -87.500 ;
        RECT -264.725 -87.780 -264.445 -87.500 ;
        RECT -254.805 -87.780 -254.525 -87.500 ;
        RECT -244.885 -87.780 -244.605 -87.500 ;
        RECT -234.965 -87.780 -234.685 -87.500 ;
        RECT -225.045 -87.780 -224.765 -87.500 ;
        RECT -215.125 -87.780 -214.845 -87.500 ;
        RECT -205.205 -87.780 -204.925 -87.500 ;
        RECT -195.285 -87.780 -195.005 -87.500 ;
        RECT -185.365 -87.780 -185.085 -87.500 ;
        RECT -175.445 -87.780 -175.165 -87.500 ;
        RECT -165.525 -87.780 -165.245 -87.500 ;
        RECT -155.605 -87.780 -155.325 -87.500 ;
        RECT -145.685 -87.780 -145.405 -87.500 ;
        RECT -135.765 -87.780 -135.485 -87.500 ;
        RECT -125.845 -87.780 -125.565 -87.500 ;
        RECT -115.925 -87.780 -115.645 -87.500 ;
        RECT -106.005 -87.780 -105.725 -87.500 ;
        RECT -96.085 -87.780 -95.805 -87.500 ;
        RECT -86.165 -87.780 -85.885 -87.500 ;
        RECT -76.245 -87.780 -75.965 -87.500 ;
        RECT -66.325 -87.780 -66.045 -87.500 ;
        RECT -56.405 -87.780 -56.125 -87.500 ;
        RECT -46.485 -87.780 -46.205 -87.500 ;
        RECT -36.565 -87.780 -36.285 -87.500 ;
        RECT -26.645 -87.780 -26.365 -87.500 ;
        RECT -16.725 -87.780 -16.445 -87.500 ;
        RECT -6.805 -87.780 -6.525 -87.500 ;
        RECT 3.115 -87.780 3.395 -87.500 ;
        RECT 13.035 -87.780 13.315 -87.500 ;
        RECT 22.955 -87.780 23.235 -87.500 ;
        RECT -279.525 -90.640 -279.245 -90.360 ;
        RECT -269.605 -90.640 -269.325 -90.360 ;
        RECT -259.685 -90.640 -259.405 -90.360 ;
        RECT -249.765 -90.640 -249.485 -90.360 ;
        RECT -239.845 -90.640 -239.565 -90.360 ;
        RECT -229.925 -90.640 -229.645 -90.360 ;
        RECT -220.005 -90.640 -219.725 -90.360 ;
        RECT -210.085 -90.640 -209.805 -90.360 ;
        RECT -200.165 -90.640 -199.885 -90.360 ;
        RECT -190.245 -90.640 -189.965 -90.360 ;
        RECT -180.325 -90.640 -180.045 -90.360 ;
        RECT -170.405 -90.640 -170.125 -90.360 ;
        RECT -160.485 -90.640 -160.205 -90.360 ;
        RECT -150.565 -90.640 -150.285 -90.360 ;
        RECT -140.645 -90.640 -140.365 -90.360 ;
        RECT -130.725 -90.640 -130.445 -90.360 ;
        RECT -120.805 -90.640 -120.525 -90.360 ;
        RECT -110.885 -90.640 -110.605 -90.360 ;
        RECT -100.965 -90.640 -100.685 -90.360 ;
        RECT -91.045 -90.640 -90.765 -90.360 ;
        RECT -81.125 -90.640 -80.845 -90.360 ;
        RECT -71.205 -90.640 -70.925 -90.360 ;
        RECT -61.285 -90.640 -61.005 -90.360 ;
        RECT -51.365 -90.640 -51.085 -90.360 ;
        RECT -41.445 -90.640 -41.165 -90.360 ;
        RECT -31.525 -90.640 -31.245 -90.360 ;
        RECT -21.605 -90.640 -21.325 -90.360 ;
        RECT -11.685 -90.640 -11.405 -90.360 ;
        RECT -1.765 -90.640 -1.485 -90.360 ;
        RECT 8.155 -90.640 8.435 -90.360 ;
        RECT 18.075 -90.640 18.355 -90.360 ;
        RECT 27.995 -90.640 28.275 -90.360 ;
        RECT -284.865 -92.180 -284.585 -91.900 ;
        RECT -283.935 -92.180 -283.655 -91.900 ;
        RECT -274.945 -92.180 -274.665 -91.900 ;
        RECT -274.015 -92.180 -273.735 -91.900 ;
        RECT -265.025 -92.180 -264.745 -91.900 ;
        RECT -264.095 -92.180 -263.815 -91.900 ;
        RECT -255.105 -92.180 -254.825 -91.900 ;
        RECT -254.175 -92.180 -253.895 -91.900 ;
        RECT -245.185 -92.180 -244.905 -91.900 ;
        RECT -244.255 -92.180 -243.975 -91.900 ;
        RECT -235.265 -92.180 -234.985 -91.900 ;
        RECT -234.335 -92.180 -234.055 -91.900 ;
        RECT -225.345 -92.180 -225.065 -91.900 ;
        RECT -224.415 -92.180 -224.135 -91.900 ;
        RECT -215.425 -92.180 -215.145 -91.900 ;
        RECT -214.495 -92.180 -214.215 -91.900 ;
        RECT -205.505 -92.180 -205.225 -91.900 ;
        RECT -204.575 -92.180 -204.295 -91.900 ;
        RECT -195.585 -92.180 -195.305 -91.900 ;
        RECT -194.655 -92.180 -194.375 -91.900 ;
        RECT -185.665 -92.180 -185.385 -91.900 ;
        RECT -184.735 -92.180 -184.455 -91.900 ;
        RECT -175.745 -92.180 -175.465 -91.900 ;
        RECT -174.815 -92.180 -174.535 -91.900 ;
        RECT -165.825 -92.180 -165.545 -91.900 ;
        RECT -164.895 -92.180 -164.615 -91.900 ;
        RECT -155.905 -92.180 -155.625 -91.900 ;
        RECT -154.975 -92.180 -154.695 -91.900 ;
        RECT -145.985 -92.180 -145.705 -91.900 ;
        RECT -145.055 -92.180 -144.775 -91.900 ;
        RECT -136.065 -92.180 -135.785 -91.900 ;
        RECT -135.135 -92.180 -134.855 -91.900 ;
        RECT -126.145 -92.180 -125.865 -91.900 ;
        RECT -125.215 -92.180 -124.935 -91.900 ;
        RECT -116.225 -92.180 -115.945 -91.900 ;
        RECT -115.295 -92.180 -115.015 -91.900 ;
        RECT -106.305 -92.180 -106.025 -91.900 ;
        RECT -105.375 -92.180 -105.095 -91.900 ;
        RECT -96.385 -92.180 -96.105 -91.900 ;
        RECT -95.455 -92.180 -95.175 -91.900 ;
        RECT -86.465 -92.180 -86.185 -91.900 ;
        RECT -85.535 -92.180 -85.255 -91.900 ;
        RECT -76.545 -92.180 -76.265 -91.900 ;
        RECT -75.615 -92.180 -75.335 -91.900 ;
        RECT -66.625 -92.180 -66.345 -91.900 ;
        RECT -65.695 -92.180 -65.415 -91.900 ;
        RECT -56.705 -92.180 -56.425 -91.900 ;
        RECT -55.775 -92.180 -55.495 -91.900 ;
        RECT -46.785 -92.180 -46.505 -91.900 ;
        RECT -45.855 -92.180 -45.575 -91.900 ;
        RECT -36.865 -92.180 -36.585 -91.900 ;
        RECT -35.935 -92.180 -35.655 -91.900 ;
        RECT -26.945 -92.180 -26.665 -91.900 ;
        RECT -26.015 -92.180 -25.735 -91.900 ;
        RECT -17.025 -92.180 -16.745 -91.900 ;
        RECT -16.095 -92.180 -15.815 -91.900 ;
        RECT -7.105 -92.180 -6.825 -91.900 ;
        RECT -6.175 -92.180 -5.895 -91.900 ;
        RECT 2.815 -92.180 3.095 -91.900 ;
        RECT 3.745 -92.180 4.025 -91.900 ;
        RECT 12.735 -92.180 13.015 -91.900 ;
        RECT 13.665 -92.180 13.945 -91.900 ;
        RECT 22.655 -92.180 22.935 -91.900 ;
        RECT 23.585 -92.180 23.865 -91.900 ;
        RECT -279.655 -174.000 -279.375 -173.720 ;
        RECT -278.725 -174.010 -278.445 -173.730 ;
        RECT -269.735 -174.000 -269.455 -173.720 ;
        RECT -268.805 -174.010 -268.525 -173.730 ;
        RECT -259.815 -174.000 -259.535 -173.720 ;
        RECT -258.885 -174.010 -258.605 -173.730 ;
        RECT -249.895 -174.000 -249.615 -173.720 ;
        RECT -248.965 -174.010 -248.685 -173.730 ;
        RECT -239.975 -174.000 -239.695 -173.720 ;
        RECT -239.045 -174.010 -238.765 -173.730 ;
        RECT -230.055 -174.000 -229.775 -173.720 ;
        RECT -229.125 -174.010 -228.845 -173.730 ;
        RECT -220.135 -174.000 -219.855 -173.720 ;
        RECT -219.205 -174.010 -218.925 -173.730 ;
        RECT -210.215 -174.000 -209.935 -173.720 ;
        RECT -209.285 -174.010 -209.005 -173.730 ;
        RECT -200.295 -174.000 -200.015 -173.720 ;
        RECT -199.365 -174.010 -199.085 -173.730 ;
        RECT -190.375 -174.000 -190.095 -173.720 ;
        RECT -189.445 -174.010 -189.165 -173.730 ;
        RECT -180.455 -174.000 -180.175 -173.720 ;
        RECT -179.525 -174.010 -179.245 -173.730 ;
        RECT -170.535 -174.000 -170.255 -173.720 ;
        RECT -169.605 -174.010 -169.325 -173.730 ;
        RECT -160.615 -174.000 -160.335 -173.720 ;
        RECT -159.685 -174.010 -159.405 -173.730 ;
        RECT -150.695 -174.000 -150.415 -173.720 ;
        RECT -149.765 -174.010 -149.485 -173.730 ;
        RECT -140.775 -174.000 -140.495 -173.720 ;
        RECT -139.845 -174.010 -139.565 -173.730 ;
        RECT -130.855 -174.000 -130.575 -173.720 ;
        RECT -129.925 -174.010 -129.645 -173.730 ;
        RECT -120.935 -174.000 -120.655 -173.720 ;
        RECT -120.005 -174.010 -119.725 -173.730 ;
        RECT -111.015 -174.000 -110.735 -173.720 ;
        RECT -110.085 -174.010 -109.805 -173.730 ;
        RECT -101.095 -174.000 -100.815 -173.720 ;
        RECT -100.165 -174.010 -99.885 -173.730 ;
        RECT -91.175 -174.000 -90.895 -173.720 ;
        RECT -90.245 -174.010 -89.965 -173.730 ;
        RECT -81.255 -174.000 -80.975 -173.720 ;
        RECT -80.325 -174.010 -80.045 -173.730 ;
        RECT -71.335 -174.000 -71.055 -173.720 ;
        RECT -70.405 -174.010 -70.125 -173.730 ;
        RECT -61.415 -174.000 -61.135 -173.720 ;
        RECT -60.485 -174.010 -60.205 -173.730 ;
        RECT -51.495 -174.000 -51.215 -173.720 ;
        RECT -50.565 -174.010 -50.285 -173.730 ;
        RECT -41.575 -174.000 -41.295 -173.720 ;
        RECT -40.645 -174.010 -40.365 -173.730 ;
        RECT -31.655 -174.000 -31.375 -173.720 ;
        RECT -30.725 -174.010 -30.445 -173.730 ;
        RECT -21.735 -174.000 -21.455 -173.720 ;
        RECT -20.805 -174.010 -20.525 -173.730 ;
        RECT -11.815 -174.000 -11.535 -173.720 ;
        RECT -10.885 -174.010 -10.605 -173.730 ;
        RECT -1.895 -174.000 -1.615 -173.720 ;
        RECT -0.965 -174.010 -0.685 -173.730 ;
        RECT 8.025 -174.000 8.305 -173.720 ;
        RECT 8.955 -174.010 9.235 -173.730 ;
        RECT 17.945 -174.000 18.225 -173.720 ;
        RECT 18.875 -174.010 19.155 -173.730 ;
        RECT 27.865 -174.000 28.145 -173.720 ;
        RECT -284.315 -175.490 -284.035 -175.210 ;
        RECT -274.395 -175.490 -274.115 -175.210 ;
        RECT -264.475 -175.490 -264.195 -175.210 ;
        RECT -254.555 -175.490 -254.275 -175.210 ;
        RECT -244.635 -175.490 -244.355 -175.210 ;
        RECT -234.715 -175.490 -234.435 -175.210 ;
        RECT -224.795 -175.490 -224.515 -175.210 ;
        RECT -214.875 -175.490 -214.595 -175.210 ;
        RECT -204.955 -175.490 -204.675 -175.210 ;
        RECT -195.035 -175.490 -194.755 -175.210 ;
        RECT -185.115 -175.490 -184.835 -175.210 ;
        RECT -175.195 -175.490 -174.915 -175.210 ;
        RECT -165.275 -175.490 -164.995 -175.210 ;
        RECT -155.355 -175.490 -155.075 -175.210 ;
        RECT -145.435 -175.490 -145.155 -175.210 ;
        RECT -135.515 -175.490 -135.235 -175.210 ;
        RECT -125.595 -175.490 -125.315 -175.210 ;
        RECT -115.675 -175.490 -115.395 -175.210 ;
        RECT -105.755 -175.490 -105.475 -175.210 ;
        RECT -95.835 -175.490 -95.555 -175.210 ;
        RECT -85.915 -175.490 -85.635 -175.210 ;
        RECT -75.995 -175.490 -75.715 -175.210 ;
        RECT -66.075 -175.490 -65.795 -175.210 ;
        RECT -56.155 -175.490 -55.875 -175.210 ;
        RECT -46.235 -175.490 -45.955 -175.210 ;
        RECT -36.315 -175.490 -36.035 -175.210 ;
        RECT -26.395 -175.490 -26.115 -175.210 ;
        RECT -16.475 -175.490 -16.195 -175.210 ;
        RECT -6.555 -175.490 -6.275 -175.210 ;
        RECT 3.365 -175.490 3.645 -175.210 ;
        RECT 13.285 -175.490 13.565 -175.210 ;
        RECT 23.205 -175.490 23.485 -175.210 ;
        RECT -279.275 -178.350 -278.995 -178.070 ;
        RECT -269.355 -178.350 -269.075 -178.070 ;
        RECT -259.435 -178.350 -259.155 -178.070 ;
        RECT -249.515 -178.350 -249.235 -178.070 ;
        RECT -239.595 -178.350 -239.315 -178.070 ;
        RECT -229.675 -178.350 -229.395 -178.070 ;
        RECT -219.755 -178.350 -219.475 -178.070 ;
        RECT -209.835 -178.350 -209.555 -178.070 ;
        RECT -199.915 -178.350 -199.635 -178.070 ;
        RECT -189.995 -178.350 -189.715 -178.070 ;
        RECT -180.075 -178.350 -179.795 -178.070 ;
        RECT -170.155 -178.350 -169.875 -178.070 ;
        RECT -160.235 -178.350 -159.955 -178.070 ;
        RECT -150.315 -178.350 -150.035 -178.070 ;
        RECT -140.395 -178.350 -140.115 -178.070 ;
        RECT -130.475 -178.350 -130.195 -178.070 ;
        RECT -120.555 -178.350 -120.275 -178.070 ;
        RECT -110.635 -178.350 -110.355 -178.070 ;
        RECT -100.715 -178.350 -100.435 -178.070 ;
        RECT -90.795 -178.350 -90.515 -178.070 ;
        RECT -80.875 -178.350 -80.595 -178.070 ;
        RECT -70.955 -178.350 -70.675 -178.070 ;
        RECT -61.035 -178.350 -60.755 -178.070 ;
        RECT -51.115 -178.350 -50.835 -178.070 ;
        RECT -41.195 -178.350 -40.915 -178.070 ;
        RECT -31.275 -178.350 -30.995 -178.070 ;
        RECT -21.355 -178.350 -21.075 -178.070 ;
        RECT -11.435 -178.350 -11.155 -178.070 ;
        RECT -1.515 -178.350 -1.235 -178.070 ;
        RECT 8.405 -178.350 8.685 -178.070 ;
        RECT 18.325 -178.350 18.605 -178.070 ;
        RECT 28.245 -178.350 28.525 -178.070 ;
        RECT -284.615 -179.890 -284.335 -179.610 ;
        RECT -283.685 -179.890 -283.405 -179.610 ;
        RECT -274.695 -179.890 -274.415 -179.610 ;
        RECT -273.765 -179.890 -273.485 -179.610 ;
        RECT -264.775 -179.890 -264.495 -179.610 ;
        RECT -263.845 -179.890 -263.565 -179.610 ;
        RECT -254.855 -179.890 -254.575 -179.610 ;
        RECT -253.925 -179.890 -253.645 -179.610 ;
        RECT -244.935 -179.890 -244.655 -179.610 ;
        RECT -244.005 -179.890 -243.725 -179.610 ;
        RECT -235.015 -179.890 -234.735 -179.610 ;
        RECT -234.085 -179.890 -233.805 -179.610 ;
        RECT -225.095 -179.890 -224.815 -179.610 ;
        RECT -224.165 -179.890 -223.885 -179.610 ;
        RECT -215.175 -179.890 -214.895 -179.610 ;
        RECT -214.245 -179.890 -213.965 -179.610 ;
        RECT -205.255 -179.890 -204.975 -179.610 ;
        RECT -204.325 -179.890 -204.045 -179.610 ;
        RECT -195.335 -179.890 -195.055 -179.610 ;
        RECT -194.405 -179.890 -194.125 -179.610 ;
        RECT -185.415 -179.890 -185.135 -179.610 ;
        RECT -184.485 -179.890 -184.205 -179.610 ;
        RECT -175.495 -179.890 -175.215 -179.610 ;
        RECT -174.565 -179.890 -174.285 -179.610 ;
        RECT -165.575 -179.890 -165.295 -179.610 ;
        RECT -164.645 -179.890 -164.365 -179.610 ;
        RECT -155.655 -179.890 -155.375 -179.610 ;
        RECT -154.725 -179.890 -154.445 -179.610 ;
        RECT -145.735 -179.890 -145.455 -179.610 ;
        RECT -144.805 -179.890 -144.525 -179.610 ;
        RECT -135.815 -179.890 -135.535 -179.610 ;
        RECT -134.885 -179.890 -134.605 -179.610 ;
        RECT -125.895 -179.890 -125.615 -179.610 ;
        RECT -124.965 -179.890 -124.685 -179.610 ;
        RECT -115.975 -179.890 -115.695 -179.610 ;
        RECT -115.045 -179.890 -114.765 -179.610 ;
        RECT -106.055 -179.890 -105.775 -179.610 ;
        RECT -105.125 -179.890 -104.845 -179.610 ;
        RECT -96.135 -179.890 -95.855 -179.610 ;
        RECT -95.205 -179.890 -94.925 -179.610 ;
        RECT -86.215 -179.890 -85.935 -179.610 ;
        RECT -85.285 -179.890 -85.005 -179.610 ;
        RECT -76.295 -179.890 -76.015 -179.610 ;
        RECT -75.365 -179.890 -75.085 -179.610 ;
        RECT -66.375 -179.890 -66.095 -179.610 ;
        RECT -65.445 -179.890 -65.165 -179.610 ;
        RECT -56.455 -179.890 -56.175 -179.610 ;
        RECT -55.525 -179.890 -55.245 -179.610 ;
        RECT -46.535 -179.890 -46.255 -179.610 ;
        RECT -45.605 -179.890 -45.325 -179.610 ;
        RECT -36.615 -179.890 -36.335 -179.610 ;
        RECT -35.685 -179.890 -35.405 -179.610 ;
        RECT -26.695 -179.890 -26.415 -179.610 ;
        RECT -25.765 -179.890 -25.485 -179.610 ;
        RECT -16.775 -179.890 -16.495 -179.610 ;
        RECT -15.845 -179.890 -15.565 -179.610 ;
        RECT -6.855 -179.890 -6.575 -179.610 ;
        RECT -5.925 -179.890 -5.645 -179.610 ;
        RECT 3.065 -179.890 3.345 -179.610 ;
        RECT 3.995 -179.890 4.275 -179.610 ;
        RECT 12.985 -179.890 13.265 -179.610 ;
        RECT 13.915 -179.890 14.195 -179.610 ;
        RECT 22.905 -179.890 23.185 -179.610 ;
        RECT 23.835 -179.890 24.115 -179.610 ;
      LAYER met3 ;
        RECT -298.750 109.690 -293.660 109.870 ;
        RECT 29.330 109.690 34.420 109.750 ;
        RECT -298.750 100.060 34.420 109.690 ;
        RECT -298.750 82.780 -293.660 100.060 ;
        RECT -291.620 82.780 -290.850 100.060 ;
        RECT -286.660 89.210 -285.890 100.060 ;
        RECT -281.700 95.140 -280.930 100.060 ;
        RECT -282.020 94.730 -280.600 95.140 ;
        RECT -281.700 90.850 -280.930 94.730 ;
        RECT -281.910 90.370 -280.710 90.850 ;
        RECT -286.980 88.800 -285.560 89.210 ;
        RECT -286.660 82.780 -285.890 88.800 ;
        RECT -281.700 82.780 -280.930 90.370 ;
        RECT -276.760 89.210 -275.990 100.060 ;
        RECT -271.780 95.230 -271.010 100.060 ;
        RECT -271.780 95.140 -271.000 95.230 ;
        RECT -272.100 94.730 -270.680 95.140 ;
        RECT -271.780 92.780 -271.000 94.730 ;
        RECT -271.820 90.850 -271.000 92.780 ;
        RECT -271.990 90.370 -270.790 90.850 ;
        RECT -277.060 88.800 -275.640 89.210 ;
        RECT -271.820 88.880 -271.000 90.370 ;
        RECT -266.810 89.210 -266.040 100.060 ;
        RECT -261.820 95.140 -261.050 100.060 ;
        RECT -262.180 94.730 -260.760 95.140 ;
        RECT -261.820 90.850 -261.050 94.730 ;
        RECT -262.070 90.370 -260.870 90.850 ;
        RECT -276.760 82.780 -275.990 88.800 ;
        RECT -271.830 85.270 -271.000 88.880 ;
        RECT -267.140 88.800 -265.720 89.210 ;
        RECT -271.830 82.780 -271.010 85.270 ;
        RECT -266.810 82.780 -266.040 88.800 ;
        RECT -261.820 82.780 -261.050 90.370 ;
        RECT -256.920 89.210 -256.150 100.060 ;
        RECT -251.930 95.140 -251.160 100.060 ;
        RECT -252.260 94.730 -250.840 95.140 ;
        RECT -251.930 90.850 -251.160 94.730 ;
        RECT -252.150 90.370 -250.950 90.850 ;
        RECT -257.220 88.800 -255.800 89.210 ;
        RECT -256.920 82.780 -256.150 88.800 ;
        RECT -251.930 82.780 -251.160 90.370 ;
        RECT -246.990 89.210 -246.220 100.060 ;
        RECT -242.020 95.140 -241.250 100.060 ;
        RECT -242.340 94.730 -240.920 95.140 ;
        RECT -242.020 90.850 -241.250 94.730 ;
        RECT -242.230 90.370 -241.030 90.850 ;
        RECT -247.300 88.800 -245.880 89.210 ;
        RECT -246.990 82.780 -246.220 88.800 ;
        RECT -242.020 82.780 -241.250 90.370 ;
        RECT -237.080 89.210 -236.310 100.060 ;
        RECT -232.120 95.140 -231.350 100.060 ;
        RECT -232.420 94.730 -231.000 95.140 ;
        RECT -232.120 90.850 -231.350 94.730 ;
        RECT -232.310 90.370 -231.110 90.850 ;
        RECT -237.380 88.800 -235.960 89.210 ;
        RECT -237.080 82.780 -236.310 88.800 ;
        RECT -232.120 82.780 -231.350 90.370 ;
        RECT -227.150 89.210 -226.380 100.060 ;
        RECT -222.180 95.140 -221.410 100.060 ;
        RECT -222.500 94.730 -221.080 95.140 ;
        RECT -222.180 90.850 -221.410 94.730 ;
        RECT -222.390 90.370 -221.190 90.850 ;
        RECT -227.460 88.800 -226.040 89.210 ;
        RECT -227.150 82.780 -226.380 88.800 ;
        RECT -222.180 82.780 -221.410 90.370 ;
        RECT -217.200 89.210 -216.430 100.060 ;
        RECT -212.240 95.140 -211.470 100.060 ;
        RECT -212.580 94.730 -211.160 95.140 ;
        RECT -212.240 90.850 -211.470 94.730 ;
        RECT -212.470 90.370 -211.270 90.850 ;
        RECT -217.540 88.800 -216.120 89.210 ;
        RECT -217.200 82.780 -216.430 88.800 ;
        RECT -212.240 82.780 -211.470 90.370 ;
        RECT -207.290 89.210 -206.520 100.060 ;
        RECT -202.350 95.140 -201.580 100.060 ;
        RECT -202.660 94.730 -201.240 95.140 ;
        RECT -202.350 90.850 -201.580 94.730 ;
        RECT -202.550 90.370 -201.350 90.850 ;
        RECT -207.620 88.800 -206.200 89.210 ;
        RECT -207.290 82.780 -206.520 88.800 ;
        RECT -202.350 82.780 -201.580 90.370 ;
        RECT -197.420 89.210 -196.650 100.060 ;
        RECT -192.420 95.140 -191.650 100.060 ;
        RECT -192.740 94.730 -191.320 95.140 ;
        RECT -192.420 90.850 -191.650 94.730 ;
        RECT -192.630 90.370 -191.430 90.850 ;
        RECT -197.700 88.800 -196.280 89.210 ;
        RECT -197.420 82.780 -196.650 88.800 ;
        RECT -192.420 82.780 -191.650 90.370 ;
        RECT -187.460 89.210 -186.690 100.060 ;
        RECT -182.510 95.140 -181.740 100.060 ;
        RECT -182.820 94.730 -181.400 95.140 ;
        RECT -182.510 90.850 -181.740 94.730 ;
        RECT -182.710 90.370 -181.510 90.850 ;
        RECT -187.780 88.800 -186.360 89.210 ;
        RECT -187.460 82.780 -186.690 88.800 ;
        RECT -182.510 82.780 -181.740 90.370 ;
        RECT -177.550 89.210 -176.780 100.060 ;
        RECT -172.560 95.140 -171.790 100.060 ;
        RECT -172.900 94.730 -171.480 95.140 ;
        RECT -172.560 90.850 -171.790 94.730 ;
        RECT -172.790 90.370 -171.590 90.850 ;
        RECT -177.860 88.800 -176.440 89.210 ;
        RECT -177.550 82.780 -176.780 88.800 ;
        RECT -172.560 82.780 -171.790 90.370 ;
        RECT -167.620 89.210 -166.850 100.060 ;
        RECT -162.620 95.140 -161.850 100.060 ;
        RECT -162.980 94.730 -161.560 95.140 ;
        RECT -162.620 90.850 -161.850 94.730 ;
        RECT -162.870 90.370 -161.670 90.850 ;
        RECT -167.940 88.800 -166.520 89.210 ;
        RECT -167.620 82.780 -166.850 88.800 ;
        RECT -162.620 82.780 -161.850 90.370 ;
        RECT -157.710 89.210 -156.940 100.060 ;
        RECT -152.760 95.140 -151.990 100.060 ;
        RECT -153.060 94.730 -151.640 95.140 ;
        RECT -152.760 90.850 -151.990 94.730 ;
        RECT -152.950 90.370 -151.750 90.850 ;
        RECT -158.020 88.800 -156.600 89.210 ;
        RECT -157.710 82.780 -156.940 88.800 ;
        RECT -152.760 82.780 -151.990 90.370 ;
        RECT -147.790 89.210 -147.020 100.060 ;
        RECT -142.830 95.140 -142.060 100.060 ;
        RECT -143.140 94.730 -141.720 95.140 ;
        RECT -142.830 90.850 -142.060 94.730 ;
        RECT -143.030 90.370 -141.830 90.850 ;
        RECT -148.100 88.800 -146.680 89.210 ;
        RECT -147.790 82.780 -147.020 88.800 ;
        RECT -142.830 82.780 -142.060 90.370 ;
        RECT -137.850 89.210 -137.080 100.060 ;
        RECT -132.920 95.140 -132.150 100.060 ;
        RECT -133.220 94.730 -131.800 95.140 ;
        RECT -132.920 90.850 -132.150 94.730 ;
        RECT -133.110 90.370 -131.910 90.850 ;
        RECT -138.180 88.800 -136.760 89.210 ;
        RECT -137.850 82.780 -137.080 88.800 ;
        RECT -132.920 82.780 -132.150 90.370 ;
        RECT -127.940 89.210 -127.170 100.060 ;
        RECT -122.960 95.140 -122.190 100.060 ;
        RECT -123.300 94.730 -121.880 95.140 ;
        RECT -122.960 90.850 -122.190 94.730 ;
        RECT -123.190 90.370 -121.990 90.850 ;
        RECT -128.260 88.800 -126.840 89.210 ;
        RECT -127.940 82.780 -127.170 88.800 ;
        RECT -122.960 82.780 -122.190 90.370 ;
        RECT -118.040 89.210 -117.270 100.060 ;
        RECT -113.080 95.140 -112.310 100.060 ;
        RECT -113.380 94.730 -111.960 95.140 ;
        RECT -113.080 90.850 -112.310 94.730 ;
        RECT -113.270 90.370 -112.070 90.850 ;
        RECT -118.340 88.800 -116.920 89.210 ;
        RECT -118.040 82.780 -117.270 88.800 ;
        RECT -113.080 82.780 -112.310 90.370 ;
        RECT -108.110 89.210 -107.340 100.060 ;
        RECT -103.150 95.140 -102.380 100.060 ;
        RECT -103.460 94.730 -102.040 95.140 ;
        RECT -103.150 90.850 -102.380 94.730 ;
        RECT -103.350 90.370 -102.150 90.850 ;
        RECT -108.420 88.800 -107.000 89.210 ;
        RECT -108.110 82.780 -107.340 88.800 ;
        RECT -103.150 82.780 -102.380 90.370 ;
        RECT -98.160 89.210 -97.390 100.060 ;
        RECT -93.210 95.140 -92.440 100.060 ;
        RECT -93.540 94.730 -92.120 95.140 ;
        RECT -93.210 90.850 -92.440 94.730 ;
        RECT -93.430 90.370 -92.230 90.850 ;
        RECT -98.500 88.800 -97.080 89.210 ;
        RECT -98.160 82.780 -97.390 88.800 ;
        RECT -93.210 82.780 -92.440 90.370 ;
        RECT -88.260 89.210 -87.490 100.060 ;
        RECT -83.270 95.140 -82.500 100.060 ;
        RECT -83.620 94.730 -82.200 95.140 ;
        RECT -83.270 90.850 -82.500 94.730 ;
        RECT -83.510 90.370 -82.310 90.850 ;
        RECT -88.580 88.800 -87.160 89.210 ;
        RECT -88.260 82.780 -87.490 88.800 ;
        RECT -83.270 82.780 -82.500 90.370 ;
        RECT -78.350 89.210 -77.580 100.060 ;
        RECT -73.390 95.140 -72.620 100.060 ;
        RECT -73.700 94.730 -72.280 95.140 ;
        RECT -73.390 90.850 -72.620 94.730 ;
        RECT -73.590 90.370 -72.390 90.850 ;
        RECT -78.660 88.800 -77.240 89.210 ;
        RECT -78.350 82.780 -77.580 88.800 ;
        RECT -73.390 82.780 -72.620 90.370 ;
        RECT -68.410 89.210 -67.640 100.060 ;
        RECT -63.430 95.140 -62.660 100.060 ;
        RECT -63.780 94.730 -62.360 95.140 ;
        RECT -63.430 90.850 -62.660 94.730 ;
        RECT -63.670 90.370 -62.470 90.850 ;
        RECT -68.740 88.800 -67.320 89.210 ;
        RECT -68.410 82.780 -67.640 88.800 ;
        RECT -63.430 82.780 -62.660 90.370 ;
        RECT -58.520 89.210 -57.750 100.060 ;
        RECT -53.520 95.140 -52.750 100.060 ;
        RECT -53.860 94.730 -52.440 95.140 ;
        RECT -53.520 90.850 -52.750 94.730 ;
        RECT -53.750 90.370 -52.550 90.850 ;
        RECT -58.820 88.800 -57.400 89.210 ;
        RECT -58.520 82.780 -57.750 88.800 ;
        RECT -53.520 82.780 -52.750 90.370 ;
        RECT -48.560 89.210 -47.790 100.060 ;
        RECT -43.630 95.140 -42.860 100.060 ;
        RECT -43.940 94.730 -42.520 95.140 ;
        RECT -43.630 90.850 -42.860 94.730 ;
        RECT -43.830 90.370 -42.630 90.850 ;
        RECT -48.900 88.800 -47.480 89.210 ;
        RECT -48.560 82.780 -47.790 88.800 ;
        RECT -43.630 82.780 -42.860 90.370 ;
        RECT -38.680 89.210 -37.910 100.060 ;
        RECT -33.700 95.140 -32.930 100.060 ;
        RECT -34.020 94.730 -32.600 95.140 ;
        RECT -33.700 90.850 -32.930 94.730 ;
        RECT -33.910 90.370 -32.710 90.850 ;
        RECT -38.980 88.800 -37.560 89.210 ;
        RECT -38.680 82.780 -37.910 88.800 ;
        RECT -33.700 82.780 -32.930 90.370 ;
        RECT -28.750 89.210 -27.980 100.060 ;
        RECT -23.800 95.140 -23.030 100.060 ;
        RECT -24.100 94.730 -22.680 95.140 ;
        RECT -23.800 90.850 -23.030 94.730 ;
        RECT -23.990 90.370 -22.790 90.850 ;
        RECT -29.060 88.800 -27.640 89.210 ;
        RECT -28.750 82.780 -27.980 88.800 ;
        RECT -23.800 82.780 -23.030 90.370 ;
        RECT -18.820 89.210 -18.050 100.060 ;
        RECT -13.870 95.140 -13.100 100.060 ;
        RECT -14.180 94.730 -12.760 95.140 ;
        RECT -13.870 90.850 -13.100 94.730 ;
        RECT -14.070 90.370 -12.870 90.850 ;
        RECT -19.140 88.800 -17.720 89.210 ;
        RECT -18.820 82.780 -18.050 88.800 ;
        RECT -13.870 82.780 -13.100 90.370 ;
        RECT -8.920 89.210 -8.150 100.060 ;
        RECT -3.940 95.140 -3.170 100.060 ;
        RECT -4.260 94.730 -2.840 95.140 ;
        RECT -3.940 90.850 -3.170 94.730 ;
        RECT -4.150 90.370 -2.950 90.850 ;
        RECT -9.220 88.800 -7.800 89.210 ;
        RECT -8.920 82.780 -8.150 88.800 ;
        RECT -3.940 82.780 -3.170 90.370 ;
        RECT 1.010 89.210 1.780 100.060 ;
        RECT 5.940 95.140 6.710 100.060 ;
        RECT 5.660 94.730 7.080 95.140 ;
        RECT 5.940 90.850 6.710 94.730 ;
        RECT 5.770 90.370 6.970 90.850 ;
        RECT 0.700 88.800 2.120 89.210 ;
        RECT 1.010 82.780 1.780 88.800 ;
        RECT 5.940 82.780 6.710 90.370 ;
        RECT 10.940 89.210 11.710 100.060 ;
        RECT 15.890 95.140 16.660 100.060 ;
        RECT 15.580 94.730 17.000 95.140 ;
        RECT 15.890 90.850 16.660 94.730 ;
        RECT 15.690 90.370 16.890 90.850 ;
        RECT 10.620 88.800 12.040 89.210 ;
        RECT 10.940 82.780 11.710 88.800 ;
        RECT 15.890 82.780 16.660 90.370 ;
        RECT 20.870 89.210 21.640 100.060 ;
        RECT 25.880 95.140 26.650 100.060 ;
        RECT 25.500 94.730 26.650 95.140 ;
        RECT 25.880 90.850 26.650 94.730 ;
        RECT 25.610 90.370 26.440 90.850 ;
        RECT 20.540 88.800 21.960 89.210 ;
        RECT 20.870 82.780 21.640 88.800 ;
        RECT 25.880 82.780 26.650 90.370 ;
        RECT 29.330 83.200 34.420 100.060 ;
        RECT 27.700 83.150 164.350 83.200 ;
        RECT 27.700 82.780 165.390 83.150 ;
        RECT -298.750 73.570 165.390 82.780 ;
        RECT -298.750 73.150 34.420 73.570 ;
        RECT -298.750 73.140 -293.660 73.150 ;
        RECT -298.500 21.980 -293.410 22.160 ;
        RECT -245.790 21.980 -216.050 73.150 ;
        RECT 29.330 73.020 34.420 73.150 ;
        RECT 29.580 21.980 34.670 22.040 ;
        RECT -298.500 12.350 34.670 21.980 ;
        RECT -298.500 -4.930 -293.410 12.350 ;
        RECT -291.370 -4.930 -290.600 12.350 ;
        RECT -286.410 1.500 -285.640 12.350 ;
        RECT -281.450 7.430 -280.680 12.350 ;
        RECT -281.770 7.020 -280.350 7.430 ;
        RECT -281.450 3.140 -280.680 7.020 ;
        RECT -281.660 2.660 -280.460 3.140 ;
        RECT -286.730 1.090 -285.310 1.500 ;
        RECT -286.410 -4.930 -285.640 1.090 ;
        RECT -281.450 -4.930 -280.680 2.660 ;
        RECT -276.510 1.500 -275.740 12.350 ;
        RECT -271.530 7.520 -270.760 12.350 ;
        RECT -271.530 7.430 -270.750 7.520 ;
        RECT -271.850 7.020 -270.430 7.430 ;
        RECT -271.530 5.070 -270.750 7.020 ;
        RECT -271.570 3.140 -270.750 5.070 ;
        RECT -271.740 2.660 -270.540 3.140 ;
        RECT -276.810 1.090 -275.390 1.500 ;
        RECT -271.570 1.170 -270.750 2.660 ;
        RECT -266.560 1.500 -265.790 12.350 ;
        RECT -261.570 7.430 -260.800 12.350 ;
        RECT -261.930 7.020 -260.510 7.430 ;
        RECT -261.570 3.140 -260.800 7.020 ;
        RECT -261.820 2.660 -260.620 3.140 ;
        RECT -276.510 -4.930 -275.740 1.090 ;
        RECT -271.580 -2.440 -270.750 1.170 ;
        RECT -266.890 1.090 -265.470 1.500 ;
        RECT -271.580 -4.930 -270.760 -2.440 ;
        RECT -266.560 -4.930 -265.790 1.090 ;
        RECT -261.570 -4.930 -260.800 2.660 ;
        RECT -256.670 1.500 -255.900 12.350 ;
        RECT -251.680 7.430 -250.910 12.350 ;
        RECT -252.010 7.020 -250.590 7.430 ;
        RECT -251.680 3.140 -250.910 7.020 ;
        RECT -251.900 2.660 -250.700 3.140 ;
        RECT -256.970 1.090 -255.550 1.500 ;
        RECT -256.670 -4.930 -255.900 1.090 ;
        RECT -251.680 -4.930 -250.910 2.660 ;
        RECT -246.740 1.500 -245.970 12.350 ;
        RECT -241.770 7.430 -241.000 12.350 ;
        RECT -242.090 7.020 -240.670 7.430 ;
        RECT -241.770 3.140 -241.000 7.020 ;
        RECT -241.980 2.660 -240.780 3.140 ;
        RECT -247.050 1.090 -245.630 1.500 ;
        RECT -246.740 -4.930 -245.970 1.090 ;
        RECT -241.770 -4.930 -241.000 2.660 ;
        RECT -236.830 1.500 -236.060 12.350 ;
        RECT -231.870 7.430 -231.100 12.350 ;
        RECT -232.170 7.020 -230.750 7.430 ;
        RECT -231.870 3.140 -231.100 7.020 ;
        RECT -232.060 2.660 -230.860 3.140 ;
        RECT -237.130 1.090 -235.710 1.500 ;
        RECT -236.830 -4.930 -236.060 1.090 ;
        RECT -231.870 -4.930 -231.100 2.660 ;
        RECT -226.900 1.500 -226.130 12.350 ;
        RECT -221.930 7.430 -221.160 12.350 ;
        RECT -222.250 7.020 -220.830 7.430 ;
        RECT -221.930 3.140 -221.160 7.020 ;
        RECT -222.140 2.660 -220.940 3.140 ;
        RECT -227.210 1.090 -225.790 1.500 ;
        RECT -226.900 -4.930 -226.130 1.090 ;
        RECT -221.930 -4.930 -221.160 2.660 ;
        RECT -216.950 1.500 -216.180 12.350 ;
        RECT -211.990 7.430 -211.220 12.350 ;
        RECT -212.330 7.020 -210.910 7.430 ;
        RECT -211.990 3.140 -211.220 7.020 ;
        RECT -212.220 2.660 -211.020 3.140 ;
        RECT -217.290 1.090 -215.870 1.500 ;
        RECT -216.950 -4.930 -216.180 1.090 ;
        RECT -211.990 -4.930 -211.220 2.660 ;
        RECT -207.040 1.500 -206.270 12.350 ;
        RECT -202.100 7.430 -201.330 12.350 ;
        RECT -202.410 7.020 -200.990 7.430 ;
        RECT -202.100 3.140 -201.330 7.020 ;
        RECT -202.300 2.660 -201.100 3.140 ;
        RECT -207.370 1.090 -205.950 1.500 ;
        RECT -207.040 -4.930 -206.270 1.090 ;
        RECT -202.100 -4.930 -201.330 2.660 ;
        RECT -197.170 1.500 -196.400 12.350 ;
        RECT -192.170 7.430 -191.400 12.350 ;
        RECT -192.490 7.020 -191.070 7.430 ;
        RECT -192.170 3.140 -191.400 7.020 ;
        RECT -192.380 2.660 -191.180 3.140 ;
        RECT -197.450 1.090 -196.030 1.500 ;
        RECT -197.170 -4.930 -196.400 1.090 ;
        RECT -192.170 -4.930 -191.400 2.660 ;
        RECT -187.210 1.500 -186.440 12.350 ;
        RECT -182.260 7.430 -181.490 12.350 ;
        RECT -182.570 7.020 -181.150 7.430 ;
        RECT -182.260 3.140 -181.490 7.020 ;
        RECT -182.460 2.660 -181.260 3.140 ;
        RECT -187.530 1.090 -186.110 1.500 ;
        RECT -187.210 -4.930 -186.440 1.090 ;
        RECT -182.260 -4.930 -181.490 2.660 ;
        RECT -177.300 1.500 -176.530 12.350 ;
        RECT -172.310 7.430 -171.540 12.350 ;
        RECT -172.650 7.020 -171.230 7.430 ;
        RECT -172.310 3.140 -171.540 7.020 ;
        RECT -172.540 2.660 -171.340 3.140 ;
        RECT -177.610 1.090 -176.190 1.500 ;
        RECT -177.300 -4.930 -176.530 1.090 ;
        RECT -172.310 -4.930 -171.540 2.660 ;
        RECT -167.370 1.500 -166.600 12.350 ;
        RECT -162.370 7.430 -161.600 12.350 ;
        RECT -162.730 7.020 -161.310 7.430 ;
        RECT -162.370 3.140 -161.600 7.020 ;
        RECT -162.620 2.660 -161.420 3.140 ;
        RECT -167.690 1.090 -166.270 1.500 ;
        RECT -167.370 -4.930 -166.600 1.090 ;
        RECT -162.370 -4.930 -161.600 2.660 ;
        RECT -157.460 1.500 -156.690 12.350 ;
        RECT -152.510 7.430 -151.740 12.350 ;
        RECT -152.810 7.020 -151.390 7.430 ;
        RECT -152.510 3.140 -151.740 7.020 ;
        RECT -152.700 2.660 -151.500 3.140 ;
        RECT -157.770 1.090 -156.350 1.500 ;
        RECT -157.460 -4.930 -156.690 1.090 ;
        RECT -152.510 -4.930 -151.740 2.660 ;
        RECT -147.540 1.500 -146.770 12.350 ;
        RECT -142.580 7.430 -141.810 12.350 ;
        RECT -142.890 7.020 -141.470 7.430 ;
        RECT -142.580 3.140 -141.810 7.020 ;
        RECT -142.780 2.660 -141.580 3.140 ;
        RECT -147.850 1.090 -146.430 1.500 ;
        RECT -147.540 -4.930 -146.770 1.090 ;
        RECT -142.580 -4.930 -141.810 2.660 ;
        RECT -137.600 1.500 -136.830 12.350 ;
        RECT -132.670 7.430 -131.900 12.350 ;
        RECT -132.970 7.020 -131.550 7.430 ;
        RECT -132.670 3.140 -131.900 7.020 ;
        RECT -132.860 2.660 -131.660 3.140 ;
        RECT -137.930 1.090 -136.510 1.500 ;
        RECT -137.600 -4.930 -136.830 1.090 ;
        RECT -132.670 -4.930 -131.900 2.660 ;
        RECT -127.690 1.500 -126.920 12.350 ;
        RECT -122.710 7.430 -121.940 12.350 ;
        RECT -123.050 7.020 -121.630 7.430 ;
        RECT -122.710 3.140 -121.940 7.020 ;
        RECT -122.940 2.660 -121.740 3.140 ;
        RECT -128.010 1.090 -126.590 1.500 ;
        RECT -127.690 -4.930 -126.920 1.090 ;
        RECT -122.710 -4.930 -121.940 2.660 ;
        RECT -117.790 1.500 -117.020 12.350 ;
        RECT -112.830 7.430 -112.060 12.350 ;
        RECT -113.130 7.020 -111.710 7.430 ;
        RECT -112.830 3.140 -112.060 7.020 ;
        RECT -113.020 2.660 -111.820 3.140 ;
        RECT -118.090 1.090 -116.670 1.500 ;
        RECT -117.790 -4.930 -117.020 1.090 ;
        RECT -112.830 -4.930 -112.060 2.660 ;
        RECT -107.860 1.500 -107.090 12.350 ;
        RECT -102.900 7.430 -102.130 12.350 ;
        RECT -103.210 7.020 -101.790 7.430 ;
        RECT -102.900 3.140 -102.130 7.020 ;
        RECT -103.100 2.660 -101.900 3.140 ;
        RECT -108.170 1.090 -106.750 1.500 ;
        RECT -107.860 -4.930 -107.090 1.090 ;
        RECT -102.900 -4.930 -102.130 2.660 ;
        RECT -97.910 1.500 -97.140 12.350 ;
        RECT -92.960 7.430 -92.190 12.350 ;
        RECT -93.290 7.020 -91.870 7.430 ;
        RECT -92.960 3.140 -92.190 7.020 ;
        RECT -93.180 2.660 -91.980 3.140 ;
        RECT -98.250 1.090 -96.830 1.500 ;
        RECT -97.910 -4.930 -97.140 1.090 ;
        RECT -92.960 -4.930 -92.190 2.660 ;
        RECT -88.010 1.500 -87.240 12.350 ;
        RECT -83.020 7.430 -82.250 12.350 ;
        RECT -83.370 7.020 -81.950 7.430 ;
        RECT -83.020 3.140 -82.250 7.020 ;
        RECT -83.260 2.660 -82.060 3.140 ;
        RECT -88.330 1.090 -86.910 1.500 ;
        RECT -88.010 -4.930 -87.240 1.090 ;
        RECT -83.020 -4.930 -82.250 2.660 ;
        RECT -78.100 1.500 -77.330 12.350 ;
        RECT -73.140 7.430 -72.370 12.350 ;
        RECT -73.450 7.020 -72.030 7.430 ;
        RECT -73.140 3.140 -72.370 7.020 ;
        RECT -73.340 2.660 -72.140 3.140 ;
        RECT -78.410 1.090 -76.990 1.500 ;
        RECT -78.100 -4.930 -77.330 1.090 ;
        RECT -73.140 -4.930 -72.370 2.660 ;
        RECT -68.160 1.500 -67.390 12.350 ;
        RECT -63.180 7.430 -62.410 12.350 ;
        RECT -63.530 7.020 -62.110 7.430 ;
        RECT -63.180 3.140 -62.410 7.020 ;
        RECT -63.420 2.660 -62.220 3.140 ;
        RECT -68.490 1.090 -67.070 1.500 ;
        RECT -68.160 -4.930 -67.390 1.090 ;
        RECT -63.180 -4.930 -62.410 2.660 ;
        RECT -58.270 1.500 -57.500 12.350 ;
        RECT -53.270 7.430 -52.500 12.350 ;
        RECT -53.610 7.020 -52.190 7.430 ;
        RECT -53.270 3.140 -52.500 7.020 ;
        RECT -53.500 2.660 -52.300 3.140 ;
        RECT -58.570 1.090 -57.150 1.500 ;
        RECT -58.270 -4.930 -57.500 1.090 ;
        RECT -53.270 -4.930 -52.500 2.660 ;
        RECT -48.310 1.500 -47.540 12.350 ;
        RECT -43.380 7.430 -42.610 12.350 ;
        RECT -43.690 7.020 -42.270 7.430 ;
        RECT -43.380 3.140 -42.610 7.020 ;
        RECT -43.580 2.660 -42.380 3.140 ;
        RECT -48.650 1.090 -47.230 1.500 ;
        RECT -48.310 -4.930 -47.540 1.090 ;
        RECT -43.380 -4.930 -42.610 2.660 ;
        RECT -38.430 1.500 -37.660 12.350 ;
        RECT -33.450 7.430 -32.680 12.350 ;
        RECT -33.770 7.020 -32.350 7.430 ;
        RECT -33.450 3.140 -32.680 7.020 ;
        RECT -33.660 2.660 -32.460 3.140 ;
        RECT -38.730 1.090 -37.310 1.500 ;
        RECT -38.430 -4.930 -37.660 1.090 ;
        RECT -33.450 -4.930 -32.680 2.660 ;
        RECT -28.500 1.500 -27.730 12.350 ;
        RECT -23.550 7.430 -22.780 12.350 ;
        RECT -23.850 7.020 -22.430 7.430 ;
        RECT -23.550 3.140 -22.780 7.020 ;
        RECT -23.740 2.660 -22.540 3.140 ;
        RECT -28.810 1.090 -27.390 1.500 ;
        RECT -28.500 -4.930 -27.730 1.090 ;
        RECT -23.550 -4.930 -22.780 2.660 ;
        RECT -18.570 1.500 -17.800 12.350 ;
        RECT -13.620 7.430 -12.850 12.350 ;
        RECT -13.930 7.020 -12.510 7.430 ;
        RECT -13.620 3.140 -12.850 7.020 ;
        RECT -13.820 2.660 -12.620 3.140 ;
        RECT -18.890 1.090 -17.470 1.500 ;
        RECT -18.570 -4.930 -17.800 1.090 ;
        RECT -13.620 -4.930 -12.850 2.660 ;
        RECT -8.670 1.500 -7.900 12.350 ;
        RECT -3.690 7.430 -2.920 12.350 ;
        RECT -4.010 7.020 -2.590 7.430 ;
        RECT -3.690 3.140 -2.920 7.020 ;
        RECT -3.900 2.660 -2.700 3.140 ;
        RECT -8.970 1.090 -7.550 1.500 ;
        RECT -8.670 -4.930 -7.900 1.090 ;
        RECT -3.690 -4.930 -2.920 2.660 ;
        RECT 1.260 1.500 2.030 12.350 ;
        RECT 6.190 7.430 6.960 12.350 ;
        RECT 5.910 7.020 7.330 7.430 ;
        RECT 6.190 3.140 6.960 7.020 ;
        RECT 6.020 2.660 7.220 3.140 ;
        RECT 0.950 1.090 2.370 1.500 ;
        RECT 1.260 -4.930 2.030 1.090 ;
        RECT 6.190 -4.930 6.960 2.660 ;
        RECT 11.190 1.500 11.960 12.350 ;
        RECT 16.140 7.430 16.910 12.350 ;
        RECT 15.830 7.020 17.250 7.430 ;
        RECT 16.140 3.140 16.910 7.020 ;
        RECT 15.940 2.660 17.140 3.140 ;
        RECT 10.870 1.090 12.290 1.500 ;
        RECT 11.190 -4.930 11.960 1.090 ;
        RECT 16.140 -4.930 16.910 2.660 ;
        RECT 21.120 1.500 21.890 12.350 ;
        RECT 26.130 7.430 26.900 12.350 ;
        RECT 25.750 7.020 26.900 7.430 ;
        RECT 26.130 3.140 26.900 7.020 ;
        RECT 25.860 2.660 26.690 3.140 ;
        RECT 20.790 1.090 22.210 1.500 ;
        RECT 21.120 -4.930 21.890 1.090 ;
        RECT 26.130 -4.930 26.900 2.660 ;
        RECT 29.580 -4.510 34.670 12.350 ;
        RECT 138.320 -4.510 165.390 73.570 ;
        RECT 27.950 -4.930 165.390 -4.510 ;
        RECT -298.500 -14.140 165.390 -4.930 ;
        RECT -298.500 -14.560 34.670 -14.140 ;
        RECT -298.500 -14.570 -293.410 -14.560 ;
        RECT -296.740 -71.370 -291.650 -71.190 ;
        RECT -176.260 -71.370 -146.520 -14.560 ;
        RECT 29.580 -14.690 34.670 -14.560 ;
        RECT 31.340 -71.370 36.430 -71.310 ;
        RECT -296.740 -81.000 36.430 -71.370 ;
        RECT -296.740 -98.280 -291.650 -81.000 ;
        RECT -289.610 -98.280 -288.840 -81.000 ;
        RECT -284.650 -91.850 -283.880 -81.000 ;
        RECT -279.690 -85.920 -278.920 -81.000 ;
        RECT -280.010 -86.330 -278.590 -85.920 ;
        RECT -279.690 -90.210 -278.920 -86.330 ;
        RECT -279.900 -90.690 -278.700 -90.210 ;
        RECT -284.970 -92.260 -283.550 -91.850 ;
        RECT -284.650 -98.280 -283.880 -92.260 ;
        RECT -279.690 -98.280 -278.920 -90.690 ;
        RECT -274.750 -91.850 -273.980 -81.000 ;
        RECT -269.770 -85.830 -269.000 -81.000 ;
        RECT -269.770 -85.920 -268.990 -85.830 ;
        RECT -270.090 -86.330 -268.670 -85.920 ;
        RECT -269.770 -88.280 -268.990 -86.330 ;
        RECT -269.810 -90.210 -268.990 -88.280 ;
        RECT -269.980 -90.690 -268.780 -90.210 ;
        RECT -275.050 -92.260 -273.630 -91.850 ;
        RECT -269.810 -92.180 -268.990 -90.690 ;
        RECT -264.800 -91.850 -264.030 -81.000 ;
        RECT -259.810 -85.920 -259.040 -81.000 ;
        RECT -260.170 -86.330 -258.750 -85.920 ;
        RECT -259.810 -90.210 -259.040 -86.330 ;
        RECT -260.060 -90.690 -258.860 -90.210 ;
        RECT -274.750 -98.280 -273.980 -92.260 ;
        RECT -269.820 -95.790 -268.990 -92.180 ;
        RECT -265.130 -92.260 -263.710 -91.850 ;
        RECT -269.820 -98.280 -269.000 -95.790 ;
        RECT -264.800 -98.280 -264.030 -92.260 ;
        RECT -259.810 -98.280 -259.040 -90.690 ;
        RECT -254.910 -91.850 -254.140 -81.000 ;
        RECT -249.920 -85.920 -249.150 -81.000 ;
        RECT -250.250 -86.330 -248.830 -85.920 ;
        RECT -249.920 -90.210 -249.150 -86.330 ;
        RECT -250.140 -90.690 -248.940 -90.210 ;
        RECT -255.210 -92.260 -253.790 -91.850 ;
        RECT -254.910 -98.280 -254.140 -92.260 ;
        RECT -249.920 -98.280 -249.150 -90.690 ;
        RECT -244.980 -91.850 -244.210 -81.000 ;
        RECT -240.010 -85.920 -239.240 -81.000 ;
        RECT -240.330 -86.330 -238.910 -85.920 ;
        RECT -240.010 -90.210 -239.240 -86.330 ;
        RECT -240.220 -90.690 -239.020 -90.210 ;
        RECT -245.290 -92.260 -243.870 -91.850 ;
        RECT -244.980 -98.280 -244.210 -92.260 ;
        RECT -240.010 -98.280 -239.240 -90.690 ;
        RECT -235.070 -91.850 -234.300 -81.000 ;
        RECT -230.110 -85.920 -229.340 -81.000 ;
        RECT -230.410 -86.330 -228.990 -85.920 ;
        RECT -230.110 -90.210 -229.340 -86.330 ;
        RECT -230.300 -90.690 -229.100 -90.210 ;
        RECT -235.370 -92.260 -233.950 -91.850 ;
        RECT -235.070 -98.280 -234.300 -92.260 ;
        RECT -230.110 -98.280 -229.340 -90.690 ;
        RECT -225.140 -91.850 -224.370 -81.000 ;
        RECT -220.170 -85.920 -219.400 -81.000 ;
        RECT -220.490 -86.330 -219.070 -85.920 ;
        RECT -220.170 -90.210 -219.400 -86.330 ;
        RECT -220.380 -90.690 -219.180 -90.210 ;
        RECT -225.450 -92.260 -224.030 -91.850 ;
        RECT -225.140 -98.280 -224.370 -92.260 ;
        RECT -220.170 -98.280 -219.400 -90.690 ;
        RECT -215.190 -91.850 -214.420 -81.000 ;
        RECT -210.230 -85.920 -209.460 -81.000 ;
        RECT -210.570 -86.330 -209.150 -85.920 ;
        RECT -210.230 -90.210 -209.460 -86.330 ;
        RECT -210.460 -90.690 -209.260 -90.210 ;
        RECT -215.530 -92.260 -214.110 -91.850 ;
        RECT -215.190 -98.280 -214.420 -92.260 ;
        RECT -210.230 -98.280 -209.460 -90.690 ;
        RECT -205.280 -91.850 -204.510 -81.000 ;
        RECT -200.340 -85.920 -199.570 -81.000 ;
        RECT -200.650 -86.330 -199.230 -85.920 ;
        RECT -200.340 -90.210 -199.570 -86.330 ;
        RECT -200.540 -90.690 -199.340 -90.210 ;
        RECT -205.610 -92.260 -204.190 -91.850 ;
        RECT -205.280 -98.280 -204.510 -92.260 ;
        RECT -200.340 -98.280 -199.570 -90.690 ;
        RECT -195.410 -91.850 -194.640 -81.000 ;
        RECT -190.410 -85.920 -189.640 -81.000 ;
        RECT -190.730 -86.330 -189.310 -85.920 ;
        RECT -190.410 -90.210 -189.640 -86.330 ;
        RECT -190.620 -90.690 -189.420 -90.210 ;
        RECT -195.690 -92.260 -194.270 -91.850 ;
        RECT -195.410 -98.280 -194.640 -92.260 ;
        RECT -190.410 -98.280 -189.640 -90.690 ;
        RECT -185.450 -91.850 -184.680 -81.000 ;
        RECT -180.500 -85.920 -179.730 -81.000 ;
        RECT -180.810 -86.330 -179.390 -85.920 ;
        RECT -180.500 -90.210 -179.730 -86.330 ;
        RECT -180.700 -90.690 -179.500 -90.210 ;
        RECT -185.770 -92.260 -184.350 -91.850 ;
        RECT -185.450 -98.280 -184.680 -92.260 ;
        RECT -180.500 -98.280 -179.730 -90.690 ;
        RECT -175.540 -91.850 -174.770 -81.000 ;
        RECT -170.550 -85.920 -169.780 -81.000 ;
        RECT -170.890 -86.330 -169.470 -85.920 ;
        RECT -170.550 -90.210 -169.780 -86.330 ;
        RECT -170.780 -90.690 -169.580 -90.210 ;
        RECT -175.850 -92.260 -174.430 -91.850 ;
        RECT -175.540 -98.280 -174.770 -92.260 ;
        RECT -170.550 -98.280 -169.780 -90.690 ;
        RECT -165.610 -91.850 -164.840 -81.000 ;
        RECT -160.610 -85.920 -159.840 -81.000 ;
        RECT -160.970 -86.330 -159.550 -85.920 ;
        RECT -160.610 -90.210 -159.840 -86.330 ;
        RECT -160.860 -90.690 -159.660 -90.210 ;
        RECT -165.930 -92.260 -164.510 -91.850 ;
        RECT -165.610 -98.280 -164.840 -92.260 ;
        RECT -160.610 -98.280 -159.840 -90.690 ;
        RECT -155.700 -91.850 -154.930 -81.000 ;
        RECT -150.750 -85.920 -149.980 -81.000 ;
        RECT -151.050 -86.330 -149.630 -85.920 ;
        RECT -150.750 -90.210 -149.980 -86.330 ;
        RECT -150.940 -90.690 -149.740 -90.210 ;
        RECT -156.010 -92.260 -154.590 -91.850 ;
        RECT -155.700 -98.280 -154.930 -92.260 ;
        RECT -150.750 -98.280 -149.980 -90.690 ;
        RECT -145.780 -91.850 -145.010 -81.000 ;
        RECT -140.820 -85.920 -140.050 -81.000 ;
        RECT -141.130 -86.330 -139.710 -85.920 ;
        RECT -140.820 -90.210 -140.050 -86.330 ;
        RECT -141.020 -90.690 -139.820 -90.210 ;
        RECT -146.090 -92.260 -144.670 -91.850 ;
        RECT -145.780 -98.280 -145.010 -92.260 ;
        RECT -140.820 -98.280 -140.050 -90.690 ;
        RECT -135.840 -91.850 -135.070 -81.000 ;
        RECT -130.910 -85.920 -130.140 -81.000 ;
        RECT -131.210 -86.330 -129.790 -85.920 ;
        RECT -130.910 -90.210 -130.140 -86.330 ;
        RECT -131.100 -90.690 -129.900 -90.210 ;
        RECT -136.170 -92.260 -134.750 -91.850 ;
        RECT -135.840 -98.280 -135.070 -92.260 ;
        RECT -130.910 -98.280 -130.140 -90.690 ;
        RECT -125.930 -91.850 -125.160 -81.000 ;
        RECT -120.950 -85.920 -120.180 -81.000 ;
        RECT -121.290 -86.330 -119.870 -85.920 ;
        RECT -120.950 -90.210 -120.180 -86.330 ;
        RECT -121.180 -90.690 -119.980 -90.210 ;
        RECT -126.250 -92.260 -124.830 -91.850 ;
        RECT -125.930 -98.280 -125.160 -92.260 ;
        RECT -120.950 -98.280 -120.180 -90.690 ;
        RECT -116.030 -91.850 -115.260 -81.000 ;
        RECT -111.070 -85.920 -110.300 -81.000 ;
        RECT -111.370 -86.330 -109.950 -85.920 ;
        RECT -111.070 -90.210 -110.300 -86.330 ;
        RECT -111.260 -90.690 -110.060 -90.210 ;
        RECT -116.330 -92.260 -114.910 -91.850 ;
        RECT -116.030 -98.280 -115.260 -92.260 ;
        RECT -111.070 -98.280 -110.300 -90.690 ;
        RECT -106.100 -91.850 -105.330 -81.000 ;
        RECT -101.140 -85.920 -100.370 -81.000 ;
        RECT -101.450 -86.330 -100.030 -85.920 ;
        RECT -101.140 -90.210 -100.370 -86.330 ;
        RECT -101.340 -90.690 -100.140 -90.210 ;
        RECT -106.410 -92.260 -104.990 -91.850 ;
        RECT -106.100 -98.280 -105.330 -92.260 ;
        RECT -101.140 -98.280 -100.370 -90.690 ;
        RECT -96.150 -91.850 -95.380 -81.000 ;
        RECT -91.200 -85.920 -90.430 -81.000 ;
        RECT -91.530 -86.330 -90.110 -85.920 ;
        RECT -91.200 -90.210 -90.430 -86.330 ;
        RECT -91.420 -90.690 -90.220 -90.210 ;
        RECT -96.490 -92.260 -95.070 -91.850 ;
        RECT -96.150 -98.280 -95.380 -92.260 ;
        RECT -91.200 -98.280 -90.430 -90.690 ;
        RECT -86.250 -91.850 -85.480 -81.000 ;
        RECT -81.260 -85.920 -80.490 -81.000 ;
        RECT -81.610 -86.330 -80.190 -85.920 ;
        RECT -81.260 -90.210 -80.490 -86.330 ;
        RECT -81.500 -90.690 -80.300 -90.210 ;
        RECT -86.570 -92.260 -85.150 -91.850 ;
        RECT -86.250 -98.280 -85.480 -92.260 ;
        RECT -81.260 -98.280 -80.490 -90.690 ;
        RECT -76.340 -91.850 -75.570 -81.000 ;
        RECT -71.380 -85.920 -70.610 -81.000 ;
        RECT -71.690 -86.330 -70.270 -85.920 ;
        RECT -71.380 -90.210 -70.610 -86.330 ;
        RECT -71.580 -90.690 -70.380 -90.210 ;
        RECT -76.650 -92.260 -75.230 -91.850 ;
        RECT -76.340 -98.280 -75.570 -92.260 ;
        RECT -71.380 -98.280 -70.610 -90.690 ;
        RECT -66.400 -91.850 -65.630 -81.000 ;
        RECT -61.420 -85.920 -60.650 -81.000 ;
        RECT -61.770 -86.330 -60.350 -85.920 ;
        RECT -61.420 -90.210 -60.650 -86.330 ;
        RECT -61.660 -90.690 -60.460 -90.210 ;
        RECT -66.730 -92.260 -65.310 -91.850 ;
        RECT -66.400 -98.280 -65.630 -92.260 ;
        RECT -61.420 -98.280 -60.650 -90.690 ;
        RECT -56.510 -91.850 -55.740 -81.000 ;
        RECT -51.510 -85.920 -50.740 -81.000 ;
        RECT -51.850 -86.330 -50.430 -85.920 ;
        RECT -51.510 -90.210 -50.740 -86.330 ;
        RECT -51.740 -90.690 -50.540 -90.210 ;
        RECT -56.810 -92.260 -55.390 -91.850 ;
        RECT -56.510 -98.280 -55.740 -92.260 ;
        RECT -51.510 -98.280 -50.740 -90.690 ;
        RECT -46.550 -91.850 -45.780 -81.000 ;
        RECT -41.620 -85.920 -40.850 -81.000 ;
        RECT -41.930 -86.330 -40.510 -85.920 ;
        RECT -41.620 -90.210 -40.850 -86.330 ;
        RECT -41.820 -90.690 -40.620 -90.210 ;
        RECT -46.890 -92.260 -45.470 -91.850 ;
        RECT -46.550 -98.280 -45.780 -92.260 ;
        RECT -41.620 -98.280 -40.850 -90.690 ;
        RECT -36.670 -91.850 -35.900 -81.000 ;
        RECT -31.690 -85.920 -30.920 -81.000 ;
        RECT -32.010 -86.330 -30.590 -85.920 ;
        RECT -31.690 -90.210 -30.920 -86.330 ;
        RECT -31.900 -90.690 -30.700 -90.210 ;
        RECT -36.970 -92.260 -35.550 -91.850 ;
        RECT -36.670 -98.280 -35.900 -92.260 ;
        RECT -31.690 -98.280 -30.920 -90.690 ;
        RECT -26.740 -91.850 -25.970 -81.000 ;
        RECT -21.790 -85.920 -21.020 -81.000 ;
        RECT -22.090 -86.330 -20.670 -85.920 ;
        RECT -21.790 -90.210 -21.020 -86.330 ;
        RECT -21.980 -90.690 -20.780 -90.210 ;
        RECT -27.050 -92.260 -25.630 -91.850 ;
        RECT -26.740 -98.280 -25.970 -92.260 ;
        RECT -21.790 -98.280 -21.020 -90.690 ;
        RECT -16.810 -91.850 -16.040 -81.000 ;
        RECT -11.860 -85.920 -11.090 -81.000 ;
        RECT -12.170 -86.330 -10.750 -85.920 ;
        RECT -11.860 -90.210 -11.090 -86.330 ;
        RECT -12.060 -90.690 -10.860 -90.210 ;
        RECT -17.130 -92.260 -15.710 -91.850 ;
        RECT -16.810 -98.280 -16.040 -92.260 ;
        RECT -11.860 -98.280 -11.090 -90.690 ;
        RECT -6.910 -91.850 -6.140 -81.000 ;
        RECT -1.930 -85.920 -1.160 -81.000 ;
        RECT -2.250 -86.330 -0.830 -85.920 ;
        RECT -1.930 -90.210 -1.160 -86.330 ;
        RECT -2.140 -90.690 -0.940 -90.210 ;
        RECT -7.210 -92.260 -5.790 -91.850 ;
        RECT -6.910 -98.280 -6.140 -92.260 ;
        RECT -1.930 -98.280 -1.160 -90.690 ;
        RECT 3.020 -91.850 3.790 -81.000 ;
        RECT 7.950 -85.920 8.720 -81.000 ;
        RECT 7.670 -86.330 9.090 -85.920 ;
        RECT 7.950 -90.210 8.720 -86.330 ;
        RECT 7.780 -90.690 8.980 -90.210 ;
        RECT 2.710 -92.260 4.130 -91.850 ;
        RECT 3.020 -98.280 3.790 -92.260 ;
        RECT 7.950 -98.280 8.720 -90.690 ;
        RECT 12.950 -91.850 13.720 -81.000 ;
        RECT 17.900 -85.920 18.670 -81.000 ;
        RECT 17.590 -86.330 19.010 -85.920 ;
        RECT 17.900 -90.210 18.670 -86.330 ;
        RECT 17.700 -90.690 18.900 -90.210 ;
        RECT 12.630 -92.260 14.050 -91.850 ;
        RECT 12.950 -98.280 13.720 -92.260 ;
        RECT 17.900 -98.280 18.670 -90.690 ;
        RECT 22.880 -91.850 23.650 -81.000 ;
        RECT 27.890 -85.920 28.660 -81.000 ;
        RECT 27.510 -86.330 28.660 -85.920 ;
        RECT 27.890 -90.210 28.660 -86.330 ;
        RECT 27.620 -90.690 28.450 -90.210 ;
        RECT 22.550 -92.260 23.970 -91.850 ;
        RECT 22.880 -98.280 23.650 -92.260 ;
        RECT 27.890 -98.280 28.660 -90.690 ;
        RECT 31.340 -97.860 36.430 -81.000 ;
        RECT 138.320 -97.860 165.390 -14.140 ;
        RECT 29.710 -98.280 166.360 -97.860 ;
        RECT -296.740 -107.490 166.360 -98.280 ;
        RECT -296.740 -107.910 36.430 -107.490 ;
        RECT -296.740 -107.920 -291.650 -107.910 ;
        RECT -296.490 -159.080 -291.400 -158.900 ;
        RECT -29.520 -159.080 -0.060 -107.910 ;
        RECT 31.340 -108.040 36.430 -107.910 ;
        RECT 31.590 -159.080 36.680 -159.020 ;
        RECT -296.490 -168.710 36.680 -159.080 ;
        RECT -296.490 -185.990 -291.400 -168.710 ;
        RECT -289.360 -185.990 -288.590 -168.710 ;
        RECT -284.400 -179.560 -283.630 -168.710 ;
        RECT -279.440 -173.630 -278.670 -168.710 ;
        RECT -279.760 -174.040 -278.340 -173.630 ;
        RECT -279.440 -177.920 -278.670 -174.040 ;
        RECT -279.650 -178.400 -278.450 -177.920 ;
        RECT -284.720 -179.970 -283.300 -179.560 ;
        RECT -284.400 -185.990 -283.630 -179.970 ;
        RECT -279.440 -185.990 -278.670 -178.400 ;
        RECT -274.500 -179.560 -273.730 -168.710 ;
        RECT -269.520 -173.540 -268.750 -168.710 ;
        RECT -269.520 -173.630 -268.740 -173.540 ;
        RECT -269.840 -174.040 -268.420 -173.630 ;
        RECT -269.520 -175.990 -268.740 -174.040 ;
        RECT -269.560 -177.920 -268.740 -175.990 ;
        RECT -269.730 -178.400 -268.530 -177.920 ;
        RECT -274.800 -179.970 -273.380 -179.560 ;
        RECT -269.560 -179.890 -268.740 -178.400 ;
        RECT -264.550 -179.560 -263.780 -168.710 ;
        RECT -259.560 -173.630 -258.790 -168.710 ;
        RECT -259.920 -174.040 -258.500 -173.630 ;
        RECT -259.560 -177.920 -258.790 -174.040 ;
        RECT -259.810 -178.400 -258.610 -177.920 ;
        RECT -274.500 -185.990 -273.730 -179.970 ;
        RECT -269.570 -183.500 -268.740 -179.890 ;
        RECT -264.880 -179.970 -263.460 -179.560 ;
        RECT -269.570 -185.990 -268.750 -183.500 ;
        RECT -264.550 -185.990 -263.780 -179.970 ;
        RECT -259.560 -185.990 -258.790 -178.400 ;
        RECT -254.660 -179.560 -253.890 -168.710 ;
        RECT -249.670 -173.630 -248.900 -168.710 ;
        RECT -250.000 -174.040 -248.580 -173.630 ;
        RECT -249.670 -177.920 -248.900 -174.040 ;
        RECT -249.890 -178.400 -248.690 -177.920 ;
        RECT -254.960 -179.970 -253.540 -179.560 ;
        RECT -254.660 -185.990 -253.890 -179.970 ;
        RECT -249.670 -185.990 -248.900 -178.400 ;
        RECT -244.730 -179.560 -243.960 -168.710 ;
        RECT -239.760 -173.630 -238.990 -168.710 ;
        RECT -240.080 -174.040 -238.660 -173.630 ;
        RECT -239.760 -177.920 -238.990 -174.040 ;
        RECT -239.970 -178.400 -238.770 -177.920 ;
        RECT -245.040 -179.970 -243.620 -179.560 ;
        RECT -244.730 -185.990 -243.960 -179.970 ;
        RECT -239.760 -185.990 -238.990 -178.400 ;
        RECT -234.820 -179.560 -234.050 -168.710 ;
        RECT -229.860 -173.630 -229.090 -168.710 ;
        RECT -230.160 -174.040 -228.740 -173.630 ;
        RECT -229.860 -177.920 -229.090 -174.040 ;
        RECT -230.050 -178.400 -228.850 -177.920 ;
        RECT -235.120 -179.970 -233.700 -179.560 ;
        RECT -234.820 -185.990 -234.050 -179.970 ;
        RECT -229.860 -185.990 -229.090 -178.400 ;
        RECT -224.890 -179.560 -224.120 -168.710 ;
        RECT -219.920 -173.630 -219.150 -168.710 ;
        RECT -220.240 -174.040 -218.820 -173.630 ;
        RECT -219.920 -177.920 -219.150 -174.040 ;
        RECT -220.130 -178.400 -218.930 -177.920 ;
        RECT -225.200 -179.970 -223.780 -179.560 ;
        RECT -224.890 -185.990 -224.120 -179.970 ;
        RECT -219.920 -185.990 -219.150 -178.400 ;
        RECT -214.940 -179.560 -214.170 -168.710 ;
        RECT -209.980 -173.630 -209.210 -168.710 ;
        RECT -210.320 -174.040 -208.900 -173.630 ;
        RECT -209.980 -177.920 -209.210 -174.040 ;
        RECT -210.210 -178.400 -209.010 -177.920 ;
        RECT -215.280 -179.970 -213.860 -179.560 ;
        RECT -214.940 -185.990 -214.170 -179.970 ;
        RECT -209.980 -185.990 -209.210 -178.400 ;
        RECT -205.030 -179.560 -204.260 -168.710 ;
        RECT -200.090 -173.630 -199.320 -168.710 ;
        RECT -200.400 -174.040 -198.980 -173.630 ;
        RECT -200.090 -177.920 -199.320 -174.040 ;
        RECT -200.290 -178.400 -199.090 -177.920 ;
        RECT -205.360 -179.970 -203.940 -179.560 ;
        RECT -205.030 -185.990 -204.260 -179.970 ;
        RECT -200.090 -185.990 -199.320 -178.400 ;
        RECT -195.160 -179.560 -194.390 -168.710 ;
        RECT -190.160 -173.630 -189.390 -168.710 ;
        RECT -190.480 -174.040 -189.060 -173.630 ;
        RECT -190.160 -177.920 -189.390 -174.040 ;
        RECT -190.370 -178.400 -189.170 -177.920 ;
        RECT -195.440 -179.970 -194.020 -179.560 ;
        RECT -195.160 -185.990 -194.390 -179.970 ;
        RECT -190.160 -185.990 -189.390 -178.400 ;
        RECT -185.200 -179.560 -184.430 -168.710 ;
        RECT -180.250 -173.630 -179.480 -168.710 ;
        RECT -180.560 -174.040 -179.140 -173.630 ;
        RECT -180.250 -177.920 -179.480 -174.040 ;
        RECT -180.450 -178.400 -179.250 -177.920 ;
        RECT -185.520 -179.970 -184.100 -179.560 ;
        RECT -185.200 -185.990 -184.430 -179.970 ;
        RECT -180.250 -185.990 -179.480 -178.400 ;
        RECT -175.290 -179.560 -174.520 -168.710 ;
        RECT -170.300 -173.630 -169.530 -168.710 ;
        RECT -170.640 -174.040 -169.220 -173.630 ;
        RECT -170.300 -177.920 -169.530 -174.040 ;
        RECT -170.530 -178.400 -169.330 -177.920 ;
        RECT -175.600 -179.970 -174.180 -179.560 ;
        RECT -175.290 -185.990 -174.520 -179.970 ;
        RECT -170.300 -185.990 -169.530 -178.400 ;
        RECT -165.360 -179.560 -164.590 -168.710 ;
        RECT -160.360 -173.630 -159.590 -168.710 ;
        RECT -160.720 -174.040 -159.300 -173.630 ;
        RECT -160.360 -177.920 -159.590 -174.040 ;
        RECT -160.610 -178.400 -159.410 -177.920 ;
        RECT -165.680 -179.970 -164.260 -179.560 ;
        RECT -165.360 -185.990 -164.590 -179.970 ;
        RECT -160.360 -185.990 -159.590 -178.400 ;
        RECT -155.450 -179.560 -154.680 -168.710 ;
        RECT -150.500 -173.630 -149.730 -168.710 ;
        RECT -150.800 -174.040 -149.380 -173.630 ;
        RECT -150.500 -177.920 -149.730 -174.040 ;
        RECT -150.690 -178.400 -149.490 -177.920 ;
        RECT -155.760 -179.970 -154.340 -179.560 ;
        RECT -155.450 -185.990 -154.680 -179.970 ;
        RECT -150.500 -185.990 -149.730 -178.400 ;
        RECT -145.530 -179.560 -144.760 -168.710 ;
        RECT -140.570 -173.630 -139.800 -168.710 ;
        RECT -140.880 -174.040 -139.460 -173.630 ;
        RECT -140.570 -177.920 -139.800 -174.040 ;
        RECT -140.770 -178.400 -139.570 -177.920 ;
        RECT -145.840 -179.970 -144.420 -179.560 ;
        RECT -145.530 -185.990 -144.760 -179.970 ;
        RECT -140.570 -185.990 -139.800 -178.400 ;
        RECT -135.590 -179.560 -134.820 -168.710 ;
        RECT -130.660 -173.630 -129.890 -168.710 ;
        RECT -130.960 -174.040 -129.540 -173.630 ;
        RECT -130.660 -177.920 -129.890 -174.040 ;
        RECT -130.850 -178.400 -129.650 -177.920 ;
        RECT -135.920 -179.970 -134.500 -179.560 ;
        RECT -135.590 -185.990 -134.820 -179.970 ;
        RECT -130.660 -185.990 -129.890 -178.400 ;
        RECT -125.680 -179.560 -124.910 -168.710 ;
        RECT -120.700 -173.630 -119.930 -168.710 ;
        RECT -121.040 -174.040 -119.620 -173.630 ;
        RECT -120.700 -177.920 -119.930 -174.040 ;
        RECT -120.930 -178.400 -119.730 -177.920 ;
        RECT -126.000 -179.970 -124.580 -179.560 ;
        RECT -125.680 -185.990 -124.910 -179.970 ;
        RECT -120.700 -185.990 -119.930 -178.400 ;
        RECT -115.780 -179.560 -115.010 -168.710 ;
        RECT -110.820 -173.630 -110.050 -168.710 ;
        RECT -111.120 -174.040 -109.700 -173.630 ;
        RECT -110.820 -177.920 -110.050 -174.040 ;
        RECT -111.010 -178.400 -109.810 -177.920 ;
        RECT -116.080 -179.970 -114.660 -179.560 ;
        RECT -115.780 -185.990 -115.010 -179.970 ;
        RECT -110.820 -185.990 -110.050 -178.400 ;
        RECT -105.850 -179.560 -105.080 -168.710 ;
        RECT -100.890 -173.630 -100.120 -168.710 ;
        RECT -101.200 -174.040 -99.780 -173.630 ;
        RECT -100.890 -177.920 -100.120 -174.040 ;
        RECT -101.090 -178.400 -99.890 -177.920 ;
        RECT -106.160 -179.970 -104.740 -179.560 ;
        RECT -105.850 -185.990 -105.080 -179.970 ;
        RECT -100.890 -185.990 -100.120 -178.400 ;
        RECT -95.900 -179.560 -95.130 -168.710 ;
        RECT -90.950 -173.630 -90.180 -168.710 ;
        RECT -91.280 -174.040 -89.860 -173.630 ;
        RECT -90.950 -177.920 -90.180 -174.040 ;
        RECT -91.170 -178.400 -89.970 -177.920 ;
        RECT -96.240 -179.970 -94.820 -179.560 ;
        RECT -95.900 -185.990 -95.130 -179.970 ;
        RECT -90.950 -185.990 -90.180 -178.400 ;
        RECT -86.000 -179.560 -85.230 -168.710 ;
        RECT -81.010 -173.630 -80.240 -168.710 ;
        RECT -81.360 -174.040 -79.940 -173.630 ;
        RECT -81.010 -177.920 -80.240 -174.040 ;
        RECT -81.250 -178.400 -80.050 -177.920 ;
        RECT -86.320 -179.970 -84.900 -179.560 ;
        RECT -86.000 -185.990 -85.230 -179.970 ;
        RECT -81.010 -185.990 -80.240 -178.400 ;
        RECT -76.090 -179.560 -75.320 -168.710 ;
        RECT -71.130 -173.630 -70.360 -168.710 ;
        RECT -71.440 -174.040 -70.020 -173.630 ;
        RECT -71.130 -177.920 -70.360 -174.040 ;
        RECT -71.330 -178.400 -70.130 -177.920 ;
        RECT -76.400 -179.970 -74.980 -179.560 ;
        RECT -76.090 -185.990 -75.320 -179.970 ;
        RECT -71.130 -185.990 -70.360 -178.400 ;
        RECT -66.150 -179.560 -65.380 -168.710 ;
        RECT -61.170 -173.630 -60.400 -168.710 ;
        RECT -61.520 -174.040 -60.100 -173.630 ;
        RECT -61.170 -177.920 -60.400 -174.040 ;
        RECT -61.410 -178.400 -60.210 -177.920 ;
        RECT -66.480 -179.970 -65.060 -179.560 ;
        RECT -66.150 -185.990 -65.380 -179.970 ;
        RECT -61.170 -185.990 -60.400 -178.400 ;
        RECT -56.260 -179.560 -55.490 -168.710 ;
        RECT -51.260 -173.630 -50.490 -168.710 ;
        RECT -51.600 -174.040 -50.180 -173.630 ;
        RECT -51.260 -177.920 -50.490 -174.040 ;
        RECT -51.490 -178.400 -50.290 -177.920 ;
        RECT -56.560 -179.970 -55.140 -179.560 ;
        RECT -56.260 -185.990 -55.490 -179.970 ;
        RECT -51.260 -185.990 -50.490 -178.400 ;
        RECT -46.300 -179.560 -45.530 -168.710 ;
        RECT -41.370 -173.630 -40.600 -168.710 ;
        RECT -41.680 -174.040 -40.260 -173.630 ;
        RECT -41.370 -177.920 -40.600 -174.040 ;
        RECT -41.570 -178.400 -40.370 -177.920 ;
        RECT -46.640 -179.970 -45.220 -179.560 ;
        RECT -46.300 -185.990 -45.530 -179.970 ;
        RECT -41.370 -185.990 -40.600 -178.400 ;
        RECT -36.420 -179.560 -35.650 -168.710 ;
        RECT -31.440 -173.630 -30.670 -168.710 ;
        RECT -31.760 -174.040 -30.340 -173.630 ;
        RECT -31.440 -177.920 -30.670 -174.040 ;
        RECT -31.650 -178.400 -30.450 -177.920 ;
        RECT -36.720 -179.970 -35.300 -179.560 ;
        RECT -36.420 -185.990 -35.650 -179.970 ;
        RECT -31.440 -185.990 -30.670 -178.400 ;
        RECT -26.490 -179.560 -25.720 -168.710 ;
        RECT -21.540 -173.630 -20.770 -168.710 ;
        RECT -21.840 -174.040 -20.420 -173.630 ;
        RECT -21.540 -177.920 -20.770 -174.040 ;
        RECT -21.730 -178.400 -20.530 -177.920 ;
        RECT -26.800 -179.970 -25.380 -179.560 ;
        RECT -26.490 -185.990 -25.720 -179.970 ;
        RECT -21.540 -185.990 -20.770 -178.400 ;
        RECT -16.560 -179.560 -15.790 -168.710 ;
        RECT -11.610 -173.630 -10.840 -168.710 ;
        RECT -11.920 -174.040 -10.500 -173.630 ;
        RECT -11.610 -177.920 -10.840 -174.040 ;
        RECT -11.810 -178.400 -10.610 -177.920 ;
        RECT -16.880 -179.970 -15.460 -179.560 ;
        RECT -16.560 -185.990 -15.790 -179.970 ;
        RECT -11.610 -185.990 -10.840 -178.400 ;
        RECT -6.660 -179.560 -5.890 -168.710 ;
        RECT -1.680 -173.630 -0.910 -168.710 ;
        RECT -2.000 -174.040 -0.580 -173.630 ;
        RECT -1.680 -177.920 -0.910 -174.040 ;
        RECT -1.890 -178.400 -0.690 -177.920 ;
        RECT -6.960 -179.970 -5.540 -179.560 ;
        RECT -6.660 -185.990 -5.890 -179.970 ;
        RECT -1.680 -185.990 -0.910 -178.400 ;
        RECT 3.270 -179.560 4.040 -168.710 ;
        RECT 8.200 -173.630 8.970 -168.710 ;
        RECT 7.920 -174.040 9.340 -173.630 ;
        RECT 8.200 -177.920 8.970 -174.040 ;
        RECT 8.030 -178.400 9.230 -177.920 ;
        RECT 2.960 -179.970 4.380 -179.560 ;
        RECT 3.270 -185.990 4.040 -179.970 ;
        RECT 8.200 -185.990 8.970 -178.400 ;
        RECT 13.200 -179.560 13.970 -168.710 ;
        RECT 18.150 -173.630 18.920 -168.710 ;
        RECT 17.840 -174.040 19.260 -173.630 ;
        RECT 18.150 -177.920 18.920 -174.040 ;
        RECT 17.950 -178.400 19.150 -177.920 ;
        RECT 12.880 -179.970 14.300 -179.560 ;
        RECT 13.200 -185.990 13.970 -179.970 ;
        RECT 18.150 -185.990 18.920 -178.400 ;
        RECT 23.130 -179.560 23.900 -168.710 ;
        RECT 28.140 -173.630 28.910 -168.710 ;
        RECT 27.760 -174.040 28.910 -173.630 ;
        RECT 28.140 -177.920 28.910 -174.040 ;
        RECT 27.870 -178.400 28.700 -177.920 ;
        RECT 22.800 -179.970 24.220 -179.560 ;
        RECT 23.130 -185.990 23.900 -179.970 ;
        RECT 28.140 -185.990 28.910 -178.400 ;
        RECT 31.590 -185.570 36.680 -168.710 ;
        RECT 138.320 -185.570 165.390 -107.490 ;
        RECT 29.960 -185.990 166.610 -185.570 ;
        RECT -296.490 -195.200 166.610 -185.990 ;
        RECT -296.490 -195.620 36.680 -195.200 ;
        RECT -296.490 -195.630 -291.400 -195.620 ;
        RECT 31.590 -195.750 36.680 -195.620 ;
        RECT 138.320 -196.620 165.390 -195.200 ;
      LAYER via3 ;
        RECT -237.115 43.280 -226.395 52.800 ;
        RECT 144.705 42.570 155.425 52.090 ;
        RECT -168.635 -44.930 -157.915 -35.410 ;
        RECT 147.055 -52.660 157.775 -43.140 ;
        RECT -20.075 -134.680 -9.355 -125.160 ;
        RECT 144.735 -144.350 155.455 -134.830 ;
      LAYER met4 ;
        RECT -240.990 40.070 -223.200 58.260 ;
        RECT 140.870 39.000 159.450 56.810 ;
        RECT -172.120 -49.690 -153.930 -30.730 ;
        RECT 142.790 -56.650 161.470 -39.040 ;
        RECT -23.180 -139.440 -5.770 -120.480 ;
        RECT 141.240 -149.110 159.920 -131.500 ;
    END
  END VPWR
  PIN o_ranQ[60]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -274.325 94.875 -272.115 95.055 ;
        RECT -274.325 94.795 -273.820 94.875 ;
        RECT -273.020 94.785 -272.115 94.875 ;
      LAYER mcon ;
        RECT -274.135 94.795 -273.965 94.965 ;
        RECT -272.770 94.795 -272.600 94.965 ;
      LAYER met1 ;
        RECT -274.020 95.060 -273.020 95.760 ;
        RECT -274.200 94.760 -272.510 95.060 ;
    END
  END o_ranQ[60]
  PIN o_ranQ[124]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -274.075 7.165 -271.865 7.345 ;
        RECT -274.075 7.085 -273.570 7.165 ;
        RECT -272.770 7.075 -271.865 7.165 ;
      LAYER mcon ;
        RECT -273.885 7.085 -273.715 7.255 ;
        RECT -272.520 7.085 -272.350 7.255 ;
      LAYER met1 ;
        RECT -273.770 7.350 -272.770 8.050 ;
        RECT -273.950 7.050 -272.260 7.350 ;
    END
  END o_ranQ[124]
  PIN o_ranQ[65]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 18.565 1.355 19.070 1.435 ;
        RECT 19.870 1.355 20.775 1.445 ;
        RECT 18.565 1.175 20.775 1.355 ;
      LAYER mcon ;
        RECT 18.755 1.265 18.925 1.435 ;
        RECT 20.120 1.265 20.290 1.435 ;
      LAYER met1 ;
        RECT 18.690 1.170 20.380 1.470 ;
        RECT 18.870 0.470 19.870 1.170 ;
    END
  END o_ranQ[65]
  PIN o_ranQ[66]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 13.605 7.165 15.815 7.345 ;
        RECT 13.605 7.085 14.110 7.165 ;
        RECT 14.910 7.075 15.815 7.165 ;
      LAYER mcon ;
        RECT 13.795 7.085 13.965 7.255 ;
        RECT 15.160 7.085 15.330 7.255 ;
      LAYER met1 ;
        RECT 13.910 7.350 14.910 8.050 ;
        RECT 13.730 7.050 15.420 7.350 ;
    END
  END o_ranQ[66]
  PIN o_ranQ[67]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 8.645 1.355 9.150 1.435 ;
        RECT 9.950 1.355 10.855 1.445 ;
        RECT 8.645 1.175 10.855 1.355 ;
      LAYER mcon ;
        RECT 8.835 1.265 9.005 1.435 ;
        RECT 10.200 1.265 10.370 1.435 ;
      LAYER met1 ;
        RECT 8.770 1.170 10.460 1.470 ;
        RECT 8.950 0.470 9.950 1.170 ;
    END
  END o_ranQ[67]
  PIN o_ranQ[64]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 23.525 7.165 25.735 7.345 ;
        RECT 23.525 7.085 24.030 7.165 ;
        RECT 24.830 7.075 25.735 7.165 ;
      LAYER mcon ;
        RECT 23.715 7.085 23.885 7.255 ;
        RECT 25.080 7.085 25.250 7.255 ;
      LAYER met1 ;
        RECT 23.830 7.350 24.830 8.050 ;
        RECT 23.650 7.050 25.340 7.350 ;
    END
  END o_ranQ[64]
  PIN o_ranQ[68]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 3.685 7.165 5.895 7.345 ;
        RECT 3.685 7.085 4.190 7.165 ;
        RECT 4.990 7.075 5.895 7.165 ;
      LAYER mcon ;
        RECT 3.875 7.085 4.045 7.255 ;
        RECT 5.240 7.085 5.410 7.255 ;
      LAYER met1 ;
        RECT 3.990 7.350 4.990 8.050 ;
        RECT 3.810 7.050 5.500 7.350 ;
    END
  END o_ranQ[68]
  PIN o_ranQ[69]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -1.275 1.355 -0.770 1.435 ;
        RECT 0.030 1.355 0.935 1.445 ;
        RECT -1.275 1.175 0.935 1.355 ;
      LAYER mcon ;
        RECT -1.085 1.265 -0.915 1.435 ;
        RECT 0.280 1.265 0.450 1.435 ;
      LAYER met1 ;
        RECT -1.150 1.170 0.540 1.470 ;
        RECT -0.970 0.470 0.030 1.170 ;
    END
  END o_ranQ[69]
  PIN o_ranQ[70]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -6.235 7.165 -4.025 7.345 ;
        RECT -6.235 7.085 -5.730 7.165 ;
        RECT -4.930 7.075 -4.025 7.165 ;
      LAYER mcon ;
        RECT -6.045 7.085 -5.875 7.255 ;
        RECT -4.680 7.085 -4.510 7.255 ;
      LAYER met1 ;
        RECT -5.930 7.350 -4.930 8.050 ;
        RECT -6.110 7.050 -4.420 7.350 ;
    END
  END o_ranQ[70]
  PIN o_ranQ[71]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -11.195 1.355 -10.690 1.435 ;
        RECT -9.890 1.355 -8.985 1.445 ;
        RECT -11.195 1.175 -8.985 1.355 ;
      LAYER mcon ;
        RECT -11.005 1.265 -10.835 1.435 ;
        RECT -9.640 1.265 -9.470 1.435 ;
      LAYER met1 ;
        RECT -11.070 1.170 -9.380 1.470 ;
        RECT -10.890 0.470 -9.890 1.170 ;
    END
  END o_ranQ[71]
  PIN o_ranQ[72]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -16.155 7.165 -13.945 7.345 ;
        RECT -16.155 7.085 -15.650 7.165 ;
        RECT -14.850 7.075 -13.945 7.165 ;
      LAYER mcon ;
        RECT -15.965 7.085 -15.795 7.255 ;
        RECT -14.600 7.085 -14.430 7.255 ;
      LAYER met1 ;
        RECT -15.850 7.350 -14.850 8.050 ;
        RECT -16.030 7.050 -14.340 7.350 ;
    END
  END o_ranQ[72]
  PIN o_ranQ[73]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -21.115 1.355 -20.610 1.435 ;
        RECT -19.810 1.355 -18.905 1.445 ;
        RECT -21.115 1.175 -18.905 1.355 ;
      LAYER mcon ;
        RECT -20.925 1.265 -20.755 1.435 ;
        RECT -19.560 1.265 -19.390 1.435 ;
      LAYER met1 ;
        RECT -20.990 1.170 -19.300 1.470 ;
        RECT -20.810 0.470 -19.810 1.170 ;
    END
  END o_ranQ[73]
  PIN o_ranQ[74]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -26.075 7.165 -23.865 7.345 ;
        RECT -26.075 7.085 -25.570 7.165 ;
        RECT -24.770 7.075 -23.865 7.165 ;
      LAYER mcon ;
        RECT -25.885 7.085 -25.715 7.255 ;
        RECT -24.520 7.085 -24.350 7.255 ;
      LAYER met1 ;
        RECT -25.770 7.350 -24.770 8.050 ;
        RECT -25.950 7.050 -24.260 7.350 ;
    END
  END o_ranQ[74]
  PIN o_ranQ[75]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -31.035 1.355 -30.530 1.435 ;
        RECT -29.730 1.355 -28.825 1.445 ;
        RECT -31.035 1.175 -28.825 1.355 ;
      LAYER mcon ;
        RECT -30.845 1.265 -30.675 1.435 ;
        RECT -29.480 1.265 -29.310 1.435 ;
      LAYER met1 ;
        RECT -30.910 1.170 -29.220 1.470 ;
        RECT -30.730 0.470 -29.730 1.170 ;
    END
  END o_ranQ[75]
  PIN o_ranQ[76]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -35.995 7.165 -33.785 7.345 ;
        RECT -35.995 7.085 -35.490 7.165 ;
        RECT -34.690 7.075 -33.785 7.165 ;
      LAYER mcon ;
        RECT -35.805 7.085 -35.635 7.255 ;
        RECT -34.440 7.085 -34.270 7.255 ;
      LAYER met1 ;
        RECT -35.690 7.350 -34.690 8.050 ;
        RECT -35.870 7.050 -34.180 7.350 ;
    END
  END o_ranQ[76]
  PIN o_ranQ[77]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -40.955 1.355 -40.450 1.435 ;
        RECT -39.650 1.355 -38.745 1.445 ;
        RECT -40.955 1.175 -38.745 1.355 ;
      LAYER mcon ;
        RECT -40.765 1.265 -40.595 1.435 ;
        RECT -39.400 1.265 -39.230 1.435 ;
      LAYER met1 ;
        RECT -40.830 1.170 -39.140 1.470 ;
        RECT -40.650 0.470 -39.650 1.170 ;
    END
  END o_ranQ[77]
  PIN o_ranQ[78]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -45.915 7.165 -43.705 7.345 ;
        RECT -45.915 7.085 -45.410 7.165 ;
        RECT -44.610 7.075 -43.705 7.165 ;
      LAYER mcon ;
        RECT -45.725 7.085 -45.555 7.255 ;
        RECT -44.360 7.085 -44.190 7.255 ;
      LAYER met1 ;
        RECT -45.610 7.350 -44.610 8.050 ;
        RECT -45.790 7.050 -44.100 7.350 ;
    END
  END o_ranQ[78]
  PIN o_ranQ[79]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -50.875 1.355 -50.370 1.435 ;
        RECT -49.570 1.355 -48.665 1.445 ;
        RECT -50.875 1.175 -48.665 1.355 ;
      LAYER mcon ;
        RECT -50.685 1.265 -50.515 1.435 ;
        RECT -49.320 1.265 -49.150 1.435 ;
      LAYER met1 ;
        RECT -50.750 1.170 -49.060 1.470 ;
        RECT -50.570 0.470 -49.570 1.170 ;
    END
  END o_ranQ[79]
  PIN o_ranQ[81]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -60.795 1.355 -60.290 1.435 ;
        RECT -59.490 1.355 -58.585 1.445 ;
        RECT -60.795 1.175 -58.585 1.355 ;
      LAYER mcon ;
        RECT -60.605 1.265 -60.435 1.435 ;
        RECT -59.240 1.265 -59.070 1.435 ;
      LAYER met1 ;
        RECT -60.670 1.170 -58.980 1.470 ;
        RECT -60.490 0.470 -59.490 1.170 ;
    END
  END o_ranQ[81]
  PIN o_ranQ[82]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -65.755 7.165 -63.545 7.345 ;
        RECT -65.755 7.085 -65.250 7.165 ;
        RECT -64.450 7.075 -63.545 7.165 ;
      LAYER mcon ;
        RECT -65.565 7.085 -65.395 7.255 ;
        RECT -64.200 7.085 -64.030 7.255 ;
      LAYER met1 ;
        RECT -65.450 7.350 -64.450 8.050 ;
        RECT -65.630 7.050 -63.940 7.350 ;
    END
  END o_ranQ[82]
  PIN o_ranQ[83]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -70.715 1.355 -70.210 1.435 ;
        RECT -69.410 1.355 -68.505 1.445 ;
        RECT -70.715 1.175 -68.505 1.355 ;
      LAYER mcon ;
        RECT -70.525 1.265 -70.355 1.435 ;
        RECT -69.160 1.265 -68.990 1.435 ;
      LAYER met1 ;
        RECT -70.590 1.170 -68.900 1.470 ;
        RECT -70.410 0.470 -69.410 1.170 ;
    END
  END o_ranQ[83]
  PIN o_ranQ[80]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -55.835 7.165 -53.625 7.345 ;
        RECT -55.835 7.085 -55.330 7.165 ;
        RECT -54.530 7.075 -53.625 7.165 ;
      LAYER mcon ;
        RECT -55.645 7.085 -55.475 7.255 ;
        RECT -54.280 7.085 -54.110 7.255 ;
      LAYER met1 ;
        RECT -55.530 7.350 -54.530 8.050 ;
        RECT -55.710 7.050 -54.020 7.350 ;
    END
  END o_ranQ[80]
  PIN o_ranQ[84]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -75.675 7.165 -73.465 7.345 ;
        RECT -75.675 7.085 -75.170 7.165 ;
        RECT -74.370 7.075 -73.465 7.165 ;
      LAYER mcon ;
        RECT -75.485 7.085 -75.315 7.255 ;
        RECT -74.120 7.085 -73.950 7.255 ;
      LAYER met1 ;
        RECT -75.370 7.350 -74.370 8.050 ;
        RECT -75.550 7.050 -73.860 7.350 ;
    END
  END o_ranQ[84]
  PIN o_ranQ[85]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -80.635 1.355 -80.130 1.435 ;
        RECT -79.330 1.355 -78.425 1.445 ;
        RECT -80.635 1.175 -78.425 1.355 ;
      LAYER mcon ;
        RECT -80.445 1.265 -80.275 1.435 ;
        RECT -79.080 1.265 -78.910 1.435 ;
      LAYER met1 ;
        RECT -80.510 1.170 -78.820 1.470 ;
        RECT -80.330 0.470 -79.330 1.170 ;
    END
  END o_ranQ[85]
  PIN o_ranQ[86]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -85.595 7.165 -83.385 7.345 ;
        RECT -85.595 7.085 -85.090 7.165 ;
        RECT -84.290 7.075 -83.385 7.165 ;
      LAYER mcon ;
        RECT -85.405 7.085 -85.235 7.255 ;
        RECT -84.040 7.085 -83.870 7.255 ;
      LAYER met1 ;
        RECT -85.290 7.350 -84.290 8.050 ;
        RECT -85.470 7.050 -83.780 7.350 ;
    END
  END o_ranQ[86]
  PIN o_ranQ[87]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -90.555 1.355 -90.050 1.435 ;
        RECT -89.250 1.355 -88.345 1.445 ;
        RECT -90.555 1.175 -88.345 1.355 ;
      LAYER mcon ;
        RECT -90.365 1.265 -90.195 1.435 ;
        RECT -89.000 1.265 -88.830 1.435 ;
      LAYER met1 ;
        RECT -90.430 1.170 -88.740 1.470 ;
        RECT -90.250 0.470 -89.250 1.170 ;
    END
  END o_ranQ[87]
  PIN o_ranQ[88]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -95.515 7.165 -93.305 7.345 ;
        RECT -95.515 7.085 -95.010 7.165 ;
        RECT -94.210 7.075 -93.305 7.165 ;
      LAYER mcon ;
        RECT -95.325 7.085 -95.155 7.255 ;
        RECT -93.960 7.085 -93.790 7.255 ;
      LAYER met1 ;
        RECT -95.210 7.350 -94.210 8.050 ;
        RECT -95.390 7.050 -93.700 7.350 ;
    END
  END o_ranQ[88]
  PIN o_ranQ[89]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -100.475 1.355 -99.970 1.435 ;
        RECT -99.170 1.355 -98.265 1.445 ;
        RECT -100.475 1.175 -98.265 1.355 ;
      LAYER mcon ;
        RECT -100.285 1.265 -100.115 1.435 ;
        RECT -98.920 1.265 -98.750 1.435 ;
      LAYER met1 ;
        RECT -100.350 1.170 -98.660 1.470 ;
        RECT -100.170 0.470 -99.170 1.170 ;
    END
  END o_ranQ[89]
  PIN o_ranQ[90]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -105.435 7.165 -103.225 7.345 ;
        RECT -105.435 7.085 -104.930 7.165 ;
        RECT -104.130 7.075 -103.225 7.165 ;
      LAYER mcon ;
        RECT -105.245 7.085 -105.075 7.255 ;
        RECT -103.880 7.085 -103.710 7.255 ;
      LAYER met1 ;
        RECT -105.130 7.350 -104.130 8.050 ;
        RECT -105.310 7.050 -103.620 7.350 ;
    END
  END o_ranQ[90]
  PIN o_ranQ[91]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -110.395 1.355 -109.890 1.435 ;
        RECT -109.090 1.355 -108.185 1.445 ;
        RECT -110.395 1.175 -108.185 1.355 ;
      LAYER mcon ;
        RECT -110.205 1.265 -110.035 1.435 ;
        RECT -108.840 1.265 -108.670 1.435 ;
      LAYER met1 ;
        RECT -110.270 1.170 -108.580 1.470 ;
        RECT -110.090 0.470 -109.090 1.170 ;
    END
  END o_ranQ[91]
  PIN o_ranQ[92]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -115.355 7.165 -113.145 7.345 ;
        RECT -115.355 7.085 -114.850 7.165 ;
        RECT -114.050 7.075 -113.145 7.165 ;
      LAYER mcon ;
        RECT -115.165 7.085 -114.995 7.255 ;
        RECT -113.800 7.085 -113.630 7.255 ;
      LAYER met1 ;
        RECT -115.050 7.350 -114.050 8.050 ;
        RECT -115.230 7.050 -113.540 7.350 ;
    END
  END o_ranQ[92]
  PIN o_ranQ[93]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -120.315 1.355 -119.810 1.435 ;
        RECT -119.010 1.355 -118.105 1.445 ;
        RECT -120.315 1.175 -118.105 1.355 ;
      LAYER mcon ;
        RECT -120.125 1.265 -119.955 1.435 ;
        RECT -118.760 1.265 -118.590 1.435 ;
      LAYER met1 ;
        RECT -120.190 1.170 -118.500 1.470 ;
        RECT -120.010 0.470 -119.010 1.170 ;
    END
  END o_ranQ[93]
  PIN o_ranQ[94]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -125.275 7.165 -123.065 7.345 ;
        RECT -125.275 7.085 -124.770 7.165 ;
        RECT -123.970 7.075 -123.065 7.165 ;
      LAYER mcon ;
        RECT -125.085 7.085 -124.915 7.255 ;
        RECT -123.720 7.085 -123.550 7.255 ;
      LAYER met1 ;
        RECT -124.970 7.350 -123.970 8.050 ;
        RECT -125.150 7.050 -123.460 7.350 ;
    END
  END o_ranQ[94]
  PIN o_ranQ[95]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -130.235 1.355 -129.730 1.435 ;
        RECT -128.930 1.355 -128.025 1.445 ;
        RECT -130.235 1.175 -128.025 1.355 ;
      LAYER mcon ;
        RECT -130.045 1.265 -129.875 1.435 ;
        RECT -128.680 1.265 -128.510 1.435 ;
      LAYER met1 ;
        RECT -130.110 1.170 -128.420 1.470 ;
        RECT -129.930 0.470 -128.930 1.170 ;
    END
  END o_ranQ[95]
  PIN o_ranQ[97]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -140.155 1.355 -139.650 1.435 ;
        RECT -138.850 1.355 -137.945 1.445 ;
        RECT -140.155 1.175 -137.945 1.355 ;
      LAYER mcon ;
        RECT -139.965 1.265 -139.795 1.435 ;
        RECT -138.600 1.265 -138.430 1.435 ;
      LAYER met1 ;
        RECT -140.030 1.170 -138.340 1.470 ;
        RECT -139.850 0.470 -138.850 1.170 ;
    END
  END o_ranQ[97]
  PIN o_ranQ[98]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -145.115 7.165 -142.905 7.345 ;
        RECT -145.115 7.085 -144.610 7.165 ;
        RECT -143.810 7.075 -142.905 7.165 ;
      LAYER mcon ;
        RECT -144.925 7.085 -144.755 7.255 ;
        RECT -143.560 7.085 -143.390 7.255 ;
      LAYER met1 ;
        RECT -144.810 7.350 -143.810 8.050 ;
        RECT -144.990 7.050 -143.300 7.350 ;
    END
  END o_ranQ[98]
  PIN o_ranQ[99]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -150.075 1.355 -149.570 1.435 ;
        RECT -148.770 1.355 -147.865 1.445 ;
        RECT -150.075 1.175 -147.865 1.355 ;
      LAYER mcon ;
        RECT -149.885 1.265 -149.715 1.435 ;
        RECT -148.520 1.265 -148.350 1.435 ;
      LAYER met1 ;
        RECT -149.950 1.170 -148.260 1.470 ;
        RECT -149.770 0.470 -148.770 1.170 ;
    END
  END o_ranQ[99]
  PIN o_ranQ[96]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -135.195 7.165 -132.985 7.345 ;
        RECT -135.195 7.085 -134.690 7.165 ;
        RECT -133.890 7.075 -132.985 7.165 ;
      LAYER mcon ;
        RECT -135.005 7.085 -134.835 7.255 ;
        RECT -133.640 7.085 -133.470 7.255 ;
      LAYER met1 ;
        RECT -134.890 7.350 -133.890 8.050 ;
        RECT -135.070 7.050 -133.380 7.350 ;
    END
  END o_ranQ[96]
  PIN o_ranQ[100]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -155.035 7.165 -152.825 7.345 ;
        RECT -155.035 7.085 -154.530 7.165 ;
        RECT -153.730 7.075 -152.825 7.165 ;
      LAYER mcon ;
        RECT -154.845 7.085 -154.675 7.255 ;
        RECT -153.480 7.085 -153.310 7.255 ;
      LAYER met1 ;
        RECT -154.730 7.350 -153.730 8.050 ;
        RECT -154.910 7.050 -153.220 7.350 ;
    END
  END o_ranQ[100]
  PIN o_ranQ[101]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -159.995 1.355 -159.490 1.435 ;
        RECT -158.690 1.355 -157.785 1.445 ;
        RECT -159.995 1.175 -157.785 1.355 ;
      LAYER mcon ;
        RECT -159.805 1.265 -159.635 1.435 ;
        RECT -158.440 1.265 -158.270 1.435 ;
      LAYER met1 ;
        RECT -159.870 1.170 -158.180 1.470 ;
        RECT -159.690 0.470 -158.690 1.170 ;
    END
  END o_ranQ[101]
  PIN o_ranQ[102]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -164.955 7.165 -162.745 7.345 ;
        RECT -164.955 7.085 -164.450 7.165 ;
        RECT -163.650 7.075 -162.745 7.165 ;
      LAYER mcon ;
        RECT -164.765 7.085 -164.595 7.255 ;
        RECT -163.400 7.085 -163.230 7.255 ;
      LAYER met1 ;
        RECT -164.650 7.350 -163.650 8.050 ;
        RECT -164.830 7.050 -163.140 7.350 ;
    END
  END o_ranQ[102]
  PIN o_ranQ[103]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -169.915 1.355 -169.410 1.435 ;
        RECT -168.610 1.355 -167.705 1.445 ;
        RECT -169.915 1.175 -167.705 1.355 ;
      LAYER mcon ;
        RECT -169.725 1.265 -169.555 1.435 ;
        RECT -168.360 1.265 -168.190 1.435 ;
      LAYER met1 ;
        RECT -169.790 1.170 -168.100 1.470 ;
        RECT -169.610 0.470 -168.610 1.170 ;
    END
  END o_ranQ[103]
  PIN o_ranQ[104]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -174.875 7.165 -172.665 7.345 ;
        RECT -174.875 7.085 -174.370 7.165 ;
        RECT -173.570 7.075 -172.665 7.165 ;
      LAYER mcon ;
        RECT -174.685 7.085 -174.515 7.255 ;
        RECT -173.320 7.085 -173.150 7.255 ;
      LAYER met1 ;
        RECT -174.570 7.350 -173.570 8.050 ;
        RECT -174.750 7.050 -173.060 7.350 ;
    END
  END o_ranQ[104]
  PIN o_ranQ[105]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -179.835 1.355 -179.330 1.435 ;
        RECT -178.530 1.355 -177.625 1.445 ;
        RECT -179.835 1.175 -177.625 1.355 ;
      LAYER mcon ;
        RECT -179.645 1.265 -179.475 1.435 ;
        RECT -178.280 1.265 -178.110 1.435 ;
      LAYER met1 ;
        RECT -179.710 1.170 -178.020 1.470 ;
        RECT -179.530 0.470 -178.530 1.170 ;
    END
  END o_ranQ[105]
  PIN o_ranQ[106]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -184.795 7.165 -182.585 7.345 ;
        RECT -184.795 7.085 -184.290 7.165 ;
        RECT -183.490 7.075 -182.585 7.165 ;
      LAYER mcon ;
        RECT -184.605 7.085 -184.435 7.255 ;
        RECT -183.240 7.085 -183.070 7.255 ;
      LAYER met1 ;
        RECT -184.490 7.350 -183.490 8.050 ;
        RECT -184.670 7.050 -182.980 7.350 ;
    END
  END o_ranQ[106]
  PIN o_ranQ[107]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -189.755 1.355 -189.250 1.435 ;
        RECT -188.450 1.355 -187.545 1.445 ;
        RECT -189.755 1.175 -187.545 1.355 ;
      LAYER mcon ;
        RECT -189.565 1.265 -189.395 1.435 ;
        RECT -188.200 1.265 -188.030 1.435 ;
      LAYER met1 ;
        RECT -189.630 1.170 -187.940 1.470 ;
        RECT -189.450 0.470 -188.450 1.170 ;
    END
  END o_ranQ[107]
  PIN o_ranQ[108]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -194.715 7.165 -192.505 7.345 ;
        RECT -194.715 7.085 -194.210 7.165 ;
        RECT -193.410 7.075 -192.505 7.165 ;
      LAYER mcon ;
        RECT -194.525 7.085 -194.355 7.255 ;
        RECT -193.160 7.085 -192.990 7.255 ;
      LAYER met1 ;
        RECT -194.410 7.350 -193.410 8.050 ;
        RECT -194.590 7.050 -192.900 7.350 ;
    END
  END o_ranQ[108]
  PIN o_ranQ[109]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -199.675 1.355 -199.170 1.435 ;
        RECT -198.370 1.355 -197.465 1.445 ;
        RECT -199.675 1.175 -197.465 1.355 ;
      LAYER mcon ;
        RECT -199.485 1.265 -199.315 1.435 ;
        RECT -198.120 1.265 -197.950 1.435 ;
      LAYER met1 ;
        RECT -199.550 1.170 -197.860 1.470 ;
        RECT -199.370 0.470 -198.370 1.170 ;
    END
  END o_ranQ[109]
  PIN o_ranQ[110]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -204.635 7.165 -202.425 7.345 ;
        RECT -204.635 7.085 -204.130 7.165 ;
        RECT -203.330 7.075 -202.425 7.165 ;
      LAYER mcon ;
        RECT -204.445 7.085 -204.275 7.255 ;
        RECT -203.080 7.085 -202.910 7.255 ;
      LAYER met1 ;
        RECT -204.330 7.350 -203.330 8.050 ;
        RECT -204.510 7.050 -202.820 7.350 ;
    END
  END o_ranQ[110]
  PIN o_ranQ[111]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -209.595 1.355 -209.090 1.435 ;
        RECT -208.290 1.355 -207.385 1.445 ;
        RECT -209.595 1.175 -207.385 1.355 ;
      LAYER mcon ;
        RECT -209.405 1.265 -209.235 1.435 ;
        RECT -208.040 1.265 -207.870 1.435 ;
      LAYER met1 ;
        RECT -209.470 1.170 -207.780 1.470 ;
        RECT -209.290 0.470 -208.290 1.170 ;
    END
  END o_ranQ[111]
  PIN o_ranQ[113]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -219.515 1.355 -219.010 1.435 ;
        RECT -218.210 1.355 -217.305 1.445 ;
        RECT -219.515 1.175 -217.305 1.355 ;
      LAYER mcon ;
        RECT -219.325 1.265 -219.155 1.435 ;
        RECT -217.960 1.265 -217.790 1.435 ;
      LAYER met1 ;
        RECT -219.390 1.170 -217.700 1.470 ;
        RECT -219.210 0.470 -218.210 1.170 ;
    END
  END o_ranQ[113]
  PIN o_ranQ[114]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -224.475 7.165 -222.265 7.345 ;
        RECT -224.475 7.085 -223.970 7.165 ;
        RECT -223.170 7.075 -222.265 7.165 ;
      LAYER mcon ;
        RECT -224.285 7.085 -224.115 7.255 ;
        RECT -222.920 7.085 -222.750 7.255 ;
      LAYER met1 ;
        RECT -224.170 7.350 -223.170 8.050 ;
        RECT -224.350 7.050 -222.660 7.350 ;
    END
  END o_ranQ[114]
  PIN o_ranQ[115]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -229.435 1.355 -228.930 1.435 ;
        RECT -228.130 1.355 -227.225 1.445 ;
        RECT -229.435 1.175 -227.225 1.355 ;
      LAYER mcon ;
        RECT -229.245 1.265 -229.075 1.435 ;
        RECT -227.880 1.265 -227.710 1.435 ;
      LAYER met1 ;
        RECT -229.310 1.170 -227.620 1.470 ;
        RECT -229.130 0.470 -228.130 1.170 ;
    END
  END o_ranQ[115]
  PIN o_ranQ[112]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -214.555 7.165 -212.345 7.345 ;
        RECT -214.555 7.085 -214.050 7.165 ;
        RECT -213.250 7.075 -212.345 7.165 ;
      LAYER mcon ;
        RECT -214.365 7.085 -214.195 7.255 ;
        RECT -213.000 7.085 -212.830 7.255 ;
      LAYER met1 ;
        RECT -214.250 7.350 -213.250 8.050 ;
        RECT -214.430 7.050 -212.740 7.350 ;
    END
  END o_ranQ[112]
  PIN o_ranQ[116]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -234.395 7.165 -232.185 7.345 ;
        RECT -234.395 7.085 -233.890 7.165 ;
        RECT -233.090 7.075 -232.185 7.165 ;
      LAYER mcon ;
        RECT -234.205 7.085 -234.035 7.255 ;
        RECT -232.840 7.085 -232.670 7.255 ;
      LAYER met1 ;
        RECT -234.090 7.350 -233.090 8.050 ;
        RECT -234.270 7.050 -232.580 7.350 ;
    END
  END o_ranQ[116]
  PIN o_ranQ[117]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -239.355 1.355 -238.850 1.435 ;
        RECT -238.050 1.355 -237.145 1.445 ;
        RECT -239.355 1.175 -237.145 1.355 ;
      LAYER mcon ;
        RECT -239.165 1.265 -238.995 1.435 ;
        RECT -237.800 1.265 -237.630 1.435 ;
      LAYER met1 ;
        RECT -239.230 1.170 -237.540 1.470 ;
        RECT -239.050 0.470 -238.050 1.170 ;
    END
  END o_ranQ[117]
  PIN o_ranQ[118]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -244.315 7.165 -242.105 7.345 ;
        RECT -244.315 7.085 -243.810 7.165 ;
        RECT -243.010 7.075 -242.105 7.165 ;
      LAYER mcon ;
        RECT -244.125 7.085 -243.955 7.255 ;
        RECT -242.760 7.085 -242.590 7.255 ;
      LAYER met1 ;
        RECT -244.010 7.350 -243.010 8.050 ;
        RECT -244.190 7.050 -242.500 7.350 ;
    END
  END o_ranQ[118]
  PIN o_ranQ[119]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -249.275 1.355 -248.770 1.435 ;
        RECT -247.970 1.355 -247.065 1.445 ;
        RECT -249.275 1.175 -247.065 1.355 ;
      LAYER mcon ;
        RECT -249.085 1.265 -248.915 1.435 ;
        RECT -247.720 1.265 -247.550 1.435 ;
      LAYER met1 ;
        RECT -249.150 1.170 -247.460 1.470 ;
        RECT -248.970 0.470 -247.970 1.170 ;
    END
  END o_ranQ[119]
  PIN o_ranQ[120]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -254.235 7.165 -252.025 7.345 ;
        RECT -254.235 7.085 -253.730 7.165 ;
        RECT -252.930 7.075 -252.025 7.165 ;
      LAYER mcon ;
        RECT -254.045 7.085 -253.875 7.255 ;
        RECT -252.680 7.085 -252.510 7.255 ;
      LAYER met1 ;
        RECT -253.930 7.350 -252.930 8.050 ;
        RECT -254.110 7.050 -252.420 7.350 ;
    END
  END o_ranQ[120]
  PIN o_ranQ[121]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -259.195 1.355 -258.690 1.435 ;
        RECT -257.890 1.355 -256.985 1.445 ;
        RECT -259.195 1.175 -256.985 1.355 ;
      LAYER mcon ;
        RECT -259.005 1.265 -258.835 1.435 ;
        RECT -257.640 1.265 -257.470 1.435 ;
      LAYER met1 ;
        RECT -259.070 1.170 -257.380 1.470 ;
        RECT -258.890 0.470 -257.890 1.170 ;
    END
  END o_ranQ[121]
  PIN o_ranQ[122]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -264.155 7.165 -261.945 7.345 ;
        RECT -264.155 7.085 -263.650 7.165 ;
        RECT -262.850 7.075 -261.945 7.165 ;
      LAYER mcon ;
        RECT -263.965 7.085 -263.795 7.255 ;
        RECT -262.600 7.085 -262.430 7.255 ;
      LAYER met1 ;
        RECT -263.850 7.350 -262.850 8.050 ;
        RECT -264.030 7.050 -262.340 7.350 ;
    END
  END o_ranQ[122]
  PIN o_ranQ[123]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -269.115 1.355 -268.610 1.435 ;
        RECT -267.810 1.355 -266.905 1.445 ;
        RECT -269.115 1.175 -266.905 1.355 ;
      LAYER mcon ;
        RECT -268.925 1.265 -268.755 1.435 ;
        RECT -267.560 1.265 -267.390 1.435 ;
      LAYER met1 ;
        RECT -268.990 1.170 -267.300 1.470 ;
        RECT -268.810 0.470 -267.810 1.170 ;
    END
  END o_ranQ[123]
  PIN o_ranQ[125]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -279.035 1.355 -278.530 1.435 ;
        RECT -277.730 1.355 -276.825 1.445 ;
        RECT -279.035 1.175 -276.825 1.355 ;
      LAYER mcon ;
        RECT -278.845 1.265 -278.675 1.435 ;
        RECT -277.480 1.265 -277.310 1.435 ;
      LAYER met1 ;
        RECT -278.910 1.170 -277.220 1.470 ;
        RECT -278.730 0.470 -277.730 1.170 ;
    END
  END o_ranQ[125]
  PIN o_ranQ[126]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -283.995 7.165 -281.785 7.345 ;
        RECT -283.995 7.085 -283.490 7.165 ;
        RECT -282.690 7.075 -281.785 7.165 ;
      LAYER mcon ;
        RECT -283.805 7.085 -283.635 7.255 ;
        RECT -282.440 7.085 -282.270 7.255 ;
      LAYER met1 ;
        RECT -283.690 7.350 -282.690 8.050 ;
        RECT -283.870 7.050 -282.180 7.350 ;
    END
  END o_ranQ[126]
  PIN o_ranQ[127]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -288.955 1.355 -288.450 1.435 ;
        RECT -287.650 1.355 -286.745 1.445 ;
        RECT -288.955 1.175 -286.745 1.355 ;
      LAYER mcon ;
        RECT -288.765 1.265 -288.595 1.435 ;
        RECT -287.400 1.265 -287.230 1.435 ;
      LAYER met1 ;
        RECT -288.830 1.170 -287.140 1.470 ;
        RECT -288.650 0.470 -287.650 1.170 ;
    END
  END o_ranQ[127]
  PIN o_ranQ[188]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -272.315 -86.185 -270.105 -86.005 ;
        RECT -272.315 -86.265 -271.810 -86.185 ;
        RECT -271.010 -86.275 -270.105 -86.185 ;
      LAYER mcon ;
        RECT -272.125 -86.265 -271.955 -86.095 ;
        RECT -270.760 -86.265 -270.590 -86.095 ;
      LAYER met1 ;
        RECT -272.010 -86.000 -271.010 -85.300 ;
        RECT -272.190 -86.300 -270.500 -86.000 ;
    END
  END o_ranQ[188]
  PIN o_ranQ[129]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 20.325 -91.995 20.830 -91.915 ;
        RECT 21.630 -91.995 22.535 -91.905 ;
        RECT 20.325 -92.175 22.535 -91.995 ;
      LAYER mcon ;
        RECT 20.515 -92.085 20.685 -91.915 ;
        RECT 21.880 -92.085 22.050 -91.915 ;
      LAYER met1 ;
        RECT 20.450 -92.180 22.140 -91.880 ;
        RECT 20.630 -92.880 21.630 -92.180 ;
    END
  END o_ranQ[129]
  PIN o_ranQ[130]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 15.365 -86.185 17.575 -86.005 ;
        RECT 15.365 -86.265 15.870 -86.185 ;
        RECT 16.670 -86.275 17.575 -86.185 ;
      LAYER mcon ;
        RECT 15.555 -86.265 15.725 -86.095 ;
        RECT 16.920 -86.265 17.090 -86.095 ;
      LAYER met1 ;
        RECT 15.670 -86.000 16.670 -85.300 ;
        RECT 15.490 -86.300 17.180 -86.000 ;
    END
  END o_ranQ[130]
  PIN o_ranQ[131]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 10.405 -91.995 10.910 -91.915 ;
        RECT 11.710 -91.995 12.615 -91.905 ;
        RECT 10.405 -92.175 12.615 -91.995 ;
      LAYER mcon ;
        RECT 10.595 -92.085 10.765 -91.915 ;
        RECT 11.960 -92.085 12.130 -91.915 ;
      LAYER met1 ;
        RECT 10.530 -92.180 12.220 -91.880 ;
        RECT 10.710 -92.880 11.710 -92.180 ;
    END
  END o_ranQ[131]
  PIN o_ranQ[128]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 25.285 -86.185 27.495 -86.005 ;
        RECT 25.285 -86.265 25.790 -86.185 ;
        RECT 26.590 -86.275 27.495 -86.185 ;
      LAYER mcon ;
        RECT 25.475 -86.265 25.645 -86.095 ;
        RECT 26.840 -86.265 27.010 -86.095 ;
      LAYER met1 ;
        RECT 25.590 -86.000 26.590 -85.300 ;
        RECT 25.410 -86.300 27.100 -86.000 ;
    END
  END o_ranQ[128]
  PIN o_ranQ[132]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 5.445 -86.185 7.655 -86.005 ;
        RECT 5.445 -86.265 5.950 -86.185 ;
        RECT 6.750 -86.275 7.655 -86.185 ;
      LAYER mcon ;
        RECT 5.635 -86.265 5.805 -86.095 ;
        RECT 7.000 -86.265 7.170 -86.095 ;
      LAYER met1 ;
        RECT 5.750 -86.000 6.750 -85.300 ;
        RECT 5.570 -86.300 7.260 -86.000 ;
    END
  END o_ranQ[132]
  PIN o_ranQ[133]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 0.485 -91.995 0.990 -91.915 ;
        RECT 1.790 -91.995 2.695 -91.905 ;
        RECT 0.485 -92.175 2.695 -91.995 ;
      LAYER mcon ;
        RECT 0.675 -92.085 0.845 -91.915 ;
        RECT 2.040 -92.085 2.210 -91.915 ;
      LAYER met1 ;
        RECT 0.610 -92.180 2.300 -91.880 ;
        RECT 0.790 -92.880 1.790 -92.180 ;
    END
  END o_ranQ[133]
  PIN o_ranQ[134]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -4.475 -86.185 -2.265 -86.005 ;
        RECT -4.475 -86.265 -3.970 -86.185 ;
        RECT -3.170 -86.275 -2.265 -86.185 ;
      LAYER mcon ;
        RECT -4.285 -86.265 -4.115 -86.095 ;
        RECT -2.920 -86.265 -2.750 -86.095 ;
      LAYER met1 ;
        RECT -4.170 -86.000 -3.170 -85.300 ;
        RECT -4.350 -86.300 -2.660 -86.000 ;
    END
  END o_ranQ[134]
  PIN o_ranQ[135]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -9.435 -91.995 -8.930 -91.915 ;
        RECT -8.130 -91.995 -7.225 -91.905 ;
        RECT -9.435 -92.175 -7.225 -91.995 ;
      LAYER mcon ;
        RECT -9.245 -92.085 -9.075 -91.915 ;
        RECT -7.880 -92.085 -7.710 -91.915 ;
      LAYER met1 ;
        RECT -9.310 -92.180 -7.620 -91.880 ;
        RECT -9.130 -92.880 -8.130 -92.180 ;
    END
  END o_ranQ[135]
  PIN o_ranQ[136]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -14.395 -86.185 -12.185 -86.005 ;
        RECT -14.395 -86.265 -13.890 -86.185 ;
        RECT -13.090 -86.275 -12.185 -86.185 ;
      LAYER mcon ;
        RECT -14.205 -86.265 -14.035 -86.095 ;
        RECT -12.840 -86.265 -12.670 -86.095 ;
      LAYER met1 ;
        RECT -14.090 -86.000 -13.090 -85.300 ;
        RECT -14.270 -86.300 -12.580 -86.000 ;
    END
  END o_ranQ[136]
  PIN o_ranQ[137]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -19.355 -91.995 -18.850 -91.915 ;
        RECT -18.050 -91.995 -17.145 -91.905 ;
        RECT -19.355 -92.175 -17.145 -91.995 ;
      LAYER mcon ;
        RECT -19.165 -92.085 -18.995 -91.915 ;
        RECT -17.800 -92.085 -17.630 -91.915 ;
      LAYER met1 ;
        RECT -19.230 -92.180 -17.540 -91.880 ;
        RECT -19.050 -92.880 -18.050 -92.180 ;
    END
  END o_ranQ[137]
  PIN o_ranQ[138]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -24.315 -86.185 -22.105 -86.005 ;
        RECT -24.315 -86.265 -23.810 -86.185 ;
        RECT -23.010 -86.275 -22.105 -86.185 ;
      LAYER mcon ;
        RECT -24.125 -86.265 -23.955 -86.095 ;
        RECT -22.760 -86.265 -22.590 -86.095 ;
      LAYER met1 ;
        RECT -24.010 -86.000 -23.010 -85.300 ;
        RECT -24.190 -86.300 -22.500 -86.000 ;
    END
  END o_ranQ[138]
  PIN o_ranQ[139]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -29.275 -91.995 -28.770 -91.915 ;
        RECT -27.970 -91.995 -27.065 -91.905 ;
        RECT -29.275 -92.175 -27.065 -91.995 ;
      LAYER mcon ;
        RECT -29.085 -92.085 -28.915 -91.915 ;
        RECT -27.720 -92.085 -27.550 -91.915 ;
      LAYER met1 ;
        RECT -29.150 -92.180 -27.460 -91.880 ;
        RECT -28.970 -92.880 -27.970 -92.180 ;
    END
  END o_ranQ[139]
  PIN o_ranQ[140]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -34.235 -86.185 -32.025 -86.005 ;
        RECT -34.235 -86.265 -33.730 -86.185 ;
        RECT -32.930 -86.275 -32.025 -86.185 ;
      LAYER mcon ;
        RECT -34.045 -86.265 -33.875 -86.095 ;
        RECT -32.680 -86.265 -32.510 -86.095 ;
      LAYER met1 ;
        RECT -33.930 -86.000 -32.930 -85.300 ;
        RECT -34.110 -86.300 -32.420 -86.000 ;
    END
  END o_ranQ[140]
  PIN o_ranQ[141]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -39.195 -91.995 -38.690 -91.915 ;
        RECT -37.890 -91.995 -36.985 -91.905 ;
        RECT -39.195 -92.175 -36.985 -91.995 ;
      LAYER mcon ;
        RECT -39.005 -92.085 -38.835 -91.915 ;
        RECT -37.640 -92.085 -37.470 -91.915 ;
      LAYER met1 ;
        RECT -39.070 -92.180 -37.380 -91.880 ;
        RECT -38.890 -92.880 -37.890 -92.180 ;
    END
  END o_ranQ[141]
  PIN o_ranQ[142]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -44.155 -86.185 -41.945 -86.005 ;
        RECT -44.155 -86.265 -43.650 -86.185 ;
        RECT -42.850 -86.275 -41.945 -86.185 ;
      LAYER mcon ;
        RECT -43.965 -86.265 -43.795 -86.095 ;
        RECT -42.600 -86.265 -42.430 -86.095 ;
      LAYER met1 ;
        RECT -43.850 -86.000 -42.850 -85.300 ;
        RECT -44.030 -86.300 -42.340 -86.000 ;
    END
  END o_ranQ[142]
  PIN o_ranQ[143]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -49.115 -91.995 -48.610 -91.915 ;
        RECT -47.810 -91.995 -46.905 -91.905 ;
        RECT -49.115 -92.175 -46.905 -91.995 ;
      LAYER mcon ;
        RECT -48.925 -92.085 -48.755 -91.915 ;
        RECT -47.560 -92.085 -47.390 -91.915 ;
      LAYER met1 ;
        RECT -48.990 -92.180 -47.300 -91.880 ;
        RECT -48.810 -92.880 -47.810 -92.180 ;
    END
  END o_ranQ[143]
  PIN o_ranQ[145]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -59.035 -91.995 -58.530 -91.915 ;
        RECT -57.730 -91.995 -56.825 -91.905 ;
        RECT -59.035 -92.175 -56.825 -91.995 ;
      LAYER mcon ;
        RECT -58.845 -92.085 -58.675 -91.915 ;
        RECT -57.480 -92.085 -57.310 -91.915 ;
      LAYER met1 ;
        RECT -58.910 -92.180 -57.220 -91.880 ;
        RECT -58.730 -92.880 -57.730 -92.180 ;
    END
  END o_ranQ[145]
  PIN o_ranQ[146]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -63.995 -86.185 -61.785 -86.005 ;
        RECT -63.995 -86.265 -63.490 -86.185 ;
        RECT -62.690 -86.275 -61.785 -86.185 ;
      LAYER mcon ;
        RECT -63.805 -86.265 -63.635 -86.095 ;
        RECT -62.440 -86.265 -62.270 -86.095 ;
      LAYER met1 ;
        RECT -63.690 -86.000 -62.690 -85.300 ;
        RECT -63.870 -86.300 -62.180 -86.000 ;
    END
  END o_ranQ[146]
  PIN o_ranQ[147]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -68.955 -91.995 -68.450 -91.915 ;
        RECT -67.650 -91.995 -66.745 -91.905 ;
        RECT -68.955 -92.175 -66.745 -91.995 ;
      LAYER mcon ;
        RECT -68.765 -92.085 -68.595 -91.915 ;
        RECT -67.400 -92.085 -67.230 -91.915 ;
      LAYER met1 ;
        RECT -68.830 -92.180 -67.140 -91.880 ;
        RECT -68.650 -92.880 -67.650 -92.180 ;
    END
  END o_ranQ[147]
  PIN o_ranQ[144]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -54.075 -86.185 -51.865 -86.005 ;
        RECT -54.075 -86.265 -53.570 -86.185 ;
        RECT -52.770 -86.275 -51.865 -86.185 ;
      LAYER mcon ;
        RECT -53.885 -86.265 -53.715 -86.095 ;
        RECT -52.520 -86.265 -52.350 -86.095 ;
      LAYER met1 ;
        RECT -53.770 -86.000 -52.770 -85.300 ;
        RECT -53.950 -86.300 -52.260 -86.000 ;
    END
  END o_ranQ[144]
  PIN o_ranQ[148]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -73.915 -86.185 -71.705 -86.005 ;
        RECT -73.915 -86.265 -73.410 -86.185 ;
        RECT -72.610 -86.275 -71.705 -86.185 ;
      LAYER mcon ;
        RECT -73.725 -86.265 -73.555 -86.095 ;
        RECT -72.360 -86.265 -72.190 -86.095 ;
      LAYER met1 ;
        RECT -73.610 -86.000 -72.610 -85.300 ;
        RECT -73.790 -86.300 -72.100 -86.000 ;
    END
  END o_ranQ[148]
  PIN o_ranQ[149]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -78.875 -91.995 -78.370 -91.915 ;
        RECT -77.570 -91.995 -76.665 -91.905 ;
        RECT -78.875 -92.175 -76.665 -91.995 ;
      LAYER mcon ;
        RECT -78.685 -92.085 -78.515 -91.915 ;
        RECT -77.320 -92.085 -77.150 -91.915 ;
      LAYER met1 ;
        RECT -78.750 -92.180 -77.060 -91.880 ;
        RECT -78.570 -92.880 -77.570 -92.180 ;
    END
  END o_ranQ[149]
  PIN o_ranQ[150]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -83.835 -86.185 -81.625 -86.005 ;
        RECT -83.835 -86.265 -83.330 -86.185 ;
        RECT -82.530 -86.275 -81.625 -86.185 ;
      LAYER mcon ;
        RECT -83.645 -86.265 -83.475 -86.095 ;
        RECT -82.280 -86.265 -82.110 -86.095 ;
      LAYER met1 ;
        RECT -83.530 -86.000 -82.530 -85.300 ;
        RECT -83.710 -86.300 -82.020 -86.000 ;
    END
  END o_ranQ[150]
  PIN o_ranQ[151]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -88.795 -91.995 -88.290 -91.915 ;
        RECT -87.490 -91.995 -86.585 -91.905 ;
        RECT -88.795 -92.175 -86.585 -91.995 ;
      LAYER mcon ;
        RECT -88.605 -92.085 -88.435 -91.915 ;
        RECT -87.240 -92.085 -87.070 -91.915 ;
      LAYER met1 ;
        RECT -88.670 -92.180 -86.980 -91.880 ;
        RECT -88.490 -92.880 -87.490 -92.180 ;
    END
  END o_ranQ[151]
  PIN o_ranQ[152]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -93.755 -86.185 -91.545 -86.005 ;
        RECT -93.755 -86.265 -93.250 -86.185 ;
        RECT -92.450 -86.275 -91.545 -86.185 ;
      LAYER mcon ;
        RECT -93.565 -86.265 -93.395 -86.095 ;
        RECT -92.200 -86.265 -92.030 -86.095 ;
      LAYER met1 ;
        RECT -93.450 -86.000 -92.450 -85.300 ;
        RECT -93.630 -86.300 -91.940 -86.000 ;
    END
  END o_ranQ[152]
  PIN o_ranQ[153]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -98.715 -91.995 -98.210 -91.915 ;
        RECT -97.410 -91.995 -96.505 -91.905 ;
        RECT -98.715 -92.175 -96.505 -91.995 ;
      LAYER mcon ;
        RECT -98.525 -92.085 -98.355 -91.915 ;
        RECT -97.160 -92.085 -96.990 -91.915 ;
      LAYER met1 ;
        RECT -98.590 -92.180 -96.900 -91.880 ;
        RECT -98.410 -92.880 -97.410 -92.180 ;
    END
  END o_ranQ[153]
  PIN o_ranQ[154]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -103.675 -86.185 -101.465 -86.005 ;
        RECT -103.675 -86.265 -103.170 -86.185 ;
        RECT -102.370 -86.275 -101.465 -86.185 ;
      LAYER mcon ;
        RECT -103.485 -86.265 -103.315 -86.095 ;
        RECT -102.120 -86.265 -101.950 -86.095 ;
      LAYER met1 ;
        RECT -103.370 -86.000 -102.370 -85.300 ;
        RECT -103.550 -86.300 -101.860 -86.000 ;
    END
  END o_ranQ[154]
  PIN o_ranQ[155]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -108.635 -91.995 -108.130 -91.915 ;
        RECT -107.330 -91.995 -106.425 -91.905 ;
        RECT -108.635 -92.175 -106.425 -91.995 ;
      LAYER mcon ;
        RECT -108.445 -92.085 -108.275 -91.915 ;
        RECT -107.080 -92.085 -106.910 -91.915 ;
      LAYER met1 ;
        RECT -108.510 -92.180 -106.820 -91.880 ;
        RECT -108.330 -92.880 -107.330 -92.180 ;
    END
  END o_ranQ[155]
  PIN o_ranQ[156]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -113.595 -86.185 -111.385 -86.005 ;
        RECT -113.595 -86.265 -113.090 -86.185 ;
        RECT -112.290 -86.275 -111.385 -86.185 ;
      LAYER mcon ;
        RECT -113.405 -86.265 -113.235 -86.095 ;
        RECT -112.040 -86.265 -111.870 -86.095 ;
      LAYER met1 ;
        RECT -113.290 -86.000 -112.290 -85.300 ;
        RECT -113.470 -86.300 -111.780 -86.000 ;
    END
  END o_ranQ[156]
  PIN o_ranQ[157]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -118.555 -91.995 -118.050 -91.915 ;
        RECT -117.250 -91.995 -116.345 -91.905 ;
        RECT -118.555 -92.175 -116.345 -91.995 ;
      LAYER mcon ;
        RECT -118.365 -92.085 -118.195 -91.915 ;
        RECT -117.000 -92.085 -116.830 -91.915 ;
      LAYER met1 ;
        RECT -118.430 -92.180 -116.740 -91.880 ;
        RECT -118.250 -92.880 -117.250 -92.180 ;
    END
  END o_ranQ[157]
  PIN o_ranQ[158]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -123.515 -86.185 -121.305 -86.005 ;
        RECT -123.515 -86.265 -123.010 -86.185 ;
        RECT -122.210 -86.275 -121.305 -86.185 ;
      LAYER mcon ;
        RECT -123.325 -86.265 -123.155 -86.095 ;
        RECT -121.960 -86.265 -121.790 -86.095 ;
      LAYER met1 ;
        RECT -123.210 -86.000 -122.210 -85.300 ;
        RECT -123.390 -86.300 -121.700 -86.000 ;
    END
  END o_ranQ[158]
  PIN o_ranQ[159]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -128.475 -91.995 -127.970 -91.915 ;
        RECT -127.170 -91.995 -126.265 -91.905 ;
        RECT -128.475 -92.175 -126.265 -91.995 ;
      LAYER mcon ;
        RECT -128.285 -92.085 -128.115 -91.915 ;
        RECT -126.920 -92.085 -126.750 -91.915 ;
      LAYER met1 ;
        RECT -128.350 -92.180 -126.660 -91.880 ;
        RECT -128.170 -92.880 -127.170 -92.180 ;
    END
  END o_ranQ[159]
  PIN o_ranQ[161]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -138.395 -91.995 -137.890 -91.915 ;
        RECT -137.090 -91.995 -136.185 -91.905 ;
        RECT -138.395 -92.175 -136.185 -91.995 ;
      LAYER mcon ;
        RECT -138.205 -92.085 -138.035 -91.915 ;
        RECT -136.840 -92.085 -136.670 -91.915 ;
      LAYER met1 ;
        RECT -138.270 -92.180 -136.580 -91.880 ;
        RECT -138.090 -92.880 -137.090 -92.180 ;
    END
  END o_ranQ[161]
  PIN o_ranQ[162]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -143.355 -86.185 -141.145 -86.005 ;
        RECT -143.355 -86.265 -142.850 -86.185 ;
        RECT -142.050 -86.275 -141.145 -86.185 ;
      LAYER mcon ;
        RECT -143.165 -86.265 -142.995 -86.095 ;
        RECT -141.800 -86.265 -141.630 -86.095 ;
      LAYER met1 ;
        RECT -143.050 -86.000 -142.050 -85.300 ;
        RECT -143.230 -86.300 -141.540 -86.000 ;
    END
  END o_ranQ[162]
  PIN o_ranQ[163]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -148.315 -91.995 -147.810 -91.915 ;
        RECT -147.010 -91.995 -146.105 -91.905 ;
        RECT -148.315 -92.175 -146.105 -91.995 ;
      LAYER mcon ;
        RECT -148.125 -92.085 -147.955 -91.915 ;
        RECT -146.760 -92.085 -146.590 -91.915 ;
      LAYER met1 ;
        RECT -148.190 -92.180 -146.500 -91.880 ;
        RECT -148.010 -92.880 -147.010 -92.180 ;
    END
  END o_ranQ[163]
  PIN o_ranQ[160]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -133.435 -86.185 -131.225 -86.005 ;
        RECT -133.435 -86.265 -132.930 -86.185 ;
        RECT -132.130 -86.275 -131.225 -86.185 ;
      LAYER mcon ;
        RECT -133.245 -86.265 -133.075 -86.095 ;
        RECT -131.880 -86.265 -131.710 -86.095 ;
      LAYER met1 ;
        RECT -133.130 -86.000 -132.130 -85.300 ;
        RECT -133.310 -86.300 -131.620 -86.000 ;
    END
  END o_ranQ[160]
  PIN o_ranQ[164]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -153.275 -86.185 -151.065 -86.005 ;
        RECT -153.275 -86.265 -152.770 -86.185 ;
        RECT -151.970 -86.275 -151.065 -86.185 ;
      LAYER mcon ;
        RECT -153.085 -86.265 -152.915 -86.095 ;
        RECT -151.720 -86.265 -151.550 -86.095 ;
      LAYER met1 ;
        RECT -152.970 -86.000 -151.970 -85.300 ;
        RECT -153.150 -86.300 -151.460 -86.000 ;
    END
  END o_ranQ[164]
  PIN o_ranQ[165]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -158.235 -91.995 -157.730 -91.915 ;
        RECT -156.930 -91.995 -156.025 -91.905 ;
        RECT -158.235 -92.175 -156.025 -91.995 ;
      LAYER mcon ;
        RECT -158.045 -92.085 -157.875 -91.915 ;
        RECT -156.680 -92.085 -156.510 -91.915 ;
      LAYER met1 ;
        RECT -158.110 -92.180 -156.420 -91.880 ;
        RECT -157.930 -92.880 -156.930 -92.180 ;
    END
  END o_ranQ[165]
  PIN o_ranQ[166]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -163.195 -86.185 -160.985 -86.005 ;
        RECT -163.195 -86.265 -162.690 -86.185 ;
        RECT -161.890 -86.275 -160.985 -86.185 ;
      LAYER mcon ;
        RECT -163.005 -86.265 -162.835 -86.095 ;
        RECT -161.640 -86.265 -161.470 -86.095 ;
      LAYER met1 ;
        RECT -162.890 -86.000 -161.890 -85.300 ;
        RECT -163.070 -86.300 -161.380 -86.000 ;
    END
  END o_ranQ[166]
  PIN o_ranQ[167]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -168.155 -91.995 -167.650 -91.915 ;
        RECT -166.850 -91.995 -165.945 -91.905 ;
        RECT -168.155 -92.175 -165.945 -91.995 ;
      LAYER mcon ;
        RECT -167.965 -92.085 -167.795 -91.915 ;
        RECT -166.600 -92.085 -166.430 -91.915 ;
      LAYER met1 ;
        RECT -168.030 -92.180 -166.340 -91.880 ;
        RECT -167.850 -92.880 -166.850 -92.180 ;
    END
  END o_ranQ[167]
  PIN o_ranQ[168]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -173.115 -86.185 -170.905 -86.005 ;
        RECT -173.115 -86.265 -172.610 -86.185 ;
        RECT -171.810 -86.275 -170.905 -86.185 ;
      LAYER mcon ;
        RECT -172.925 -86.265 -172.755 -86.095 ;
        RECT -171.560 -86.265 -171.390 -86.095 ;
      LAYER met1 ;
        RECT -172.810 -86.000 -171.810 -85.300 ;
        RECT -172.990 -86.300 -171.300 -86.000 ;
    END
  END o_ranQ[168]
  PIN o_ranQ[169]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -178.075 -91.995 -177.570 -91.915 ;
        RECT -176.770 -91.995 -175.865 -91.905 ;
        RECT -178.075 -92.175 -175.865 -91.995 ;
      LAYER mcon ;
        RECT -177.885 -92.085 -177.715 -91.915 ;
        RECT -176.520 -92.085 -176.350 -91.915 ;
      LAYER met1 ;
        RECT -177.950 -92.180 -176.260 -91.880 ;
        RECT -177.770 -92.880 -176.770 -92.180 ;
    END
  END o_ranQ[169]
  PIN o_ranQ[170]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -183.035 -86.185 -180.825 -86.005 ;
        RECT -183.035 -86.265 -182.530 -86.185 ;
        RECT -181.730 -86.275 -180.825 -86.185 ;
      LAYER mcon ;
        RECT -182.845 -86.265 -182.675 -86.095 ;
        RECT -181.480 -86.265 -181.310 -86.095 ;
      LAYER met1 ;
        RECT -182.730 -86.000 -181.730 -85.300 ;
        RECT -182.910 -86.300 -181.220 -86.000 ;
    END
  END o_ranQ[170]
  PIN o_ranQ[171]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -187.995 -91.995 -187.490 -91.915 ;
        RECT -186.690 -91.995 -185.785 -91.905 ;
        RECT -187.995 -92.175 -185.785 -91.995 ;
      LAYER mcon ;
        RECT -187.805 -92.085 -187.635 -91.915 ;
        RECT -186.440 -92.085 -186.270 -91.915 ;
      LAYER met1 ;
        RECT -187.870 -92.180 -186.180 -91.880 ;
        RECT -187.690 -92.880 -186.690 -92.180 ;
    END
  END o_ranQ[171]
  PIN o_ranQ[172]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -192.955 -86.185 -190.745 -86.005 ;
        RECT -192.955 -86.265 -192.450 -86.185 ;
        RECT -191.650 -86.275 -190.745 -86.185 ;
      LAYER mcon ;
        RECT -192.765 -86.265 -192.595 -86.095 ;
        RECT -191.400 -86.265 -191.230 -86.095 ;
      LAYER met1 ;
        RECT -192.650 -86.000 -191.650 -85.300 ;
        RECT -192.830 -86.300 -191.140 -86.000 ;
    END
  END o_ranQ[172]
  PIN o_ranQ[173]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -197.915 -91.995 -197.410 -91.915 ;
        RECT -196.610 -91.995 -195.705 -91.905 ;
        RECT -197.915 -92.175 -195.705 -91.995 ;
      LAYER mcon ;
        RECT -197.725 -92.085 -197.555 -91.915 ;
        RECT -196.360 -92.085 -196.190 -91.915 ;
      LAYER met1 ;
        RECT -197.790 -92.180 -196.100 -91.880 ;
        RECT -197.610 -92.880 -196.610 -92.180 ;
    END
  END o_ranQ[173]
  PIN o_ranQ[174]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -202.875 -86.185 -200.665 -86.005 ;
        RECT -202.875 -86.265 -202.370 -86.185 ;
        RECT -201.570 -86.275 -200.665 -86.185 ;
      LAYER mcon ;
        RECT -202.685 -86.265 -202.515 -86.095 ;
        RECT -201.320 -86.265 -201.150 -86.095 ;
      LAYER met1 ;
        RECT -202.570 -86.000 -201.570 -85.300 ;
        RECT -202.750 -86.300 -201.060 -86.000 ;
    END
  END o_ranQ[174]
  PIN o_ranQ[175]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -207.835 -91.995 -207.330 -91.915 ;
        RECT -206.530 -91.995 -205.625 -91.905 ;
        RECT -207.835 -92.175 -205.625 -91.995 ;
      LAYER mcon ;
        RECT -207.645 -92.085 -207.475 -91.915 ;
        RECT -206.280 -92.085 -206.110 -91.915 ;
      LAYER met1 ;
        RECT -207.710 -92.180 -206.020 -91.880 ;
        RECT -207.530 -92.880 -206.530 -92.180 ;
    END
  END o_ranQ[175]
  PIN o_ranQ[177]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -217.755 -91.995 -217.250 -91.915 ;
        RECT -216.450 -91.995 -215.545 -91.905 ;
        RECT -217.755 -92.175 -215.545 -91.995 ;
      LAYER mcon ;
        RECT -217.565 -92.085 -217.395 -91.915 ;
        RECT -216.200 -92.085 -216.030 -91.915 ;
      LAYER met1 ;
        RECT -217.630 -92.180 -215.940 -91.880 ;
        RECT -217.450 -92.880 -216.450 -92.180 ;
    END
  END o_ranQ[177]
  PIN o_ranQ[178]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -222.715 -86.185 -220.505 -86.005 ;
        RECT -222.715 -86.265 -222.210 -86.185 ;
        RECT -221.410 -86.275 -220.505 -86.185 ;
      LAYER mcon ;
        RECT -222.525 -86.265 -222.355 -86.095 ;
        RECT -221.160 -86.265 -220.990 -86.095 ;
      LAYER met1 ;
        RECT -222.410 -86.000 -221.410 -85.300 ;
        RECT -222.590 -86.300 -220.900 -86.000 ;
    END
  END o_ranQ[178]
  PIN o_ranQ[179]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -227.675 -91.995 -227.170 -91.915 ;
        RECT -226.370 -91.995 -225.465 -91.905 ;
        RECT -227.675 -92.175 -225.465 -91.995 ;
      LAYER mcon ;
        RECT -227.485 -92.085 -227.315 -91.915 ;
        RECT -226.120 -92.085 -225.950 -91.915 ;
      LAYER met1 ;
        RECT -227.550 -92.180 -225.860 -91.880 ;
        RECT -227.370 -92.880 -226.370 -92.180 ;
    END
  END o_ranQ[179]
  PIN o_ranQ[176]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -212.795 -86.185 -210.585 -86.005 ;
        RECT -212.795 -86.265 -212.290 -86.185 ;
        RECT -211.490 -86.275 -210.585 -86.185 ;
      LAYER mcon ;
        RECT -212.605 -86.265 -212.435 -86.095 ;
        RECT -211.240 -86.265 -211.070 -86.095 ;
      LAYER met1 ;
        RECT -212.490 -86.000 -211.490 -85.300 ;
        RECT -212.670 -86.300 -210.980 -86.000 ;
    END
  END o_ranQ[176]
  PIN o_ranQ[180]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -232.635 -86.185 -230.425 -86.005 ;
        RECT -232.635 -86.265 -232.130 -86.185 ;
        RECT -231.330 -86.275 -230.425 -86.185 ;
      LAYER mcon ;
        RECT -232.445 -86.265 -232.275 -86.095 ;
        RECT -231.080 -86.265 -230.910 -86.095 ;
      LAYER met1 ;
        RECT -232.330 -86.000 -231.330 -85.300 ;
        RECT -232.510 -86.300 -230.820 -86.000 ;
    END
  END o_ranQ[180]
  PIN o_ranQ[181]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -237.595 -91.995 -237.090 -91.915 ;
        RECT -236.290 -91.995 -235.385 -91.905 ;
        RECT -237.595 -92.175 -235.385 -91.995 ;
      LAYER mcon ;
        RECT -237.405 -92.085 -237.235 -91.915 ;
        RECT -236.040 -92.085 -235.870 -91.915 ;
      LAYER met1 ;
        RECT -237.470 -92.180 -235.780 -91.880 ;
        RECT -237.290 -92.880 -236.290 -92.180 ;
    END
  END o_ranQ[181]
  PIN o_ranQ[182]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -242.555 -86.185 -240.345 -86.005 ;
        RECT -242.555 -86.265 -242.050 -86.185 ;
        RECT -241.250 -86.275 -240.345 -86.185 ;
      LAYER mcon ;
        RECT -242.365 -86.265 -242.195 -86.095 ;
        RECT -241.000 -86.265 -240.830 -86.095 ;
      LAYER met1 ;
        RECT -242.250 -86.000 -241.250 -85.300 ;
        RECT -242.430 -86.300 -240.740 -86.000 ;
    END
  END o_ranQ[182]
  PIN o_ranQ[183]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -247.515 -91.995 -247.010 -91.915 ;
        RECT -246.210 -91.995 -245.305 -91.905 ;
        RECT -247.515 -92.175 -245.305 -91.995 ;
      LAYER mcon ;
        RECT -247.325 -92.085 -247.155 -91.915 ;
        RECT -245.960 -92.085 -245.790 -91.915 ;
      LAYER met1 ;
        RECT -247.390 -92.180 -245.700 -91.880 ;
        RECT -247.210 -92.880 -246.210 -92.180 ;
    END
  END o_ranQ[183]
  PIN o_ranQ[184]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -252.475 -86.185 -250.265 -86.005 ;
        RECT -252.475 -86.265 -251.970 -86.185 ;
        RECT -251.170 -86.275 -250.265 -86.185 ;
      LAYER mcon ;
        RECT -252.285 -86.265 -252.115 -86.095 ;
        RECT -250.920 -86.265 -250.750 -86.095 ;
      LAYER met1 ;
        RECT -252.170 -86.000 -251.170 -85.300 ;
        RECT -252.350 -86.300 -250.660 -86.000 ;
    END
  END o_ranQ[184]
  PIN o_ranQ[185]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -257.435 -91.995 -256.930 -91.915 ;
        RECT -256.130 -91.995 -255.225 -91.905 ;
        RECT -257.435 -92.175 -255.225 -91.995 ;
      LAYER mcon ;
        RECT -257.245 -92.085 -257.075 -91.915 ;
        RECT -255.880 -92.085 -255.710 -91.915 ;
      LAYER met1 ;
        RECT -257.310 -92.180 -255.620 -91.880 ;
        RECT -257.130 -92.880 -256.130 -92.180 ;
    END
  END o_ranQ[185]
  PIN o_ranQ[186]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -262.395 -86.185 -260.185 -86.005 ;
        RECT -262.395 -86.265 -261.890 -86.185 ;
        RECT -261.090 -86.275 -260.185 -86.185 ;
      LAYER mcon ;
        RECT -262.205 -86.265 -262.035 -86.095 ;
        RECT -260.840 -86.265 -260.670 -86.095 ;
      LAYER met1 ;
        RECT -262.090 -86.000 -261.090 -85.300 ;
        RECT -262.270 -86.300 -260.580 -86.000 ;
    END
  END o_ranQ[186]
  PIN o_ranQ[187]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -267.355 -91.995 -266.850 -91.915 ;
        RECT -266.050 -91.995 -265.145 -91.905 ;
        RECT -267.355 -92.175 -265.145 -91.995 ;
      LAYER mcon ;
        RECT -267.165 -92.085 -266.995 -91.915 ;
        RECT -265.800 -92.085 -265.630 -91.915 ;
      LAYER met1 ;
        RECT -267.230 -92.180 -265.540 -91.880 ;
        RECT -267.050 -92.880 -266.050 -92.180 ;
    END
  END o_ranQ[187]
  PIN o_ranQ[189]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -277.275 -91.995 -276.770 -91.915 ;
        RECT -275.970 -91.995 -275.065 -91.905 ;
        RECT -277.275 -92.175 -275.065 -91.995 ;
      LAYER mcon ;
        RECT -277.085 -92.085 -276.915 -91.915 ;
        RECT -275.720 -92.085 -275.550 -91.915 ;
      LAYER met1 ;
        RECT -277.150 -92.180 -275.460 -91.880 ;
        RECT -276.970 -92.880 -275.970 -92.180 ;
    END
  END o_ranQ[189]
  PIN o_ranQ[190]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -282.235 -86.185 -280.025 -86.005 ;
        RECT -282.235 -86.265 -281.730 -86.185 ;
        RECT -280.930 -86.275 -280.025 -86.185 ;
      LAYER mcon ;
        RECT -282.045 -86.265 -281.875 -86.095 ;
        RECT -280.680 -86.265 -280.510 -86.095 ;
      LAYER met1 ;
        RECT -281.930 -86.000 -280.930 -85.300 ;
        RECT -282.110 -86.300 -280.420 -86.000 ;
    END
  END o_ranQ[190]
  PIN o_ranQ[191]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -287.195 -91.995 -286.690 -91.915 ;
        RECT -285.890 -91.995 -284.985 -91.905 ;
        RECT -287.195 -92.175 -284.985 -91.995 ;
      LAYER mcon ;
        RECT -287.005 -92.085 -286.835 -91.915 ;
        RECT -285.640 -92.085 -285.470 -91.915 ;
      LAYER met1 ;
        RECT -287.070 -92.180 -285.380 -91.880 ;
        RECT -286.890 -92.880 -285.890 -92.180 ;
    END
  END o_ranQ[191]
  PIN o_ranQ[252]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -272.065 -173.895 -269.855 -173.715 ;
        RECT -272.065 -173.975 -271.560 -173.895 ;
        RECT -270.760 -173.985 -269.855 -173.895 ;
      LAYER mcon ;
        RECT -271.875 -173.975 -271.705 -173.805 ;
        RECT -270.510 -173.975 -270.340 -173.805 ;
      LAYER met1 ;
        RECT -271.760 -173.710 -270.760 -173.010 ;
        RECT -271.940 -174.010 -270.250 -173.710 ;
    END
  END o_ranQ[252]
  PIN o_ranQ[193]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 20.575 -179.705 21.080 -179.625 ;
        RECT 21.880 -179.705 22.785 -179.615 ;
        RECT 20.575 -179.885 22.785 -179.705 ;
      LAYER mcon ;
        RECT 20.765 -179.795 20.935 -179.625 ;
        RECT 22.130 -179.795 22.300 -179.625 ;
      LAYER met1 ;
        RECT 20.700 -179.890 22.390 -179.590 ;
        RECT 20.880 -180.590 21.880 -179.890 ;
    END
  END o_ranQ[193]
  PIN o_ranQ[194]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 15.615 -173.895 17.825 -173.715 ;
        RECT 15.615 -173.975 16.120 -173.895 ;
        RECT 16.920 -173.985 17.825 -173.895 ;
      LAYER mcon ;
        RECT 15.805 -173.975 15.975 -173.805 ;
        RECT 17.170 -173.975 17.340 -173.805 ;
      LAYER met1 ;
        RECT 15.920 -173.710 16.920 -173.010 ;
        RECT 15.740 -174.010 17.430 -173.710 ;
    END
  END o_ranQ[194]
  PIN o_ranQ[195]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 10.655 -179.705 11.160 -179.625 ;
        RECT 11.960 -179.705 12.865 -179.615 ;
        RECT 10.655 -179.885 12.865 -179.705 ;
      LAYER mcon ;
        RECT 10.845 -179.795 11.015 -179.625 ;
        RECT 12.210 -179.795 12.380 -179.625 ;
      LAYER met1 ;
        RECT 10.780 -179.890 12.470 -179.590 ;
        RECT 10.960 -180.590 11.960 -179.890 ;
    END
  END o_ranQ[195]
  PIN o_ranQ[192]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 25.535 -173.895 27.745 -173.715 ;
        RECT 25.535 -173.975 26.040 -173.895 ;
        RECT 26.840 -173.985 27.745 -173.895 ;
      LAYER mcon ;
        RECT 25.725 -173.975 25.895 -173.805 ;
        RECT 27.090 -173.975 27.260 -173.805 ;
      LAYER met1 ;
        RECT 25.840 -173.710 26.840 -173.010 ;
        RECT 25.660 -174.010 27.350 -173.710 ;
    END
  END o_ranQ[192]
  PIN o_ranQ[196]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 5.695 -173.895 7.905 -173.715 ;
        RECT 5.695 -173.975 6.200 -173.895 ;
        RECT 7.000 -173.985 7.905 -173.895 ;
      LAYER mcon ;
        RECT 5.885 -173.975 6.055 -173.805 ;
        RECT 7.250 -173.975 7.420 -173.805 ;
      LAYER met1 ;
        RECT 6.000 -173.710 7.000 -173.010 ;
        RECT 5.820 -174.010 7.510 -173.710 ;
    END
  END o_ranQ[196]
  PIN o_ranQ[197]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 0.735 -179.705 1.240 -179.625 ;
        RECT 2.040 -179.705 2.945 -179.615 ;
        RECT 0.735 -179.885 2.945 -179.705 ;
      LAYER mcon ;
        RECT 0.925 -179.795 1.095 -179.625 ;
        RECT 2.290 -179.795 2.460 -179.625 ;
      LAYER met1 ;
        RECT 0.860 -179.890 2.550 -179.590 ;
        RECT 1.040 -180.590 2.040 -179.890 ;
    END
  END o_ranQ[197]
  PIN o_ranQ[198]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -4.225 -173.895 -2.015 -173.715 ;
        RECT -4.225 -173.975 -3.720 -173.895 ;
        RECT -2.920 -173.985 -2.015 -173.895 ;
      LAYER mcon ;
        RECT -4.035 -173.975 -3.865 -173.805 ;
        RECT -2.670 -173.975 -2.500 -173.805 ;
      LAYER met1 ;
        RECT -3.920 -173.710 -2.920 -173.010 ;
        RECT -4.100 -174.010 -2.410 -173.710 ;
    END
  END o_ranQ[198]
  PIN o_ranQ[199]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -9.185 -179.705 -8.680 -179.625 ;
        RECT -7.880 -179.705 -6.975 -179.615 ;
        RECT -9.185 -179.885 -6.975 -179.705 ;
      LAYER mcon ;
        RECT -8.995 -179.795 -8.825 -179.625 ;
        RECT -7.630 -179.795 -7.460 -179.625 ;
      LAYER met1 ;
        RECT -9.060 -179.890 -7.370 -179.590 ;
        RECT -8.880 -180.590 -7.880 -179.890 ;
    END
  END o_ranQ[199]
  PIN o_ranQ[200]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -14.145 -173.895 -11.935 -173.715 ;
        RECT -14.145 -173.975 -13.640 -173.895 ;
        RECT -12.840 -173.985 -11.935 -173.895 ;
      LAYER mcon ;
        RECT -13.955 -173.975 -13.785 -173.805 ;
        RECT -12.590 -173.975 -12.420 -173.805 ;
      LAYER met1 ;
        RECT -13.840 -173.710 -12.840 -173.010 ;
        RECT -14.020 -174.010 -12.330 -173.710 ;
    END
  END o_ranQ[200]
  PIN o_ranQ[201]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -19.105 -179.705 -18.600 -179.625 ;
        RECT -17.800 -179.705 -16.895 -179.615 ;
        RECT -19.105 -179.885 -16.895 -179.705 ;
      LAYER mcon ;
        RECT -18.915 -179.795 -18.745 -179.625 ;
        RECT -17.550 -179.795 -17.380 -179.625 ;
      LAYER met1 ;
        RECT -18.980 -179.890 -17.290 -179.590 ;
        RECT -18.800 -180.590 -17.800 -179.890 ;
    END
  END o_ranQ[201]
  PIN o_ranQ[202]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -24.065 -173.895 -21.855 -173.715 ;
        RECT -24.065 -173.975 -23.560 -173.895 ;
        RECT -22.760 -173.985 -21.855 -173.895 ;
      LAYER mcon ;
        RECT -23.875 -173.975 -23.705 -173.805 ;
        RECT -22.510 -173.975 -22.340 -173.805 ;
      LAYER met1 ;
        RECT -23.760 -173.710 -22.760 -173.010 ;
        RECT -23.940 -174.010 -22.250 -173.710 ;
    END
  END o_ranQ[202]
  PIN o_ranQ[203]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -29.025 -179.705 -28.520 -179.625 ;
        RECT -27.720 -179.705 -26.815 -179.615 ;
        RECT -29.025 -179.885 -26.815 -179.705 ;
      LAYER mcon ;
        RECT -28.835 -179.795 -28.665 -179.625 ;
        RECT -27.470 -179.795 -27.300 -179.625 ;
      LAYER met1 ;
        RECT -28.900 -179.890 -27.210 -179.590 ;
        RECT -28.720 -180.590 -27.720 -179.890 ;
    END
  END o_ranQ[203]
  PIN o_ranQ[204]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -33.985 -173.895 -31.775 -173.715 ;
        RECT -33.985 -173.975 -33.480 -173.895 ;
        RECT -32.680 -173.985 -31.775 -173.895 ;
      LAYER mcon ;
        RECT -33.795 -173.975 -33.625 -173.805 ;
        RECT -32.430 -173.975 -32.260 -173.805 ;
      LAYER met1 ;
        RECT -33.680 -173.710 -32.680 -173.010 ;
        RECT -33.860 -174.010 -32.170 -173.710 ;
    END
  END o_ranQ[204]
  PIN o_ranQ[205]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -38.945 -179.705 -38.440 -179.625 ;
        RECT -37.640 -179.705 -36.735 -179.615 ;
        RECT -38.945 -179.885 -36.735 -179.705 ;
      LAYER mcon ;
        RECT -38.755 -179.795 -38.585 -179.625 ;
        RECT -37.390 -179.795 -37.220 -179.625 ;
      LAYER met1 ;
        RECT -38.820 -179.890 -37.130 -179.590 ;
        RECT -38.640 -180.590 -37.640 -179.890 ;
    END
  END o_ranQ[205]
  PIN o_ranQ[206]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -43.905 -173.895 -41.695 -173.715 ;
        RECT -43.905 -173.975 -43.400 -173.895 ;
        RECT -42.600 -173.985 -41.695 -173.895 ;
      LAYER mcon ;
        RECT -43.715 -173.975 -43.545 -173.805 ;
        RECT -42.350 -173.975 -42.180 -173.805 ;
      LAYER met1 ;
        RECT -43.600 -173.710 -42.600 -173.010 ;
        RECT -43.780 -174.010 -42.090 -173.710 ;
    END
  END o_ranQ[206]
  PIN o_ranQ[207]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -48.865 -179.705 -48.360 -179.625 ;
        RECT -47.560 -179.705 -46.655 -179.615 ;
        RECT -48.865 -179.885 -46.655 -179.705 ;
      LAYER mcon ;
        RECT -48.675 -179.795 -48.505 -179.625 ;
        RECT -47.310 -179.795 -47.140 -179.625 ;
      LAYER met1 ;
        RECT -48.740 -179.890 -47.050 -179.590 ;
        RECT -48.560 -180.590 -47.560 -179.890 ;
    END
  END o_ranQ[207]
  PIN o_ranQ[209]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -58.785 -179.705 -58.280 -179.625 ;
        RECT -57.480 -179.705 -56.575 -179.615 ;
        RECT -58.785 -179.885 -56.575 -179.705 ;
      LAYER mcon ;
        RECT -58.595 -179.795 -58.425 -179.625 ;
        RECT -57.230 -179.795 -57.060 -179.625 ;
      LAYER met1 ;
        RECT -58.660 -179.890 -56.970 -179.590 ;
        RECT -58.480 -180.590 -57.480 -179.890 ;
    END
  END o_ranQ[209]
  PIN o_ranQ[210]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -63.745 -173.895 -61.535 -173.715 ;
        RECT -63.745 -173.975 -63.240 -173.895 ;
        RECT -62.440 -173.985 -61.535 -173.895 ;
      LAYER mcon ;
        RECT -63.555 -173.975 -63.385 -173.805 ;
        RECT -62.190 -173.975 -62.020 -173.805 ;
      LAYER met1 ;
        RECT -63.440 -173.710 -62.440 -173.010 ;
        RECT -63.620 -174.010 -61.930 -173.710 ;
    END
  END o_ranQ[210]
  PIN o_ranQ[211]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -68.705 -179.705 -68.200 -179.625 ;
        RECT -67.400 -179.705 -66.495 -179.615 ;
        RECT -68.705 -179.885 -66.495 -179.705 ;
      LAYER mcon ;
        RECT -68.515 -179.795 -68.345 -179.625 ;
        RECT -67.150 -179.795 -66.980 -179.625 ;
      LAYER met1 ;
        RECT -68.580 -179.890 -66.890 -179.590 ;
        RECT -68.400 -180.590 -67.400 -179.890 ;
    END
  END o_ranQ[211]
  PIN o_ranQ[208]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -53.825 -173.895 -51.615 -173.715 ;
        RECT -53.825 -173.975 -53.320 -173.895 ;
        RECT -52.520 -173.985 -51.615 -173.895 ;
      LAYER mcon ;
        RECT -53.635 -173.975 -53.465 -173.805 ;
        RECT -52.270 -173.975 -52.100 -173.805 ;
      LAYER met1 ;
        RECT -53.520 -173.710 -52.520 -173.010 ;
        RECT -53.700 -174.010 -52.010 -173.710 ;
    END
  END o_ranQ[208]
  PIN o_ranQ[212]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -73.665 -173.895 -71.455 -173.715 ;
        RECT -73.665 -173.975 -73.160 -173.895 ;
        RECT -72.360 -173.985 -71.455 -173.895 ;
      LAYER mcon ;
        RECT -73.475 -173.975 -73.305 -173.805 ;
        RECT -72.110 -173.975 -71.940 -173.805 ;
      LAYER met1 ;
        RECT -73.360 -173.710 -72.360 -173.010 ;
        RECT -73.540 -174.010 -71.850 -173.710 ;
    END
  END o_ranQ[212]
  PIN o_ranQ[213]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -78.625 -179.705 -78.120 -179.625 ;
        RECT -77.320 -179.705 -76.415 -179.615 ;
        RECT -78.625 -179.885 -76.415 -179.705 ;
      LAYER mcon ;
        RECT -78.435 -179.795 -78.265 -179.625 ;
        RECT -77.070 -179.795 -76.900 -179.625 ;
      LAYER met1 ;
        RECT -78.500 -179.890 -76.810 -179.590 ;
        RECT -78.320 -180.590 -77.320 -179.890 ;
    END
  END o_ranQ[213]
  PIN o_ranQ[214]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -83.585 -173.895 -81.375 -173.715 ;
        RECT -83.585 -173.975 -83.080 -173.895 ;
        RECT -82.280 -173.985 -81.375 -173.895 ;
      LAYER mcon ;
        RECT -83.395 -173.975 -83.225 -173.805 ;
        RECT -82.030 -173.975 -81.860 -173.805 ;
      LAYER met1 ;
        RECT -83.280 -173.710 -82.280 -173.010 ;
        RECT -83.460 -174.010 -81.770 -173.710 ;
    END
  END o_ranQ[214]
  PIN o_ranQ[215]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -88.545 -179.705 -88.040 -179.625 ;
        RECT -87.240 -179.705 -86.335 -179.615 ;
        RECT -88.545 -179.885 -86.335 -179.705 ;
      LAYER mcon ;
        RECT -88.355 -179.795 -88.185 -179.625 ;
        RECT -86.990 -179.795 -86.820 -179.625 ;
      LAYER met1 ;
        RECT -88.420 -179.890 -86.730 -179.590 ;
        RECT -88.240 -180.590 -87.240 -179.890 ;
    END
  END o_ranQ[215]
  PIN o_ranQ[216]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -93.505 -173.895 -91.295 -173.715 ;
        RECT -93.505 -173.975 -93.000 -173.895 ;
        RECT -92.200 -173.985 -91.295 -173.895 ;
      LAYER mcon ;
        RECT -93.315 -173.975 -93.145 -173.805 ;
        RECT -91.950 -173.975 -91.780 -173.805 ;
      LAYER met1 ;
        RECT -93.200 -173.710 -92.200 -173.010 ;
        RECT -93.380 -174.010 -91.690 -173.710 ;
    END
  END o_ranQ[216]
  PIN o_ranQ[217]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -98.465 -179.705 -97.960 -179.625 ;
        RECT -97.160 -179.705 -96.255 -179.615 ;
        RECT -98.465 -179.885 -96.255 -179.705 ;
      LAYER mcon ;
        RECT -98.275 -179.795 -98.105 -179.625 ;
        RECT -96.910 -179.795 -96.740 -179.625 ;
      LAYER met1 ;
        RECT -98.340 -179.890 -96.650 -179.590 ;
        RECT -98.160 -180.590 -97.160 -179.890 ;
    END
  END o_ranQ[217]
  PIN o_ranQ[218]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -103.425 -173.895 -101.215 -173.715 ;
        RECT -103.425 -173.975 -102.920 -173.895 ;
        RECT -102.120 -173.985 -101.215 -173.895 ;
      LAYER mcon ;
        RECT -103.235 -173.975 -103.065 -173.805 ;
        RECT -101.870 -173.975 -101.700 -173.805 ;
      LAYER met1 ;
        RECT -103.120 -173.710 -102.120 -173.010 ;
        RECT -103.300 -174.010 -101.610 -173.710 ;
    END
  END o_ranQ[218]
  PIN o_ranQ[219]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -108.385 -179.705 -107.880 -179.625 ;
        RECT -107.080 -179.705 -106.175 -179.615 ;
        RECT -108.385 -179.885 -106.175 -179.705 ;
      LAYER mcon ;
        RECT -108.195 -179.795 -108.025 -179.625 ;
        RECT -106.830 -179.795 -106.660 -179.625 ;
      LAYER met1 ;
        RECT -108.260 -179.890 -106.570 -179.590 ;
        RECT -108.080 -180.590 -107.080 -179.890 ;
    END
  END o_ranQ[219]
  PIN o_ranQ[220]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -113.345 -173.895 -111.135 -173.715 ;
        RECT -113.345 -173.975 -112.840 -173.895 ;
        RECT -112.040 -173.985 -111.135 -173.895 ;
      LAYER mcon ;
        RECT -113.155 -173.975 -112.985 -173.805 ;
        RECT -111.790 -173.975 -111.620 -173.805 ;
      LAYER met1 ;
        RECT -113.040 -173.710 -112.040 -173.010 ;
        RECT -113.220 -174.010 -111.530 -173.710 ;
    END
  END o_ranQ[220]
  PIN o_ranQ[221]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -118.305 -179.705 -117.800 -179.625 ;
        RECT -117.000 -179.705 -116.095 -179.615 ;
        RECT -118.305 -179.885 -116.095 -179.705 ;
      LAYER mcon ;
        RECT -118.115 -179.795 -117.945 -179.625 ;
        RECT -116.750 -179.795 -116.580 -179.625 ;
      LAYER met1 ;
        RECT -118.180 -179.890 -116.490 -179.590 ;
        RECT -118.000 -180.590 -117.000 -179.890 ;
    END
  END o_ranQ[221]
  PIN o_ranQ[222]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -123.265 -173.895 -121.055 -173.715 ;
        RECT -123.265 -173.975 -122.760 -173.895 ;
        RECT -121.960 -173.985 -121.055 -173.895 ;
      LAYER mcon ;
        RECT -123.075 -173.975 -122.905 -173.805 ;
        RECT -121.710 -173.975 -121.540 -173.805 ;
      LAYER met1 ;
        RECT -122.960 -173.710 -121.960 -173.010 ;
        RECT -123.140 -174.010 -121.450 -173.710 ;
    END
  END o_ranQ[222]
  PIN o_ranQ[223]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -128.225 -179.705 -127.720 -179.625 ;
        RECT -126.920 -179.705 -126.015 -179.615 ;
        RECT -128.225 -179.885 -126.015 -179.705 ;
      LAYER mcon ;
        RECT -128.035 -179.795 -127.865 -179.625 ;
        RECT -126.670 -179.795 -126.500 -179.625 ;
      LAYER met1 ;
        RECT -128.100 -179.890 -126.410 -179.590 ;
        RECT -127.920 -180.590 -126.920 -179.890 ;
    END
  END o_ranQ[223]
  PIN o_ranQ[225]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -138.145 -179.705 -137.640 -179.625 ;
        RECT -136.840 -179.705 -135.935 -179.615 ;
        RECT -138.145 -179.885 -135.935 -179.705 ;
      LAYER mcon ;
        RECT -137.955 -179.795 -137.785 -179.625 ;
        RECT -136.590 -179.795 -136.420 -179.625 ;
      LAYER met1 ;
        RECT -138.020 -179.890 -136.330 -179.590 ;
        RECT -137.840 -180.590 -136.840 -179.890 ;
    END
  END o_ranQ[225]
  PIN o_ranQ[226]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -143.105 -173.895 -140.895 -173.715 ;
        RECT -143.105 -173.975 -142.600 -173.895 ;
        RECT -141.800 -173.985 -140.895 -173.895 ;
      LAYER mcon ;
        RECT -142.915 -173.975 -142.745 -173.805 ;
        RECT -141.550 -173.975 -141.380 -173.805 ;
      LAYER met1 ;
        RECT -142.800 -173.710 -141.800 -173.010 ;
        RECT -142.980 -174.010 -141.290 -173.710 ;
    END
  END o_ranQ[226]
  PIN o_ranQ[227]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -148.065 -179.705 -147.560 -179.625 ;
        RECT -146.760 -179.705 -145.855 -179.615 ;
        RECT -148.065 -179.885 -145.855 -179.705 ;
      LAYER mcon ;
        RECT -147.875 -179.795 -147.705 -179.625 ;
        RECT -146.510 -179.795 -146.340 -179.625 ;
      LAYER met1 ;
        RECT -147.940 -179.890 -146.250 -179.590 ;
        RECT -147.760 -180.590 -146.760 -179.890 ;
    END
  END o_ranQ[227]
  PIN o_ranQ[224]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -133.185 -173.895 -130.975 -173.715 ;
        RECT -133.185 -173.975 -132.680 -173.895 ;
        RECT -131.880 -173.985 -130.975 -173.895 ;
      LAYER mcon ;
        RECT -132.995 -173.975 -132.825 -173.805 ;
        RECT -131.630 -173.975 -131.460 -173.805 ;
      LAYER met1 ;
        RECT -132.880 -173.710 -131.880 -173.010 ;
        RECT -133.060 -174.010 -131.370 -173.710 ;
    END
  END o_ranQ[224]
  PIN o_ranQ[228]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -153.025 -173.895 -150.815 -173.715 ;
        RECT -153.025 -173.975 -152.520 -173.895 ;
        RECT -151.720 -173.985 -150.815 -173.895 ;
      LAYER mcon ;
        RECT -152.835 -173.975 -152.665 -173.805 ;
        RECT -151.470 -173.975 -151.300 -173.805 ;
      LAYER met1 ;
        RECT -152.720 -173.710 -151.720 -173.010 ;
        RECT -152.900 -174.010 -151.210 -173.710 ;
    END
  END o_ranQ[228]
  PIN o_ranQ[229]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -157.985 -179.705 -157.480 -179.625 ;
        RECT -156.680 -179.705 -155.775 -179.615 ;
        RECT -157.985 -179.885 -155.775 -179.705 ;
      LAYER mcon ;
        RECT -157.795 -179.795 -157.625 -179.625 ;
        RECT -156.430 -179.795 -156.260 -179.625 ;
      LAYER met1 ;
        RECT -157.860 -179.890 -156.170 -179.590 ;
        RECT -157.680 -180.590 -156.680 -179.890 ;
    END
  END o_ranQ[229]
  PIN o_ranQ[230]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -162.945 -173.895 -160.735 -173.715 ;
        RECT -162.945 -173.975 -162.440 -173.895 ;
        RECT -161.640 -173.985 -160.735 -173.895 ;
      LAYER mcon ;
        RECT -162.755 -173.975 -162.585 -173.805 ;
        RECT -161.390 -173.975 -161.220 -173.805 ;
      LAYER met1 ;
        RECT -162.640 -173.710 -161.640 -173.010 ;
        RECT -162.820 -174.010 -161.130 -173.710 ;
    END
  END o_ranQ[230]
  PIN o_ranQ[231]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -167.905 -179.705 -167.400 -179.625 ;
        RECT -166.600 -179.705 -165.695 -179.615 ;
        RECT -167.905 -179.885 -165.695 -179.705 ;
      LAYER mcon ;
        RECT -167.715 -179.795 -167.545 -179.625 ;
        RECT -166.350 -179.795 -166.180 -179.625 ;
      LAYER met1 ;
        RECT -167.780 -179.890 -166.090 -179.590 ;
        RECT -167.600 -180.590 -166.600 -179.890 ;
    END
  END o_ranQ[231]
  PIN o_ranQ[232]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -172.865 -173.895 -170.655 -173.715 ;
        RECT -172.865 -173.975 -172.360 -173.895 ;
        RECT -171.560 -173.985 -170.655 -173.895 ;
      LAYER mcon ;
        RECT -172.675 -173.975 -172.505 -173.805 ;
        RECT -171.310 -173.975 -171.140 -173.805 ;
      LAYER met1 ;
        RECT -172.560 -173.710 -171.560 -173.010 ;
        RECT -172.740 -174.010 -171.050 -173.710 ;
    END
  END o_ranQ[232]
  PIN o_ranQ[233]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -177.825 -179.705 -177.320 -179.625 ;
        RECT -176.520 -179.705 -175.615 -179.615 ;
        RECT -177.825 -179.885 -175.615 -179.705 ;
      LAYER mcon ;
        RECT -177.635 -179.795 -177.465 -179.625 ;
        RECT -176.270 -179.795 -176.100 -179.625 ;
      LAYER met1 ;
        RECT -177.700 -179.890 -176.010 -179.590 ;
        RECT -177.520 -180.590 -176.520 -179.890 ;
    END
  END o_ranQ[233]
  PIN o_ranQ[234]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -182.785 -173.895 -180.575 -173.715 ;
        RECT -182.785 -173.975 -182.280 -173.895 ;
        RECT -181.480 -173.985 -180.575 -173.895 ;
      LAYER mcon ;
        RECT -182.595 -173.975 -182.425 -173.805 ;
        RECT -181.230 -173.975 -181.060 -173.805 ;
      LAYER met1 ;
        RECT -182.480 -173.710 -181.480 -173.010 ;
        RECT -182.660 -174.010 -180.970 -173.710 ;
    END
  END o_ranQ[234]
  PIN o_ranQ[235]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -187.745 -179.705 -187.240 -179.625 ;
        RECT -186.440 -179.705 -185.535 -179.615 ;
        RECT -187.745 -179.885 -185.535 -179.705 ;
      LAYER mcon ;
        RECT -187.555 -179.795 -187.385 -179.625 ;
        RECT -186.190 -179.795 -186.020 -179.625 ;
      LAYER met1 ;
        RECT -187.620 -179.890 -185.930 -179.590 ;
        RECT -187.440 -180.590 -186.440 -179.890 ;
    END
  END o_ranQ[235]
  PIN o_ranQ[236]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -192.705 -173.895 -190.495 -173.715 ;
        RECT -192.705 -173.975 -192.200 -173.895 ;
        RECT -191.400 -173.985 -190.495 -173.895 ;
      LAYER mcon ;
        RECT -192.515 -173.975 -192.345 -173.805 ;
        RECT -191.150 -173.975 -190.980 -173.805 ;
      LAYER met1 ;
        RECT -192.400 -173.710 -191.400 -173.010 ;
        RECT -192.580 -174.010 -190.890 -173.710 ;
    END
  END o_ranQ[236]
  PIN o_ranQ[237]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -197.665 -179.705 -197.160 -179.625 ;
        RECT -196.360 -179.705 -195.455 -179.615 ;
        RECT -197.665 -179.885 -195.455 -179.705 ;
      LAYER mcon ;
        RECT -197.475 -179.795 -197.305 -179.625 ;
        RECT -196.110 -179.795 -195.940 -179.625 ;
      LAYER met1 ;
        RECT -197.540 -179.890 -195.850 -179.590 ;
        RECT -197.360 -180.590 -196.360 -179.890 ;
    END
  END o_ranQ[237]
  PIN o_ranQ[238]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -202.625 -173.895 -200.415 -173.715 ;
        RECT -202.625 -173.975 -202.120 -173.895 ;
        RECT -201.320 -173.985 -200.415 -173.895 ;
      LAYER mcon ;
        RECT -202.435 -173.975 -202.265 -173.805 ;
        RECT -201.070 -173.975 -200.900 -173.805 ;
      LAYER met1 ;
        RECT -202.320 -173.710 -201.320 -173.010 ;
        RECT -202.500 -174.010 -200.810 -173.710 ;
    END
  END o_ranQ[238]
  PIN o_ranQ[239]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -207.585 -179.705 -207.080 -179.625 ;
        RECT -206.280 -179.705 -205.375 -179.615 ;
        RECT -207.585 -179.885 -205.375 -179.705 ;
      LAYER mcon ;
        RECT -207.395 -179.795 -207.225 -179.625 ;
        RECT -206.030 -179.795 -205.860 -179.625 ;
      LAYER met1 ;
        RECT -207.460 -179.890 -205.770 -179.590 ;
        RECT -207.280 -180.590 -206.280 -179.890 ;
    END
  END o_ranQ[239]
  PIN o_ranQ[241]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -217.505 -179.705 -217.000 -179.625 ;
        RECT -216.200 -179.705 -215.295 -179.615 ;
        RECT -217.505 -179.885 -215.295 -179.705 ;
      LAYER mcon ;
        RECT -217.315 -179.795 -217.145 -179.625 ;
        RECT -215.950 -179.795 -215.780 -179.625 ;
      LAYER met1 ;
        RECT -217.380 -179.890 -215.690 -179.590 ;
        RECT -217.200 -180.590 -216.200 -179.890 ;
    END
  END o_ranQ[241]
  PIN o_ranQ[242]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -222.465 -173.895 -220.255 -173.715 ;
        RECT -222.465 -173.975 -221.960 -173.895 ;
        RECT -221.160 -173.985 -220.255 -173.895 ;
      LAYER mcon ;
        RECT -222.275 -173.975 -222.105 -173.805 ;
        RECT -220.910 -173.975 -220.740 -173.805 ;
      LAYER met1 ;
        RECT -222.160 -173.710 -221.160 -173.010 ;
        RECT -222.340 -174.010 -220.650 -173.710 ;
    END
  END o_ranQ[242]
  PIN o_ranQ[243]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -227.425 -179.705 -226.920 -179.625 ;
        RECT -226.120 -179.705 -225.215 -179.615 ;
        RECT -227.425 -179.885 -225.215 -179.705 ;
      LAYER mcon ;
        RECT -227.235 -179.795 -227.065 -179.625 ;
        RECT -225.870 -179.795 -225.700 -179.625 ;
      LAYER met1 ;
        RECT -227.300 -179.890 -225.610 -179.590 ;
        RECT -227.120 -180.590 -226.120 -179.890 ;
    END
  END o_ranQ[243]
  PIN o_ranQ[240]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -212.545 -173.895 -210.335 -173.715 ;
        RECT -212.545 -173.975 -212.040 -173.895 ;
        RECT -211.240 -173.985 -210.335 -173.895 ;
      LAYER mcon ;
        RECT -212.355 -173.975 -212.185 -173.805 ;
        RECT -210.990 -173.975 -210.820 -173.805 ;
      LAYER met1 ;
        RECT -212.240 -173.710 -211.240 -173.010 ;
        RECT -212.420 -174.010 -210.730 -173.710 ;
    END
  END o_ranQ[240]
  PIN o_ranQ[244]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -232.385 -173.895 -230.175 -173.715 ;
        RECT -232.385 -173.975 -231.880 -173.895 ;
        RECT -231.080 -173.985 -230.175 -173.895 ;
      LAYER mcon ;
        RECT -232.195 -173.975 -232.025 -173.805 ;
        RECT -230.830 -173.975 -230.660 -173.805 ;
      LAYER met1 ;
        RECT -232.080 -173.710 -231.080 -173.010 ;
        RECT -232.260 -174.010 -230.570 -173.710 ;
    END
  END o_ranQ[244]
  PIN o_ranQ[245]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -237.345 -179.705 -236.840 -179.625 ;
        RECT -236.040 -179.705 -235.135 -179.615 ;
        RECT -237.345 -179.885 -235.135 -179.705 ;
      LAYER mcon ;
        RECT -237.155 -179.795 -236.985 -179.625 ;
        RECT -235.790 -179.795 -235.620 -179.625 ;
      LAYER met1 ;
        RECT -237.220 -179.890 -235.530 -179.590 ;
        RECT -237.040 -180.590 -236.040 -179.890 ;
    END
  END o_ranQ[245]
  PIN o_ranQ[246]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -242.305 -173.895 -240.095 -173.715 ;
        RECT -242.305 -173.975 -241.800 -173.895 ;
        RECT -241.000 -173.985 -240.095 -173.895 ;
      LAYER mcon ;
        RECT -242.115 -173.975 -241.945 -173.805 ;
        RECT -240.750 -173.975 -240.580 -173.805 ;
      LAYER met1 ;
        RECT -242.000 -173.710 -241.000 -173.010 ;
        RECT -242.180 -174.010 -240.490 -173.710 ;
    END
  END o_ranQ[246]
  PIN o_ranQ[247]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -247.265 -179.705 -246.760 -179.625 ;
        RECT -245.960 -179.705 -245.055 -179.615 ;
        RECT -247.265 -179.885 -245.055 -179.705 ;
      LAYER mcon ;
        RECT -247.075 -179.795 -246.905 -179.625 ;
        RECT -245.710 -179.795 -245.540 -179.625 ;
      LAYER met1 ;
        RECT -247.140 -179.890 -245.450 -179.590 ;
        RECT -246.960 -180.590 -245.960 -179.890 ;
    END
  END o_ranQ[247]
  PIN o_ranQ[248]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -252.225 -173.895 -250.015 -173.715 ;
        RECT -252.225 -173.975 -251.720 -173.895 ;
        RECT -250.920 -173.985 -250.015 -173.895 ;
      LAYER mcon ;
        RECT -252.035 -173.975 -251.865 -173.805 ;
        RECT -250.670 -173.975 -250.500 -173.805 ;
      LAYER met1 ;
        RECT -251.920 -173.710 -250.920 -173.010 ;
        RECT -252.100 -174.010 -250.410 -173.710 ;
    END
  END o_ranQ[248]
  PIN o_ranQ[249]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -257.185 -179.705 -256.680 -179.625 ;
        RECT -255.880 -179.705 -254.975 -179.615 ;
        RECT -257.185 -179.885 -254.975 -179.705 ;
      LAYER mcon ;
        RECT -256.995 -179.795 -256.825 -179.625 ;
        RECT -255.630 -179.795 -255.460 -179.625 ;
      LAYER met1 ;
        RECT -257.060 -179.890 -255.370 -179.590 ;
        RECT -256.880 -180.590 -255.880 -179.890 ;
    END
  END o_ranQ[249]
  PIN o_ranQ[250]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -262.145 -173.895 -259.935 -173.715 ;
        RECT -262.145 -173.975 -261.640 -173.895 ;
        RECT -260.840 -173.985 -259.935 -173.895 ;
      LAYER mcon ;
        RECT -261.955 -173.975 -261.785 -173.805 ;
        RECT -260.590 -173.975 -260.420 -173.805 ;
      LAYER met1 ;
        RECT -261.840 -173.710 -260.840 -173.010 ;
        RECT -262.020 -174.010 -260.330 -173.710 ;
    END
  END o_ranQ[250]
  PIN o_ranQ[251]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -267.105 -179.705 -266.600 -179.625 ;
        RECT -265.800 -179.705 -264.895 -179.615 ;
        RECT -267.105 -179.885 -264.895 -179.705 ;
      LAYER mcon ;
        RECT -266.915 -179.795 -266.745 -179.625 ;
        RECT -265.550 -179.795 -265.380 -179.625 ;
      LAYER met1 ;
        RECT -266.980 -179.890 -265.290 -179.590 ;
        RECT -266.800 -180.590 -265.800 -179.890 ;
    END
  END o_ranQ[251]
  PIN o_ranQ[253]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -277.025 -179.705 -276.520 -179.625 ;
        RECT -275.720 -179.705 -274.815 -179.615 ;
        RECT -277.025 -179.885 -274.815 -179.705 ;
      LAYER mcon ;
        RECT -276.835 -179.795 -276.665 -179.625 ;
        RECT -275.470 -179.795 -275.300 -179.625 ;
      LAYER met1 ;
        RECT -276.900 -179.890 -275.210 -179.590 ;
        RECT -276.720 -180.590 -275.720 -179.890 ;
    END
  END o_ranQ[253]
  PIN o_ranQ[254]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -281.985 -173.895 -279.775 -173.715 ;
        RECT -281.985 -173.975 -281.480 -173.895 ;
        RECT -280.680 -173.985 -279.775 -173.895 ;
      LAYER mcon ;
        RECT -281.795 -173.975 -281.625 -173.805 ;
        RECT -280.430 -173.975 -280.260 -173.805 ;
      LAYER met1 ;
        RECT -281.680 -173.710 -280.680 -173.010 ;
        RECT -281.860 -174.010 -280.170 -173.710 ;
    END
  END o_ranQ[254]
  PIN o_ranQ[255]
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -286.945 -179.705 -286.440 -179.625 ;
        RECT -285.640 -179.705 -284.735 -179.615 ;
        RECT -286.945 -179.885 -284.735 -179.705 ;
      LAYER mcon ;
        RECT -286.755 -179.795 -286.585 -179.625 ;
        RECT -285.390 -179.795 -285.220 -179.625 ;
      LAYER met1 ;
        RECT -286.820 -179.890 -285.130 -179.590 ;
        RECT -286.640 -180.590 -285.640 -179.890 ;
    END
  END o_ranQ[255]
  OBS
      LAYER nwell ;
        RECT -290.950 95.095 -289.345 95.330 ;
        RECT -291.650 93.570 -289.345 95.095 ;
      LAYER pwell ;
        RECT -288.925 93.765 -288.145 95.135 ;
        RECT -284.395 93.765 -283.615 95.135 ;
        RECT -279.005 93.765 -278.225 95.135 ;
        RECT -274.475 93.765 -273.695 95.135 ;
        RECT -269.085 93.765 -268.305 95.135 ;
        RECT -264.555 93.765 -263.775 95.135 ;
        RECT -259.165 93.765 -258.385 95.135 ;
        RECT -254.635 93.765 -253.855 95.135 ;
        RECT -249.245 93.765 -248.465 95.135 ;
        RECT -244.715 93.765 -243.935 95.135 ;
        RECT -239.325 93.765 -238.545 95.135 ;
        RECT -234.795 93.765 -234.015 95.135 ;
        RECT -229.405 93.765 -228.625 95.135 ;
        RECT -224.875 93.765 -224.095 95.135 ;
        RECT -219.485 93.765 -218.705 95.135 ;
        RECT -214.955 93.765 -214.175 95.135 ;
        RECT -209.565 93.765 -208.785 95.135 ;
        RECT -205.035 93.765 -204.255 95.135 ;
        RECT -199.645 93.765 -198.865 95.135 ;
        RECT -195.115 93.765 -194.335 95.135 ;
        RECT -189.725 93.765 -188.945 95.135 ;
        RECT -185.195 93.765 -184.415 95.135 ;
        RECT -179.805 93.765 -179.025 95.135 ;
        RECT -175.275 93.765 -174.495 95.135 ;
        RECT -169.885 93.765 -169.105 95.135 ;
        RECT -165.355 93.765 -164.575 95.135 ;
        RECT -159.965 93.765 -159.185 95.135 ;
        RECT -155.435 93.765 -154.655 95.135 ;
        RECT -150.045 93.765 -149.265 95.135 ;
        RECT -145.515 93.765 -144.735 95.135 ;
        RECT -140.125 93.765 -139.345 95.135 ;
        RECT -135.595 93.765 -134.815 95.135 ;
        RECT -130.205 93.765 -129.425 95.135 ;
        RECT -125.675 93.765 -124.895 95.135 ;
        RECT -120.285 93.765 -119.505 95.135 ;
        RECT -115.755 93.765 -114.975 95.135 ;
        RECT -110.365 93.765 -109.585 95.135 ;
        RECT -105.835 93.765 -105.055 95.135 ;
        RECT -100.445 93.765 -99.665 95.135 ;
        RECT -95.915 93.765 -95.135 95.135 ;
        RECT -90.525 93.765 -89.745 95.135 ;
        RECT -85.995 93.765 -85.215 95.135 ;
        RECT -80.605 93.765 -79.825 95.135 ;
        RECT -76.075 93.765 -75.295 95.135 ;
        RECT -70.685 93.765 -69.905 95.135 ;
        RECT -66.155 93.765 -65.375 95.135 ;
        RECT -60.765 93.765 -59.985 95.135 ;
        RECT -56.235 93.765 -55.455 95.135 ;
        RECT -50.845 93.765 -50.065 95.135 ;
        RECT -46.315 93.765 -45.535 95.135 ;
        RECT -40.925 93.765 -40.145 95.135 ;
        RECT -36.395 93.765 -35.615 95.135 ;
        RECT -31.005 93.765 -30.225 95.135 ;
        RECT -26.475 93.765 -25.695 95.135 ;
        RECT -21.085 93.765 -20.305 95.135 ;
        RECT -16.555 93.765 -15.775 95.135 ;
        RECT -11.165 93.765 -10.385 95.135 ;
        RECT -6.635 93.765 -5.855 95.135 ;
        RECT -1.245 93.765 -0.465 95.135 ;
        RECT 3.285 93.765 4.065 95.135 ;
        RECT 8.675 93.765 9.455 95.135 ;
        RECT 13.205 93.765 13.985 95.135 ;
        RECT 18.595 93.765 19.375 95.135 ;
        RECT 23.125 93.765 23.905 95.135 ;
      LAYER nwell ;
        RECT -291.650 93.510 -290.810 93.570 ;
      LAYER pwell ;
        RECT -290.975 93.140 -289.625 93.225 ;
        RECT -291.445 92.355 -289.625 93.140 ;
        RECT -290.975 92.315 -289.625 92.355 ;
        RECT 24.605 93.140 25.955 93.225 ;
        RECT 24.605 92.355 26.425 93.140 ;
        RECT 24.605 92.315 25.955 92.355 ;
      LAYER nwell ;
        RECT -291.650 90.420 -289.430 92.025 ;
      LAYER pwell ;
        RECT -289.355 90.015 -288.575 90.175 ;
        RECT -290.145 89.230 -288.575 90.015 ;
        RECT -289.355 88.805 -288.575 89.230 ;
        RECT -283.965 88.805 -283.185 90.175 ;
        RECT -279.435 88.805 -278.655 90.175 ;
        RECT -274.045 88.805 -273.265 90.175 ;
        RECT -269.515 88.805 -268.735 90.175 ;
        RECT -264.125 88.805 -263.345 90.175 ;
        RECT -259.595 88.805 -258.815 90.175 ;
        RECT -254.205 88.805 -253.425 90.175 ;
        RECT -249.675 88.805 -248.895 90.175 ;
        RECT -244.285 88.805 -243.505 90.175 ;
        RECT -239.755 88.805 -238.975 90.175 ;
        RECT -234.365 88.805 -233.585 90.175 ;
        RECT -229.835 88.805 -229.055 90.175 ;
        RECT -224.445 88.805 -223.665 90.175 ;
        RECT -219.915 88.805 -219.135 90.175 ;
        RECT -214.525 88.805 -213.745 90.175 ;
        RECT -209.995 88.805 -209.215 90.175 ;
        RECT -204.605 88.805 -203.825 90.175 ;
        RECT -200.075 88.805 -199.295 90.175 ;
        RECT -194.685 88.805 -193.905 90.175 ;
        RECT -190.155 88.805 -189.375 90.175 ;
        RECT -184.765 88.805 -183.985 90.175 ;
        RECT -180.235 88.805 -179.455 90.175 ;
        RECT -174.845 88.805 -174.065 90.175 ;
        RECT -170.315 88.805 -169.535 90.175 ;
        RECT -164.925 88.805 -164.145 90.175 ;
        RECT -160.395 88.805 -159.615 90.175 ;
        RECT -155.005 88.805 -154.225 90.175 ;
        RECT -150.475 88.805 -149.695 90.175 ;
        RECT -145.085 88.805 -144.305 90.175 ;
        RECT -140.555 88.805 -139.775 90.175 ;
        RECT -135.165 88.805 -134.385 90.175 ;
        RECT -130.635 88.805 -129.855 90.175 ;
        RECT -125.245 88.805 -124.465 90.175 ;
        RECT -120.715 88.805 -119.935 90.175 ;
        RECT -115.325 88.805 -114.545 90.175 ;
        RECT -110.795 88.805 -110.015 90.175 ;
        RECT -105.405 88.805 -104.625 90.175 ;
        RECT -100.875 88.805 -100.095 90.175 ;
        RECT -95.485 88.805 -94.705 90.175 ;
        RECT -90.955 88.805 -90.175 90.175 ;
        RECT -85.565 88.805 -84.785 90.175 ;
        RECT -81.035 88.805 -80.255 90.175 ;
        RECT -75.645 88.805 -74.865 90.175 ;
        RECT -71.115 88.805 -70.335 90.175 ;
        RECT -65.725 88.805 -64.945 90.175 ;
        RECT -61.195 88.805 -60.415 90.175 ;
        RECT -55.805 88.805 -55.025 90.175 ;
        RECT -51.275 88.805 -50.495 90.175 ;
        RECT -45.885 88.805 -45.105 90.175 ;
        RECT -41.355 88.805 -40.575 90.175 ;
        RECT -35.965 88.805 -35.185 90.175 ;
        RECT -31.435 88.805 -30.655 90.175 ;
        RECT -26.045 88.805 -25.265 90.175 ;
        RECT -21.515 88.805 -20.735 90.175 ;
        RECT -16.125 88.805 -15.345 90.175 ;
        RECT -11.595 88.805 -10.815 90.175 ;
        RECT -6.205 88.805 -5.425 90.175 ;
        RECT -1.675 88.805 -0.895 90.175 ;
        RECT 3.715 88.805 4.495 90.175 ;
        RECT 8.245 88.805 9.025 90.175 ;
        RECT 13.635 88.805 14.415 90.175 ;
        RECT 18.165 88.805 18.945 90.175 ;
        RECT 23.555 90.015 24.335 90.175 ;
        RECT 23.555 89.230 25.125 90.015 ;
        RECT 23.555 88.805 24.335 89.230 ;
      LAYER nwell ;
        RECT -290.700 7.385 -289.095 7.620 ;
        RECT -291.400 5.860 -289.095 7.385 ;
      LAYER pwell ;
        RECT -288.675 6.055 -287.895 7.425 ;
        RECT -284.145 6.055 -283.365 7.425 ;
        RECT -278.755 6.055 -277.975 7.425 ;
        RECT -274.225 6.055 -273.445 7.425 ;
        RECT -268.835 6.055 -268.055 7.425 ;
        RECT -264.305 6.055 -263.525 7.425 ;
        RECT -258.915 6.055 -258.135 7.425 ;
        RECT -254.385 6.055 -253.605 7.425 ;
        RECT -248.995 6.055 -248.215 7.425 ;
        RECT -244.465 6.055 -243.685 7.425 ;
        RECT -239.075 6.055 -238.295 7.425 ;
        RECT -234.545 6.055 -233.765 7.425 ;
        RECT -229.155 6.055 -228.375 7.425 ;
        RECT -224.625 6.055 -223.845 7.425 ;
        RECT -219.235 6.055 -218.455 7.425 ;
        RECT -214.705 6.055 -213.925 7.425 ;
        RECT -209.315 6.055 -208.535 7.425 ;
        RECT -204.785 6.055 -204.005 7.425 ;
        RECT -199.395 6.055 -198.615 7.425 ;
        RECT -194.865 6.055 -194.085 7.425 ;
        RECT -189.475 6.055 -188.695 7.425 ;
        RECT -184.945 6.055 -184.165 7.425 ;
        RECT -179.555 6.055 -178.775 7.425 ;
        RECT -175.025 6.055 -174.245 7.425 ;
        RECT -169.635 6.055 -168.855 7.425 ;
        RECT -165.105 6.055 -164.325 7.425 ;
        RECT -159.715 6.055 -158.935 7.425 ;
        RECT -155.185 6.055 -154.405 7.425 ;
        RECT -149.795 6.055 -149.015 7.425 ;
        RECT -145.265 6.055 -144.485 7.425 ;
        RECT -139.875 6.055 -139.095 7.425 ;
        RECT -135.345 6.055 -134.565 7.425 ;
        RECT -129.955 6.055 -129.175 7.425 ;
        RECT -125.425 6.055 -124.645 7.425 ;
        RECT -120.035 6.055 -119.255 7.425 ;
        RECT -115.505 6.055 -114.725 7.425 ;
        RECT -110.115 6.055 -109.335 7.425 ;
        RECT -105.585 6.055 -104.805 7.425 ;
        RECT -100.195 6.055 -99.415 7.425 ;
        RECT -95.665 6.055 -94.885 7.425 ;
        RECT -90.275 6.055 -89.495 7.425 ;
        RECT -85.745 6.055 -84.965 7.425 ;
        RECT -80.355 6.055 -79.575 7.425 ;
        RECT -75.825 6.055 -75.045 7.425 ;
        RECT -70.435 6.055 -69.655 7.425 ;
        RECT -65.905 6.055 -65.125 7.425 ;
        RECT -60.515 6.055 -59.735 7.425 ;
        RECT -55.985 6.055 -55.205 7.425 ;
        RECT -50.595 6.055 -49.815 7.425 ;
        RECT -46.065 6.055 -45.285 7.425 ;
        RECT -40.675 6.055 -39.895 7.425 ;
        RECT -36.145 6.055 -35.365 7.425 ;
        RECT -30.755 6.055 -29.975 7.425 ;
        RECT -26.225 6.055 -25.445 7.425 ;
        RECT -20.835 6.055 -20.055 7.425 ;
        RECT -16.305 6.055 -15.525 7.425 ;
        RECT -10.915 6.055 -10.135 7.425 ;
        RECT -6.385 6.055 -5.605 7.425 ;
        RECT -0.995 6.055 -0.215 7.425 ;
        RECT 3.535 6.055 4.315 7.425 ;
        RECT 8.925 6.055 9.705 7.425 ;
        RECT 13.455 6.055 14.235 7.425 ;
        RECT 18.845 6.055 19.625 7.425 ;
        RECT 23.375 6.055 24.155 7.425 ;
      LAYER nwell ;
        RECT -291.400 5.800 -290.560 5.860 ;
      LAYER pwell ;
        RECT -290.725 5.430 -289.375 5.515 ;
        RECT -291.195 4.645 -289.375 5.430 ;
        RECT -290.725 4.605 -289.375 4.645 ;
        RECT 24.855 5.430 26.205 5.515 ;
        RECT 24.855 4.645 26.675 5.430 ;
        RECT 24.855 4.605 26.205 4.645 ;
      LAYER nwell ;
        RECT -291.400 2.710 -289.180 4.315 ;
      LAYER pwell ;
        RECT -289.105 2.305 -288.325 2.465 ;
        RECT -289.895 1.520 -288.325 2.305 ;
        RECT -289.105 1.095 -288.325 1.520 ;
        RECT -283.715 1.095 -282.935 2.465 ;
        RECT -279.185 1.095 -278.405 2.465 ;
        RECT -273.795 1.095 -273.015 2.465 ;
        RECT -269.265 1.095 -268.485 2.465 ;
        RECT -263.875 1.095 -263.095 2.465 ;
        RECT -259.345 1.095 -258.565 2.465 ;
        RECT -253.955 1.095 -253.175 2.465 ;
        RECT -249.425 1.095 -248.645 2.465 ;
        RECT -244.035 1.095 -243.255 2.465 ;
        RECT -239.505 1.095 -238.725 2.465 ;
        RECT -234.115 1.095 -233.335 2.465 ;
        RECT -229.585 1.095 -228.805 2.465 ;
        RECT -224.195 1.095 -223.415 2.465 ;
        RECT -219.665 1.095 -218.885 2.465 ;
        RECT -214.275 1.095 -213.495 2.465 ;
        RECT -209.745 1.095 -208.965 2.465 ;
        RECT -204.355 1.095 -203.575 2.465 ;
        RECT -199.825 1.095 -199.045 2.465 ;
        RECT -194.435 1.095 -193.655 2.465 ;
        RECT -189.905 1.095 -189.125 2.465 ;
        RECT -184.515 1.095 -183.735 2.465 ;
        RECT -179.985 1.095 -179.205 2.465 ;
        RECT -174.595 1.095 -173.815 2.465 ;
        RECT -170.065 1.095 -169.285 2.465 ;
        RECT -164.675 1.095 -163.895 2.465 ;
        RECT -160.145 1.095 -159.365 2.465 ;
        RECT -154.755 1.095 -153.975 2.465 ;
        RECT -150.225 1.095 -149.445 2.465 ;
        RECT -144.835 1.095 -144.055 2.465 ;
        RECT -140.305 1.095 -139.525 2.465 ;
        RECT -134.915 1.095 -134.135 2.465 ;
        RECT -130.385 1.095 -129.605 2.465 ;
        RECT -124.995 1.095 -124.215 2.465 ;
        RECT -120.465 1.095 -119.685 2.465 ;
        RECT -115.075 1.095 -114.295 2.465 ;
        RECT -110.545 1.095 -109.765 2.465 ;
        RECT -105.155 1.095 -104.375 2.465 ;
        RECT -100.625 1.095 -99.845 2.465 ;
        RECT -95.235 1.095 -94.455 2.465 ;
        RECT -90.705 1.095 -89.925 2.465 ;
        RECT -85.315 1.095 -84.535 2.465 ;
        RECT -80.785 1.095 -80.005 2.465 ;
        RECT -75.395 1.095 -74.615 2.465 ;
        RECT -70.865 1.095 -70.085 2.465 ;
        RECT -65.475 1.095 -64.695 2.465 ;
        RECT -60.945 1.095 -60.165 2.465 ;
        RECT -55.555 1.095 -54.775 2.465 ;
        RECT -51.025 1.095 -50.245 2.465 ;
        RECT -45.635 1.095 -44.855 2.465 ;
        RECT -41.105 1.095 -40.325 2.465 ;
        RECT -35.715 1.095 -34.935 2.465 ;
        RECT -31.185 1.095 -30.405 2.465 ;
        RECT -25.795 1.095 -25.015 2.465 ;
        RECT -21.265 1.095 -20.485 2.465 ;
        RECT -15.875 1.095 -15.095 2.465 ;
        RECT -11.345 1.095 -10.565 2.465 ;
        RECT -5.955 1.095 -5.175 2.465 ;
        RECT -1.425 1.095 -0.645 2.465 ;
        RECT 3.965 1.095 4.745 2.465 ;
        RECT 8.495 1.095 9.275 2.465 ;
        RECT 13.885 1.095 14.665 2.465 ;
        RECT 18.415 1.095 19.195 2.465 ;
        RECT 23.805 2.305 24.585 2.465 ;
        RECT 23.805 1.520 25.375 2.305 ;
        RECT 23.805 1.095 24.585 1.520 ;
      LAYER nwell ;
        RECT -288.940 -85.965 -287.335 -85.730 ;
        RECT -289.640 -87.490 -287.335 -85.965 ;
      LAYER pwell ;
        RECT -286.915 -87.295 -286.135 -85.925 ;
        RECT -282.385 -87.295 -281.605 -85.925 ;
        RECT -276.995 -87.295 -276.215 -85.925 ;
        RECT -272.465 -87.295 -271.685 -85.925 ;
        RECT -267.075 -87.295 -266.295 -85.925 ;
        RECT -262.545 -87.295 -261.765 -85.925 ;
        RECT -257.155 -87.295 -256.375 -85.925 ;
        RECT -252.625 -87.295 -251.845 -85.925 ;
        RECT -247.235 -87.295 -246.455 -85.925 ;
        RECT -242.705 -87.295 -241.925 -85.925 ;
        RECT -237.315 -87.295 -236.535 -85.925 ;
        RECT -232.785 -87.295 -232.005 -85.925 ;
        RECT -227.395 -87.295 -226.615 -85.925 ;
        RECT -222.865 -87.295 -222.085 -85.925 ;
        RECT -217.475 -87.295 -216.695 -85.925 ;
        RECT -212.945 -87.295 -212.165 -85.925 ;
        RECT -207.555 -87.295 -206.775 -85.925 ;
        RECT -203.025 -87.295 -202.245 -85.925 ;
        RECT -197.635 -87.295 -196.855 -85.925 ;
        RECT -193.105 -87.295 -192.325 -85.925 ;
        RECT -187.715 -87.295 -186.935 -85.925 ;
        RECT -183.185 -87.295 -182.405 -85.925 ;
        RECT -177.795 -87.295 -177.015 -85.925 ;
        RECT -173.265 -87.295 -172.485 -85.925 ;
        RECT -167.875 -87.295 -167.095 -85.925 ;
        RECT -163.345 -87.295 -162.565 -85.925 ;
        RECT -157.955 -87.295 -157.175 -85.925 ;
        RECT -153.425 -87.295 -152.645 -85.925 ;
        RECT -148.035 -87.295 -147.255 -85.925 ;
        RECT -143.505 -87.295 -142.725 -85.925 ;
        RECT -138.115 -87.295 -137.335 -85.925 ;
        RECT -133.585 -87.295 -132.805 -85.925 ;
        RECT -128.195 -87.295 -127.415 -85.925 ;
        RECT -123.665 -87.295 -122.885 -85.925 ;
        RECT -118.275 -87.295 -117.495 -85.925 ;
        RECT -113.745 -87.295 -112.965 -85.925 ;
        RECT -108.355 -87.295 -107.575 -85.925 ;
        RECT -103.825 -87.295 -103.045 -85.925 ;
        RECT -98.435 -87.295 -97.655 -85.925 ;
        RECT -93.905 -87.295 -93.125 -85.925 ;
        RECT -88.515 -87.295 -87.735 -85.925 ;
        RECT -83.985 -87.295 -83.205 -85.925 ;
        RECT -78.595 -87.295 -77.815 -85.925 ;
        RECT -74.065 -87.295 -73.285 -85.925 ;
        RECT -68.675 -87.295 -67.895 -85.925 ;
        RECT -64.145 -87.295 -63.365 -85.925 ;
        RECT -58.755 -87.295 -57.975 -85.925 ;
        RECT -54.225 -87.295 -53.445 -85.925 ;
        RECT -48.835 -87.295 -48.055 -85.925 ;
        RECT -44.305 -87.295 -43.525 -85.925 ;
        RECT -38.915 -87.295 -38.135 -85.925 ;
        RECT -34.385 -87.295 -33.605 -85.925 ;
        RECT -28.995 -87.295 -28.215 -85.925 ;
        RECT -24.465 -87.295 -23.685 -85.925 ;
        RECT -19.075 -87.295 -18.295 -85.925 ;
        RECT -14.545 -87.295 -13.765 -85.925 ;
        RECT -9.155 -87.295 -8.375 -85.925 ;
        RECT -4.625 -87.295 -3.845 -85.925 ;
        RECT 0.765 -87.295 1.545 -85.925 ;
        RECT 5.295 -87.295 6.075 -85.925 ;
        RECT 10.685 -87.295 11.465 -85.925 ;
        RECT 15.215 -87.295 15.995 -85.925 ;
        RECT 20.605 -87.295 21.385 -85.925 ;
        RECT 25.135 -87.295 25.915 -85.925 ;
      LAYER nwell ;
        RECT -289.640 -87.550 -288.800 -87.490 ;
      LAYER pwell ;
        RECT -288.965 -87.920 -287.615 -87.835 ;
        RECT -289.435 -88.705 -287.615 -87.920 ;
        RECT -288.965 -88.745 -287.615 -88.705 ;
        RECT 26.615 -87.920 27.965 -87.835 ;
        RECT 26.615 -88.705 28.435 -87.920 ;
        RECT 26.615 -88.745 27.965 -88.705 ;
      LAYER nwell ;
        RECT -289.640 -90.640 -287.420 -89.035 ;
      LAYER pwell ;
        RECT -287.345 -91.045 -286.565 -90.885 ;
        RECT -288.135 -91.830 -286.565 -91.045 ;
        RECT -287.345 -92.255 -286.565 -91.830 ;
        RECT -281.955 -92.255 -281.175 -90.885 ;
        RECT -277.425 -92.255 -276.645 -90.885 ;
        RECT -272.035 -92.255 -271.255 -90.885 ;
        RECT -267.505 -92.255 -266.725 -90.885 ;
        RECT -262.115 -92.255 -261.335 -90.885 ;
        RECT -257.585 -92.255 -256.805 -90.885 ;
        RECT -252.195 -92.255 -251.415 -90.885 ;
        RECT -247.665 -92.255 -246.885 -90.885 ;
        RECT -242.275 -92.255 -241.495 -90.885 ;
        RECT -237.745 -92.255 -236.965 -90.885 ;
        RECT -232.355 -92.255 -231.575 -90.885 ;
        RECT -227.825 -92.255 -227.045 -90.885 ;
        RECT -222.435 -92.255 -221.655 -90.885 ;
        RECT -217.905 -92.255 -217.125 -90.885 ;
        RECT -212.515 -92.255 -211.735 -90.885 ;
        RECT -207.985 -92.255 -207.205 -90.885 ;
        RECT -202.595 -92.255 -201.815 -90.885 ;
        RECT -198.065 -92.255 -197.285 -90.885 ;
        RECT -192.675 -92.255 -191.895 -90.885 ;
        RECT -188.145 -92.255 -187.365 -90.885 ;
        RECT -182.755 -92.255 -181.975 -90.885 ;
        RECT -178.225 -92.255 -177.445 -90.885 ;
        RECT -172.835 -92.255 -172.055 -90.885 ;
        RECT -168.305 -92.255 -167.525 -90.885 ;
        RECT -162.915 -92.255 -162.135 -90.885 ;
        RECT -158.385 -92.255 -157.605 -90.885 ;
        RECT -152.995 -92.255 -152.215 -90.885 ;
        RECT -148.465 -92.255 -147.685 -90.885 ;
        RECT -143.075 -92.255 -142.295 -90.885 ;
        RECT -138.545 -92.255 -137.765 -90.885 ;
        RECT -133.155 -92.255 -132.375 -90.885 ;
        RECT -128.625 -92.255 -127.845 -90.885 ;
        RECT -123.235 -92.255 -122.455 -90.885 ;
        RECT -118.705 -92.255 -117.925 -90.885 ;
        RECT -113.315 -92.255 -112.535 -90.885 ;
        RECT -108.785 -92.255 -108.005 -90.885 ;
        RECT -103.395 -92.255 -102.615 -90.885 ;
        RECT -98.865 -92.255 -98.085 -90.885 ;
        RECT -93.475 -92.255 -92.695 -90.885 ;
        RECT -88.945 -92.255 -88.165 -90.885 ;
        RECT -83.555 -92.255 -82.775 -90.885 ;
        RECT -79.025 -92.255 -78.245 -90.885 ;
        RECT -73.635 -92.255 -72.855 -90.885 ;
        RECT -69.105 -92.255 -68.325 -90.885 ;
        RECT -63.715 -92.255 -62.935 -90.885 ;
        RECT -59.185 -92.255 -58.405 -90.885 ;
        RECT -53.795 -92.255 -53.015 -90.885 ;
        RECT -49.265 -92.255 -48.485 -90.885 ;
        RECT -43.875 -92.255 -43.095 -90.885 ;
        RECT -39.345 -92.255 -38.565 -90.885 ;
        RECT -33.955 -92.255 -33.175 -90.885 ;
        RECT -29.425 -92.255 -28.645 -90.885 ;
        RECT -24.035 -92.255 -23.255 -90.885 ;
        RECT -19.505 -92.255 -18.725 -90.885 ;
        RECT -14.115 -92.255 -13.335 -90.885 ;
        RECT -9.585 -92.255 -8.805 -90.885 ;
        RECT -4.195 -92.255 -3.415 -90.885 ;
        RECT 0.335 -92.255 1.115 -90.885 ;
        RECT 5.725 -92.255 6.505 -90.885 ;
        RECT 10.255 -92.255 11.035 -90.885 ;
        RECT 15.645 -92.255 16.425 -90.885 ;
        RECT 20.175 -92.255 20.955 -90.885 ;
        RECT 25.565 -91.045 26.345 -90.885 ;
        RECT 25.565 -91.830 27.135 -91.045 ;
        RECT 25.565 -92.255 26.345 -91.830 ;
      LAYER nwell ;
        RECT -288.690 -173.675 -287.085 -173.440 ;
        RECT -289.390 -175.200 -287.085 -173.675 ;
      LAYER pwell ;
        RECT -286.665 -175.005 -285.885 -173.635 ;
        RECT -282.135 -175.005 -281.355 -173.635 ;
        RECT -276.745 -175.005 -275.965 -173.635 ;
        RECT -272.215 -175.005 -271.435 -173.635 ;
        RECT -266.825 -175.005 -266.045 -173.635 ;
        RECT -262.295 -175.005 -261.515 -173.635 ;
        RECT -256.905 -175.005 -256.125 -173.635 ;
        RECT -252.375 -175.005 -251.595 -173.635 ;
        RECT -246.985 -175.005 -246.205 -173.635 ;
        RECT -242.455 -175.005 -241.675 -173.635 ;
        RECT -237.065 -175.005 -236.285 -173.635 ;
        RECT -232.535 -175.005 -231.755 -173.635 ;
        RECT -227.145 -175.005 -226.365 -173.635 ;
        RECT -222.615 -175.005 -221.835 -173.635 ;
        RECT -217.225 -175.005 -216.445 -173.635 ;
        RECT -212.695 -175.005 -211.915 -173.635 ;
        RECT -207.305 -175.005 -206.525 -173.635 ;
        RECT -202.775 -175.005 -201.995 -173.635 ;
        RECT -197.385 -175.005 -196.605 -173.635 ;
        RECT -192.855 -175.005 -192.075 -173.635 ;
        RECT -187.465 -175.005 -186.685 -173.635 ;
        RECT -182.935 -175.005 -182.155 -173.635 ;
        RECT -177.545 -175.005 -176.765 -173.635 ;
        RECT -173.015 -175.005 -172.235 -173.635 ;
        RECT -167.625 -175.005 -166.845 -173.635 ;
        RECT -163.095 -175.005 -162.315 -173.635 ;
        RECT -157.705 -175.005 -156.925 -173.635 ;
        RECT -153.175 -175.005 -152.395 -173.635 ;
        RECT -147.785 -175.005 -147.005 -173.635 ;
        RECT -143.255 -175.005 -142.475 -173.635 ;
        RECT -137.865 -175.005 -137.085 -173.635 ;
        RECT -133.335 -175.005 -132.555 -173.635 ;
        RECT -127.945 -175.005 -127.165 -173.635 ;
        RECT -123.415 -175.005 -122.635 -173.635 ;
        RECT -118.025 -175.005 -117.245 -173.635 ;
        RECT -113.495 -175.005 -112.715 -173.635 ;
        RECT -108.105 -175.005 -107.325 -173.635 ;
        RECT -103.575 -175.005 -102.795 -173.635 ;
        RECT -98.185 -175.005 -97.405 -173.635 ;
        RECT -93.655 -175.005 -92.875 -173.635 ;
        RECT -88.265 -175.005 -87.485 -173.635 ;
        RECT -83.735 -175.005 -82.955 -173.635 ;
        RECT -78.345 -175.005 -77.565 -173.635 ;
        RECT -73.815 -175.005 -73.035 -173.635 ;
        RECT -68.425 -175.005 -67.645 -173.635 ;
        RECT -63.895 -175.005 -63.115 -173.635 ;
        RECT -58.505 -175.005 -57.725 -173.635 ;
        RECT -53.975 -175.005 -53.195 -173.635 ;
        RECT -48.585 -175.005 -47.805 -173.635 ;
        RECT -44.055 -175.005 -43.275 -173.635 ;
        RECT -38.665 -175.005 -37.885 -173.635 ;
        RECT -34.135 -175.005 -33.355 -173.635 ;
        RECT -28.745 -175.005 -27.965 -173.635 ;
        RECT -24.215 -175.005 -23.435 -173.635 ;
        RECT -18.825 -175.005 -18.045 -173.635 ;
        RECT -14.295 -175.005 -13.515 -173.635 ;
        RECT -8.905 -175.005 -8.125 -173.635 ;
        RECT -4.375 -175.005 -3.595 -173.635 ;
        RECT 1.015 -175.005 1.795 -173.635 ;
        RECT 5.545 -175.005 6.325 -173.635 ;
        RECT 10.935 -175.005 11.715 -173.635 ;
        RECT 15.465 -175.005 16.245 -173.635 ;
        RECT 20.855 -175.005 21.635 -173.635 ;
        RECT 25.385 -175.005 26.165 -173.635 ;
      LAYER nwell ;
        RECT -289.390 -175.260 -288.550 -175.200 ;
      LAYER pwell ;
        RECT -288.715 -175.630 -287.365 -175.545 ;
        RECT -289.185 -176.415 -287.365 -175.630 ;
        RECT -288.715 -176.455 -287.365 -176.415 ;
        RECT 26.865 -175.630 28.215 -175.545 ;
        RECT 26.865 -176.415 28.685 -175.630 ;
        RECT 26.865 -176.455 28.215 -176.415 ;
      LAYER nwell ;
        RECT -289.390 -178.350 -287.170 -176.745 ;
      LAYER pwell ;
        RECT -287.095 -178.755 -286.315 -178.595 ;
        RECT -287.885 -179.540 -286.315 -178.755 ;
        RECT -287.095 -179.965 -286.315 -179.540 ;
        RECT -281.705 -179.965 -280.925 -178.595 ;
        RECT -277.175 -179.965 -276.395 -178.595 ;
        RECT -271.785 -179.965 -271.005 -178.595 ;
        RECT -267.255 -179.965 -266.475 -178.595 ;
        RECT -261.865 -179.965 -261.085 -178.595 ;
        RECT -257.335 -179.965 -256.555 -178.595 ;
        RECT -251.945 -179.965 -251.165 -178.595 ;
        RECT -247.415 -179.965 -246.635 -178.595 ;
        RECT -242.025 -179.965 -241.245 -178.595 ;
        RECT -237.495 -179.965 -236.715 -178.595 ;
        RECT -232.105 -179.965 -231.325 -178.595 ;
        RECT -227.575 -179.965 -226.795 -178.595 ;
        RECT -222.185 -179.965 -221.405 -178.595 ;
        RECT -217.655 -179.965 -216.875 -178.595 ;
        RECT -212.265 -179.965 -211.485 -178.595 ;
        RECT -207.735 -179.965 -206.955 -178.595 ;
        RECT -202.345 -179.965 -201.565 -178.595 ;
        RECT -197.815 -179.965 -197.035 -178.595 ;
        RECT -192.425 -179.965 -191.645 -178.595 ;
        RECT -187.895 -179.965 -187.115 -178.595 ;
        RECT -182.505 -179.965 -181.725 -178.595 ;
        RECT -177.975 -179.965 -177.195 -178.595 ;
        RECT -172.585 -179.965 -171.805 -178.595 ;
        RECT -168.055 -179.965 -167.275 -178.595 ;
        RECT -162.665 -179.965 -161.885 -178.595 ;
        RECT -158.135 -179.965 -157.355 -178.595 ;
        RECT -152.745 -179.965 -151.965 -178.595 ;
        RECT -148.215 -179.965 -147.435 -178.595 ;
        RECT -142.825 -179.965 -142.045 -178.595 ;
        RECT -138.295 -179.965 -137.515 -178.595 ;
        RECT -132.905 -179.965 -132.125 -178.595 ;
        RECT -128.375 -179.965 -127.595 -178.595 ;
        RECT -122.985 -179.965 -122.205 -178.595 ;
        RECT -118.455 -179.965 -117.675 -178.595 ;
        RECT -113.065 -179.965 -112.285 -178.595 ;
        RECT -108.535 -179.965 -107.755 -178.595 ;
        RECT -103.145 -179.965 -102.365 -178.595 ;
        RECT -98.615 -179.965 -97.835 -178.595 ;
        RECT -93.225 -179.965 -92.445 -178.595 ;
        RECT -88.695 -179.965 -87.915 -178.595 ;
        RECT -83.305 -179.965 -82.525 -178.595 ;
        RECT -78.775 -179.965 -77.995 -178.595 ;
        RECT -73.385 -179.965 -72.605 -178.595 ;
        RECT -68.855 -179.965 -68.075 -178.595 ;
        RECT -63.465 -179.965 -62.685 -178.595 ;
        RECT -58.935 -179.965 -58.155 -178.595 ;
        RECT -53.545 -179.965 -52.765 -178.595 ;
        RECT -49.015 -179.965 -48.235 -178.595 ;
        RECT -43.625 -179.965 -42.845 -178.595 ;
        RECT -39.095 -179.965 -38.315 -178.595 ;
        RECT -33.705 -179.965 -32.925 -178.595 ;
        RECT -29.175 -179.965 -28.395 -178.595 ;
        RECT -23.785 -179.965 -23.005 -178.595 ;
        RECT -19.255 -179.965 -18.475 -178.595 ;
        RECT -13.865 -179.965 -13.085 -178.595 ;
        RECT -9.335 -179.965 -8.555 -178.595 ;
        RECT -3.945 -179.965 -3.165 -178.595 ;
        RECT 0.585 -179.965 1.365 -178.595 ;
        RECT 5.975 -179.965 6.755 -178.595 ;
        RECT 10.505 -179.965 11.285 -178.595 ;
        RECT 15.895 -179.965 16.675 -178.595 ;
        RECT 20.425 -179.965 21.205 -178.595 ;
        RECT 25.815 -178.755 26.595 -178.595 ;
        RECT 25.815 -179.540 27.385 -178.755 ;
        RECT 25.815 -179.965 26.595 -179.540 ;
      LAYER li1 ;
        RECT -290.845 94.990 -290.675 95.140 ;
        RECT -291.460 94.820 -290.675 94.990 ;
        RECT -291.375 93.655 -291.085 94.820 ;
        RECT -290.845 94.615 -290.675 94.820 ;
        RECT -290.505 94.875 -288.295 95.055 ;
        RECT -290.505 94.785 -289.600 94.875 ;
        RECT -288.800 94.795 -288.295 94.875 ;
        RECT -280.585 94.875 -278.375 95.055 ;
        RECT -280.585 94.785 -279.680 94.875 ;
        RECT -278.880 94.795 -278.375 94.875 ;
        RECT -270.665 94.875 -268.455 95.055 ;
        RECT -270.665 94.785 -269.760 94.875 ;
        RECT -268.960 94.795 -268.455 94.875 ;
        RECT -260.745 94.875 -258.535 95.055 ;
        RECT -260.745 94.785 -259.840 94.875 ;
        RECT -259.040 94.795 -258.535 94.875 ;
        RECT -250.825 94.875 -248.615 95.055 ;
        RECT -250.825 94.785 -249.920 94.875 ;
        RECT -249.120 94.795 -248.615 94.875 ;
        RECT -240.905 94.875 -238.695 95.055 ;
        RECT -240.905 94.785 -240.000 94.875 ;
        RECT -239.200 94.795 -238.695 94.875 ;
        RECT -230.985 94.875 -228.775 95.055 ;
        RECT -230.985 94.785 -230.080 94.875 ;
        RECT -229.280 94.795 -228.775 94.875 ;
        RECT -221.065 94.875 -218.855 95.055 ;
        RECT -221.065 94.785 -220.160 94.875 ;
        RECT -219.360 94.795 -218.855 94.875 ;
        RECT -211.145 94.875 -208.935 95.055 ;
        RECT -211.145 94.785 -210.240 94.875 ;
        RECT -209.440 94.795 -208.935 94.875 ;
        RECT -201.225 94.875 -199.015 95.055 ;
        RECT -201.225 94.785 -200.320 94.875 ;
        RECT -199.520 94.795 -199.015 94.875 ;
        RECT -191.305 94.875 -189.095 95.055 ;
        RECT -191.305 94.785 -190.400 94.875 ;
        RECT -189.600 94.795 -189.095 94.875 ;
        RECT -181.385 94.875 -179.175 95.055 ;
        RECT -181.385 94.785 -180.480 94.875 ;
        RECT -179.680 94.795 -179.175 94.875 ;
        RECT -171.465 94.875 -169.255 95.055 ;
        RECT -171.465 94.785 -170.560 94.875 ;
        RECT -169.760 94.795 -169.255 94.875 ;
        RECT -161.545 94.875 -159.335 95.055 ;
        RECT -161.545 94.785 -160.640 94.875 ;
        RECT -159.840 94.795 -159.335 94.875 ;
        RECT -151.625 94.875 -149.415 95.055 ;
        RECT -151.625 94.785 -150.720 94.875 ;
        RECT -149.920 94.795 -149.415 94.875 ;
        RECT -141.705 94.875 -139.495 95.055 ;
        RECT -141.705 94.785 -140.800 94.875 ;
        RECT -140.000 94.795 -139.495 94.875 ;
        RECT -131.785 94.875 -129.575 95.055 ;
        RECT -131.785 94.785 -130.880 94.875 ;
        RECT -130.080 94.795 -129.575 94.875 ;
        RECT -121.865 94.875 -119.655 95.055 ;
        RECT -121.865 94.785 -120.960 94.875 ;
        RECT -120.160 94.795 -119.655 94.875 ;
        RECT -111.945 94.875 -109.735 95.055 ;
        RECT -111.945 94.785 -111.040 94.875 ;
        RECT -110.240 94.795 -109.735 94.875 ;
        RECT -102.025 94.875 -99.815 95.055 ;
        RECT -102.025 94.785 -101.120 94.875 ;
        RECT -100.320 94.795 -99.815 94.875 ;
        RECT -92.105 94.875 -89.895 95.055 ;
        RECT -92.105 94.785 -91.200 94.875 ;
        RECT -90.400 94.795 -89.895 94.875 ;
        RECT -82.185 94.875 -79.975 95.055 ;
        RECT -82.185 94.785 -81.280 94.875 ;
        RECT -80.480 94.795 -79.975 94.875 ;
        RECT -72.265 94.875 -70.055 95.055 ;
        RECT -72.265 94.785 -71.360 94.875 ;
        RECT -70.560 94.795 -70.055 94.875 ;
        RECT -62.345 94.875 -60.135 95.055 ;
        RECT -62.345 94.785 -61.440 94.875 ;
        RECT -60.640 94.795 -60.135 94.875 ;
        RECT -52.425 94.875 -50.215 95.055 ;
        RECT -52.425 94.785 -51.520 94.875 ;
        RECT -50.720 94.795 -50.215 94.875 ;
        RECT -42.505 94.875 -40.295 95.055 ;
        RECT -42.505 94.785 -41.600 94.875 ;
        RECT -40.800 94.795 -40.295 94.875 ;
        RECT -32.585 94.875 -30.375 95.055 ;
        RECT -32.585 94.785 -31.680 94.875 ;
        RECT -30.880 94.795 -30.375 94.875 ;
        RECT -22.665 94.875 -20.455 95.055 ;
        RECT -22.665 94.785 -21.760 94.875 ;
        RECT -20.960 94.795 -20.455 94.875 ;
        RECT -12.745 94.875 -10.535 95.055 ;
        RECT -12.745 94.785 -11.840 94.875 ;
        RECT -11.040 94.795 -10.535 94.875 ;
        RECT -2.825 94.875 -0.615 95.055 ;
        RECT -2.825 94.785 -1.920 94.875 ;
        RECT -1.120 94.795 -0.615 94.875 ;
        RECT 7.095 94.875 9.305 95.055 ;
        RECT 7.095 94.785 8.000 94.875 ;
        RECT 8.800 94.795 9.305 94.875 ;
        RECT 17.015 94.875 19.225 95.055 ;
        RECT 17.015 94.785 17.920 94.875 ;
        RECT 18.720 94.795 19.225 94.875 ;
        RECT -290.845 94.285 -289.915 94.615 ;
        RECT -289.430 94.600 -289.100 94.705 ;
        RECT -283.440 94.600 -283.110 94.705 ;
        RECT -279.510 94.600 -279.180 94.705 ;
        RECT -273.520 94.600 -273.190 94.705 ;
        RECT -269.590 94.600 -269.260 94.705 ;
        RECT -263.600 94.600 -263.270 94.705 ;
        RECT -259.670 94.600 -259.340 94.705 ;
        RECT -253.680 94.600 -253.350 94.705 ;
        RECT -249.750 94.600 -249.420 94.705 ;
        RECT -243.760 94.600 -243.430 94.705 ;
        RECT -239.830 94.600 -239.500 94.705 ;
        RECT -233.840 94.600 -233.510 94.705 ;
        RECT -229.910 94.600 -229.580 94.705 ;
        RECT -223.920 94.600 -223.590 94.705 ;
        RECT -219.990 94.600 -219.660 94.705 ;
        RECT -214.000 94.600 -213.670 94.705 ;
        RECT -210.070 94.600 -209.740 94.705 ;
        RECT -204.080 94.600 -203.750 94.705 ;
        RECT -200.150 94.600 -199.820 94.705 ;
        RECT -194.160 94.600 -193.830 94.705 ;
        RECT -190.230 94.600 -189.900 94.705 ;
        RECT -184.240 94.600 -183.910 94.705 ;
        RECT -180.310 94.600 -179.980 94.705 ;
        RECT -174.320 94.600 -173.990 94.705 ;
        RECT -170.390 94.600 -170.060 94.705 ;
        RECT -164.400 94.600 -164.070 94.705 ;
        RECT -160.470 94.600 -160.140 94.705 ;
        RECT -154.480 94.600 -154.150 94.705 ;
        RECT -150.550 94.600 -150.220 94.705 ;
        RECT -144.560 94.600 -144.230 94.705 ;
        RECT -140.630 94.600 -140.300 94.705 ;
        RECT -134.640 94.600 -134.310 94.705 ;
        RECT -130.710 94.600 -130.380 94.705 ;
        RECT -124.720 94.600 -124.390 94.705 ;
        RECT -120.790 94.600 -120.460 94.705 ;
        RECT -114.800 94.600 -114.470 94.705 ;
        RECT -110.870 94.600 -110.540 94.705 ;
        RECT -104.880 94.600 -104.550 94.705 ;
        RECT -100.950 94.600 -100.620 94.705 ;
        RECT -94.960 94.600 -94.630 94.705 ;
        RECT -91.030 94.600 -90.700 94.705 ;
        RECT -85.040 94.600 -84.710 94.705 ;
        RECT -81.110 94.600 -80.780 94.705 ;
        RECT -75.120 94.600 -74.790 94.705 ;
        RECT -71.190 94.600 -70.860 94.705 ;
        RECT -65.200 94.600 -64.870 94.705 ;
        RECT -61.270 94.600 -60.940 94.705 ;
        RECT -55.280 94.600 -54.950 94.705 ;
        RECT -51.350 94.600 -51.020 94.705 ;
        RECT -45.360 94.600 -45.030 94.705 ;
        RECT -41.430 94.600 -41.100 94.705 ;
        RECT -35.440 94.600 -35.110 94.705 ;
        RECT -31.510 94.600 -31.180 94.705 ;
        RECT -25.520 94.600 -25.190 94.705 ;
        RECT -21.590 94.600 -21.260 94.705 ;
        RECT -15.600 94.600 -15.270 94.705 ;
        RECT -11.670 94.600 -11.340 94.705 ;
        RECT -5.680 94.600 -5.350 94.705 ;
        RECT -1.750 94.600 -1.420 94.705 ;
        RECT 4.240 94.600 4.570 94.705 ;
        RECT 8.170 94.600 8.500 94.705 ;
        RECT 14.160 94.600 14.490 94.705 ;
        RECT 18.090 94.600 18.420 94.705 ;
        RECT 24.080 94.600 24.410 94.705 ;
        RECT -289.745 94.430 -288.675 94.600 ;
        RECT -290.845 93.760 -290.675 94.285 ;
        RECT -289.745 94.105 -289.575 94.430 ;
        RECT -290.505 93.925 -289.575 94.105 ;
        RECT -289.395 93.865 -289.025 94.205 ;
        RECT -288.845 94.105 -288.675 94.430 ;
        RECT -283.865 94.430 -282.795 94.600 ;
        RECT -283.865 94.105 -283.695 94.430 ;
        RECT -288.845 93.935 -288.295 94.105 ;
        RECT -284.245 93.935 -283.695 94.105 ;
        RECT -283.515 93.865 -283.145 94.205 ;
        RECT -282.965 94.105 -282.795 94.430 ;
        RECT -279.825 94.430 -278.755 94.600 ;
        RECT -279.825 94.105 -279.655 94.430 ;
        RECT -282.965 93.925 -282.035 94.105 ;
        RECT -280.585 93.925 -279.655 94.105 ;
        RECT -279.475 93.865 -279.105 94.205 ;
        RECT -278.925 94.105 -278.755 94.430 ;
        RECT -273.945 94.430 -272.875 94.600 ;
        RECT -273.945 94.105 -273.775 94.430 ;
        RECT -278.925 93.935 -278.375 94.105 ;
        RECT -274.325 93.935 -273.775 94.105 ;
        RECT -273.595 93.865 -273.225 94.205 ;
        RECT -273.045 94.105 -272.875 94.430 ;
        RECT -269.905 94.430 -268.835 94.600 ;
        RECT -269.905 94.105 -269.735 94.430 ;
        RECT -273.045 93.925 -272.115 94.105 ;
        RECT -270.665 93.925 -269.735 94.105 ;
        RECT -269.555 93.865 -269.185 94.205 ;
        RECT -269.005 94.105 -268.835 94.430 ;
        RECT -264.025 94.430 -262.955 94.600 ;
        RECT -264.025 94.105 -263.855 94.430 ;
        RECT -269.005 93.935 -268.455 94.105 ;
        RECT -264.405 93.935 -263.855 94.105 ;
        RECT -263.675 93.865 -263.305 94.205 ;
        RECT -263.125 94.105 -262.955 94.430 ;
        RECT -259.985 94.430 -258.915 94.600 ;
        RECT -259.985 94.105 -259.815 94.430 ;
        RECT -263.125 93.925 -262.195 94.105 ;
        RECT -260.745 93.925 -259.815 94.105 ;
        RECT -259.635 93.865 -259.265 94.205 ;
        RECT -259.085 94.105 -258.915 94.430 ;
        RECT -254.105 94.430 -253.035 94.600 ;
        RECT -254.105 94.105 -253.935 94.430 ;
        RECT -259.085 93.935 -258.535 94.105 ;
        RECT -254.485 93.935 -253.935 94.105 ;
        RECT -253.755 93.865 -253.385 94.205 ;
        RECT -253.205 94.105 -253.035 94.430 ;
        RECT -250.065 94.430 -248.995 94.600 ;
        RECT -250.065 94.105 -249.895 94.430 ;
        RECT -253.205 93.925 -252.275 94.105 ;
        RECT -250.825 93.925 -249.895 94.105 ;
        RECT -249.715 93.865 -249.345 94.205 ;
        RECT -249.165 94.105 -248.995 94.430 ;
        RECT -244.185 94.430 -243.115 94.600 ;
        RECT -244.185 94.105 -244.015 94.430 ;
        RECT -249.165 93.935 -248.615 94.105 ;
        RECT -244.565 93.935 -244.015 94.105 ;
        RECT -243.835 93.865 -243.465 94.205 ;
        RECT -243.285 94.105 -243.115 94.430 ;
        RECT -240.145 94.430 -239.075 94.600 ;
        RECT -240.145 94.105 -239.975 94.430 ;
        RECT -243.285 93.925 -242.355 94.105 ;
        RECT -240.905 93.925 -239.975 94.105 ;
        RECT -239.795 93.865 -239.425 94.205 ;
        RECT -239.245 94.105 -239.075 94.430 ;
        RECT -234.265 94.430 -233.195 94.600 ;
        RECT -234.265 94.105 -234.095 94.430 ;
        RECT -239.245 93.935 -238.695 94.105 ;
        RECT -234.645 93.935 -234.095 94.105 ;
        RECT -233.915 93.865 -233.545 94.205 ;
        RECT -233.365 94.105 -233.195 94.430 ;
        RECT -230.225 94.430 -229.155 94.600 ;
        RECT -230.225 94.105 -230.055 94.430 ;
        RECT -233.365 93.925 -232.435 94.105 ;
        RECT -230.985 93.925 -230.055 94.105 ;
        RECT -229.875 93.865 -229.505 94.205 ;
        RECT -229.325 94.105 -229.155 94.430 ;
        RECT -224.345 94.430 -223.275 94.600 ;
        RECT -224.345 94.105 -224.175 94.430 ;
        RECT -229.325 93.935 -228.775 94.105 ;
        RECT -224.725 93.935 -224.175 94.105 ;
        RECT -223.995 93.865 -223.625 94.205 ;
        RECT -223.445 94.105 -223.275 94.430 ;
        RECT -220.305 94.430 -219.235 94.600 ;
        RECT -220.305 94.105 -220.135 94.430 ;
        RECT -223.445 93.925 -222.515 94.105 ;
        RECT -221.065 93.925 -220.135 94.105 ;
        RECT -219.955 93.865 -219.585 94.205 ;
        RECT -219.405 94.105 -219.235 94.430 ;
        RECT -214.425 94.430 -213.355 94.600 ;
        RECT -214.425 94.105 -214.255 94.430 ;
        RECT -219.405 93.935 -218.855 94.105 ;
        RECT -214.805 93.935 -214.255 94.105 ;
        RECT -214.075 93.865 -213.705 94.205 ;
        RECT -213.525 94.105 -213.355 94.430 ;
        RECT -210.385 94.430 -209.315 94.600 ;
        RECT -210.385 94.105 -210.215 94.430 ;
        RECT -213.525 93.925 -212.595 94.105 ;
        RECT -211.145 93.925 -210.215 94.105 ;
        RECT -210.035 93.865 -209.665 94.205 ;
        RECT -209.485 94.105 -209.315 94.430 ;
        RECT -204.505 94.430 -203.435 94.600 ;
        RECT -204.505 94.105 -204.335 94.430 ;
        RECT -209.485 93.935 -208.935 94.105 ;
        RECT -204.885 93.935 -204.335 94.105 ;
        RECT -204.155 93.865 -203.785 94.205 ;
        RECT -203.605 94.105 -203.435 94.430 ;
        RECT -200.465 94.430 -199.395 94.600 ;
        RECT -200.465 94.105 -200.295 94.430 ;
        RECT -203.605 93.925 -202.675 94.105 ;
        RECT -201.225 93.925 -200.295 94.105 ;
        RECT -200.115 93.865 -199.745 94.205 ;
        RECT -199.565 94.105 -199.395 94.430 ;
        RECT -194.585 94.430 -193.515 94.600 ;
        RECT -194.585 94.105 -194.415 94.430 ;
        RECT -199.565 93.935 -199.015 94.105 ;
        RECT -194.965 93.935 -194.415 94.105 ;
        RECT -194.235 93.865 -193.865 94.205 ;
        RECT -193.685 94.105 -193.515 94.430 ;
        RECT -190.545 94.430 -189.475 94.600 ;
        RECT -190.545 94.105 -190.375 94.430 ;
        RECT -193.685 93.925 -192.755 94.105 ;
        RECT -191.305 93.925 -190.375 94.105 ;
        RECT -190.195 93.865 -189.825 94.205 ;
        RECT -189.645 94.105 -189.475 94.430 ;
        RECT -184.665 94.430 -183.595 94.600 ;
        RECT -184.665 94.105 -184.495 94.430 ;
        RECT -189.645 93.935 -189.095 94.105 ;
        RECT -185.045 93.935 -184.495 94.105 ;
        RECT -184.315 93.865 -183.945 94.205 ;
        RECT -183.765 94.105 -183.595 94.430 ;
        RECT -180.625 94.430 -179.555 94.600 ;
        RECT -180.625 94.105 -180.455 94.430 ;
        RECT -183.765 93.925 -182.835 94.105 ;
        RECT -181.385 93.925 -180.455 94.105 ;
        RECT -180.275 93.865 -179.905 94.205 ;
        RECT -179.725 94.105 -179.555 94.430 ;
        RECT -174.745 94.430 -173.675 94.600 ;
        RECT -174.745 94.105 -174.575 94.430 ;
        RECT -179.725 93.935 -179.175 94.105 ;
        RECT -175.125 93.935 -174.575 94.105 ;
        RECT -174.395 93.865 -174.025 94.205 ;
        RECT -173.845 94.105 -173.675 94.430 ;
        RECT -170.705 94.430 -169.635 94.600 ;
        RECT -170.705 94.105 -170.535 94.430 ;
        RECT -173.845 93.925 -172.915 94.105 ;
        RECT -171.465 93.925 -170.535 94.105 ;
        RECT -170.355 93.865 -169.985 94.205 ;
        RECT -169.805 94.105 -169.635 94.430 ;
        RECT -164.825 94.430 -163.755 94.600 ;
        RECT -164.825 94.105 -164.655 94.430 ;
        RECT -169.805 93.935 -169.255 94.105 ;
        RECT -165.205 93.935 -164.655 94.105 ;
        RECT -164.475 93.865 -164.105 94.205 ;
        RECT -163.925 94.105 -163.755 94.430 ;
        RECT -160.785 94.430 -159.715 94.600 ;
        RECT -160.785 94.105 -160.615 94.430 ;
        RECT -163.925 93.925 -162.995 94.105 ;
        RECT -161.545 93.925 -160.615 94.105 ;
        RECT -160.435 93.865 -160.065 94.205 ;
        RECT -159.885 94.105 -159.715 94.430 ;
        RECT -154.905 94.430 -153.835 94.600 ;
        RECT -154.905 94.105 -154.735 94.430 ;
        RECT -159.885 93.935 -159.335 94.105 ;
        RECT -155.285 93.935 -154.735 94.105 ;
        RECT -154.555 93.865 -154.185 94.205 ;
        RECT -154.005 94.105 -153.835 94.430 ;
        RECT -150.865 94.430 -149.795 94.600 ;
        RECT -150.865 94.105 -150.695 94.430 ;
        RECT -154.005 93.925 -153.075 94.105 ;
        RECT -151.625 93.925 -150.695 94.105 ;
        RECT -150.515 93.865 -150.145 94.205 ;
        RECT -149.965 94.105 -149.795 94.430 ;
        RECT -144.985 94.430 -143.915 94.600 ;
        RECT -144.985 94.105 -144.815 94.430 ;
        RECT -149.965 93.935 -149.415 94.105 ;
        RECT -145.365 93.935 -144.815 94.105 ;
        RECT -144.635 93.865 -144.265 94.205 ;
        RECT -144.085 94.105 -143.915 94.430 ;
        RECT -140.945 94.430 -139.875 94.600 ;
        RECT -140.945 94.105 -140.775 94.430 ;
        RECT -144.085 93.925 -143.155 94.105 ;
        RECT -141.705 93.925 -140.775 94.105 ;
        RECT -140.595 93.865 -140.225 94.205 ;
        RECT -140.045 94.105 -139.875 94.430 ;
        RECT -135.065 94.430 -133.995 94.600 ;
        RECT -135.065 94.105 -134.895 94.430 ;
        RECT -140.045 93.935 -139.495 94.105 ;
        RECT -135.445 93.935 -134.895 94.105 ;
        RECT -134.715 93.865 -134.345 94.205 ;
        RECT -134.165 94.105 -133.995 94.430 ;
        RECT -131.025 94.430 -129.955 94.600 ;
        RECT -131.025 94.105 -130.855 94.430 ;
        RECT -134.165 93.925 -133.235 94.105 ;
        RECT -131.785 93.925 -130.855 94.105 ;
        RECT -130.675 93.865 -130.305 94.205 ;
        RECT -130.125 94.105 -129.955 94.430 ;
        RECT -125.145 94.430 -124.075 94.600 ;
        RECT -125.145 94.105 -124.975 94.430 ;
        RECT -130.125 93.935 -129.575 94.105 ;
        RECT -125.525 93.935 -124.975 94.105 ;
        RECT -124.795 93.865 -124.425 94.205 ;
        RECT -124.245 94.105 -124.075 94.430 ;
        RECT -121.105 94.430 -120.035 94.600 ;
        RECT -121.105 94.105 -120.935 94.430 ;
        RECT -124.245 93.925 -123.315 94.105 ;
        RECT -121.865 93.925 -120.935 94.105 ;
        RECT -120.755 93.865 -120.385 94.205 ;
        RECT -120.205 94.105 -120.035 94.430 ;
        RECT -115.225 94.430 -114.155 94.600 ;
        RECT -115.225 94.105 -115.055 94.430 ;
        RECT -120.205 93.935 -119.655 94.105 ;
        RECT -115.605 93.935 -115.055 94.105 ;
        RECT -114.875 93.865 -114.505 94.205 ;
        RECT -114.325 94.105 -114.155 94.430 ;
        RECT -111.185 94.430 -110.115 94.600 ;
        RECT -111.185 94.105 -111.015 94.430 ;
        RECT -114.325 93.925 -113.395 94.105 ;
        RECT -111.945 93.925 -111.015 94.105 ;
        RECT -110.835 93.865 -110.465 94.205 ;
        RECT -110.285 94.105 -110.115 94.430 ;
        RECT -105.305 94.430 -104.235 94.600 ;
        RECT -105.305 94.105 -105.135 94.430 ;
        RECT -110.285 93.935 -109.735 94.105 ;
        RECT -105.685 93.935 -105.135 94.105 ;
        RECT -104.955 93.865 -104.585 94.205 ;
        RECT -104.405 94.105 -104.235 94.430 ;
        RECT -101.265 94.430 -100.195 94.600 ;
        RECT -101.265 94.105 -101.095 94.430 ;
        RECT -104.405 93.925 -103.475 94.105 ;
        RECT -102.025 93.925 -101.095 94.105 ;
        RECT -100.915 93.865 -100.545 94.205 ;
        RECT -100.365 94.105 -100.195 94.430 ;
        RECT -95.385 94.430 -94.315 94.600 ;
        RECT -95.385 94.105 -95.215 94.430 ;
        RECT -100.365 93.935 -99.815 94.105 ;
        RECT -95.765 93.935 -95.215 94.105 ;
        RECT -95.035 93.865 -94.665 94.205 ;
        RECT -94.485 94.105 -94.315 94.430 ;
        RECT -91.345 94.430 -90.275 94.600 ;
        RECT -91.345 94.105 -91.175 94.430 ;
        RECT -94.485 93.925 -93.555 94.105 ;
        RECT -92.105 93.925 -91.175 94.105 ;
        RECT -90.995 93.865 -90.625 94.205 ;
        RECT -90.445 94.105 -90.275 94.430 ;
        RECT -85.465 94.430 -84.395 94.600 ;
        RECT -85.465 94.105 -85.295 94.430 ;
        RECT -90.445 93.935 -89.895 94.105 ;
        RECT -85.845 93.935 -85.295 94.105 ;
        RECT -85.115 93.865 -84.745 94.205 ;
        RECT -84.565 94.105 -84.395 94.430 ;
        RECT -81.425 94.430 -80.355 94.600 ;
        RECT -81.425 94.105 -81.255 94.430 ;
        RECT -84.565 93.925 -83.635 94.105 ;
        RECT -82.185 93.925 -81.255 94.105 ;
        RECT -81.075 93.865 -80.705 94.205 ;
        RECT -80.525 94.105 -80.355 94.430 ;
        RECT -75.545 94.430 -74.475 94.600 ;
        RECT -75.545 94.105 -75.375 94.430 ;
        RECT -80.525 93.935 -79.975 94.105 ;
        RECT -75.925 93.935 -75.375 94.105 ;
        RECT -75.195 93.865 -74.825 94.205 ;
        RECT -74.645 94.105 -74.475 94.430 ;
        RECT -71.505 94.430 -70.435 94.600 ;
        RECT -71.505 94.105 -71.335 94.430 ;
        RECT -74.645 93.925 -73.715 94.105 ;
        RECT -72.265 93.925 -71.335 94.105 ;
        RECT -71.155 93.865 -70.785 94.205 ;
        RECT -70.605 94.105 -70.435 94.430 ;
        RECT -65.625 94.430 -64.555 94.600 ;
        RECT -65.625 94.105 -65.455 94.430 ;
        RECT -70.605 93.935 -70.055 94.105 ;
        RECT -66.005 93.935 -65.455 94.105 ;
        RECT -65.275 93.865 -64.905 94.205 ;
        RECT -64.725 94.105 -64.555 94.430 ;
        RECT -61.585 94.430 -60.515 94.600 ;
        RECT -61.585 94.105 -61.415 94.430 ;
        RECT -64.725 93.925 -63.795 94.105 ;
        RECT -62.345 93.925 -61.415 94.105 ;
        RECT -61.235 93.865 -60.865 94.205 ;
        RECT -60.685 94.105 -60.515 94.430 ;
        RECT -55.705 94.430 -54.635 94.600 ;
        RECT -55.705 94.105 -55.535 94.430 ;
        RECT -60.685 93.935 -60.135 94.105 ;
        RECT -56.085 93.935 -55.535 94.105 ;
        RECT -55.355 93.865 -54.985 94.205 ;
        RECT -54.805 94.105 -54.635 94.430 ;
        RECT -51.665 94.430 -50.595 94.600 ;
        RECT -51.665 94.105 -51.495 94.430 ;
        RECT -54.805 93.925 -53.875 94.105 ;
        RECT -52.425 93.925 -51.495 94.105 ;
        RECT -51.315 93.865 -50.945 94.205 ;
        RECT -50.765 94.105 -50.595 94.430 ;
        RECT -45.785 94.430 -44.715 94.600 ;
        RECT -45.785 94.105 -45.615 94.430 ;
        RECT -50.765 93.935 -50.215 94.105 ;
        RECT -46.165 93.935 -45.615 94.105 ;
        RECT -45.435 93.865 -45.065 94.205 ;
        RECT -44.885 94.105 -44.715 94.430 ;
        RECT -41.745 94.430 -40.675 94.600 ;
        RECT -41.745 94.105 -41.575 94.430 ;
        RECT -44.885 93.925 -43.955 94.105 ;
        RECT -42.505 93.925 -41.575 94.105 ;
        RECT -41.395 93.865 -41.025 94.205 ;
        RECT -40.845 94.105 -40.675 94.430 ;
        RECT -35.865 94.430 -34.795 94.600 ;
        RECT -35.865 94.105 -35.695 94.430 ;
        RECT -40.845 93.935 -40.295 94.105 ;
        RECT -36.245 93.935 -35.695 94.105 ;
        RECT -35.515 93.865 -35.145 94.205 ;
        RECT -34.965 94.105 -34.795 94.430 ;
        RECT -31.825 94.430 -30.755 94.600 ;
        RECT -31.825 94.105 -31.655 94.430 ;
        RECT -34.965 93.925 -34.035 94.105 ;
        RECT -32.585 93.925 -31.655 94.105 ;
        RECT -31.475 93.865 -31.105 94.205 ;
        RECT -30.925 94.105 -30.755 94.430 ;
        RECT -25.945 94.430 -24.875 94.600 ;
        RECT -25.945 94.105 -25.775 94.430 ;
        RECT -30.925 93.935 -30.375 94.105 ;
        RECT -26.325 93.935 -25.775 94.105 ;
        RECT -25.595 93.865 -25.225 94.205 ;
        RECT -25.045 94.105 -24.875 94.430 ;
        RECT -21.905 94.430 -20.835 94.600 ;
        RECT -21.905 94.105 -21.735 94.430 ;
        RECT -25.045 93.925 -24.115 94.105 ;
        RECT -22.665 93.925 -21.735 94.105 ;
        RECT -21.555 93.865 -21.185 94.205 ;
        RECT -21.005 94.105 -20.835 94.430 ;
        RECT -16.025 94.430 -14.955 94.600 ;
        RECT -16.025 94.105 -15.855 94.430 ;
        RECT -21.005 93.935 -20.455 94.105 ;
        RECT -16.405 93.935 -15.855 94.105 ;
        RECT -15.675 93.865 -15.305 94.205 ;
        RECT -15.125 94.105 -14.955 94.430 ;
        RECT -11.985 94.430 -10.915 94.600 ;
        RECT -11.985 94.105 -11.815 94.430 ;
        RECT -15.125 93.925 -14.195 94.105 ;
        RECT -12.745 93.925 -11.815 94.105 ;
        RECT -11.635 93.865 -11.265 94.205 ;
        RECT -11.085 94.105 -10.915 94.430 ;
        RECT -6.105 94.430 -5.035 94.600 ;
        RECT -6.105 94.105 -5.935 94.430 ;
        RECT -11.085 93.935 -10.535 94.105 ;
        RECT -6.485 93.935 -5.935 94.105 ;
        RECT -5.755 93.865 -5.385 94.205 ;
        RECT -5.205 94.105 -5.035 94.430 ;
        RECT -2.065 94.430 -0.995 94.600 ;
        RECT -2.065 94.105 -1.895 94.430 ;
        RECT -5.205 93.925 -4.275 94.105 ;
        RECT -2.825 93.925 -1.895 94.105 ;
        RECT -1.715 93.865 -1.345 94.205 ;
        RECT -1.165 94.105 -0.995 94.430 ;
        RECT 3.815 94.430 4.885 94.600 ;
        RECT 3.815 94.105 3.985 94.430 ;
        RECT -1.165 93.935 -0.615 94.105 ;
        RECT 3.435 93.935 3.985 94.105 ;
        RECT 4.165 93.865 4.535 94.205 ;
        RECT 4.715 94.105 4.885 94.430 ;
        RECT 7.855 94.430 8.925 94.600 ;
        RECT 7.855 94.105 8.025 94.430 ;
        RECT 4.715 93.925 5.645 94.105 ;
        RECT 7.095 93.925 8.025 94.105 ;
        RECT 8.205 93.865 8.575 94.205 ;
        RECT 8.755 94.105 8.925 94.430 ;
        RECT 13.735 94.430 14.805 94.600 ;
        RECT 13.735 94.105 13.905 94.430 ;
        RECT 8.755 93.935 9.305 94.105 ;
        RECT 13.355 93.935 13.905 94.105 ;
        RECT 14.085 93.865 14.455 94.205 ;
        RECT 14.635 94.105 14.805 94.430 ;
        RECT 17.775 94.430 18.845 94.600 ;
        RECT 17.775 94.105 17.945 94.430 ;
        RECT 14.635 93.925 15.565 94.105 ;
        RECT 17.015 93.925 17.945 94.105 ;
        RECT 18.125 93.865 18.495 94.205 ;
        RECT 18.675 94.105 18.845 94.430 ;
        RECT 23.655 94.430 24.725 94.600 ;
        RECT 23.655 94.105 23.825 94.430 ;
        RECT 18.675 93.935 19.225 94.105 ;
        RECT 23.275 93.935 23.825 94.105 ;
        RECT 24.005 93.865 24.375 94.205 ;
        RECT 24.555 94.105 24.725 94.430 ;
        RECT 24.555 93.925 25.485 94.105 ;
        RECT -291.460 93.245 -289.620 93.415 ;
        RECT 24.600 93.245 26.440 93.415 ;
        RECT -291.375 92.520 -291.085 93.245 ;
        RECT -290.915 92.445 -290.605 93.245 ;
        RECT -290.400 92.445 -289.705 93.075 ;
        RECT -291.375 90.695 -291.085 91.860 ;
        RECT -290.400 91.845 -290.230 92.445 ;
        RECT -290.060 92.005 -289.725 92.255 ;
        RECT -287.365 92.095 -287.035 93.075 ;
        RECT -285.505 92.095 -285.175 93.075 ;
        RECT -282.835 92.445 -282.140 93.075 ;
        RECT -290.915 90.695 -290.635 91.835 ;
        RECT -290.465 90.865 -290.135 91.845 ;
        RECT -289.965 90.695 -289.705 91.835 ;
        RECT -287.775 91.685 -287.440 91.935 ;
        RECT -287.270 91.495 -287.100 92.095 ;
        RECT -287.795 90.865 -287.100 91.495 ;
        RECT -285.440 91.495 -285.270 92.095 ;
        RECT -282.815 92.005 -282.480 92.255 ;
        RECT -285.100 91.685 -284.765 91.935 ;
        RECT -282.310 91.845 -282.140 92.445 ;
        RECT -280.480 92.445 -279.785 93.075 ;
        RECT -280.480 91.845 -280.310 92.445 ;
        RECT -280.140 92.005 -279.805 92.255 ;
        RECT -277.445 92.095 -277.115 93.075 ;
        RECT -275.585 92.095 -275.255 93.075 ;
        RECT -272.915 92.445 -272.220 93.075 ;
        RECT -285.440 90.865 -284.745 91.495 ;
        RECT -282.405 90.865 -282.075 91.845 ;
        RECT -280.545 90.865 -280.215 91.845 ;
        RECT -277.855 91.685 -277.520 91.935 ;
        RECT -277.350 91.495 -277.180 92.095 ;
        RECT -277.875 90.865 -277.180 91.495 ;
        RECT -275.520 91.495 -275.350 92.095 ;
        RECT -272.895 92.005 -272.560 92.255 ;
        RECT -275.180 91.685 -274.845 91.935 ;
        RECT -272.390 91.845 -272.220 92.445 ;
        RECT -270.560 92.445 -269.865 93.075 ;
        RECT -270.560 91.845 -270.390 92.445 ;
        RECT -270.220 92.005 -269.885 92.255 ;
        RECT -267.525 92.095 -267.195 93.075 ;
        RECT -265.665 92.095 -265.335 93.075 ;
        RECT -262.995 92.445 -262.300 93.075 ;
        RECT -275.520 90.865 -274.825 91.495 ;
        RECT -272.485 90.865 -272.155 91.845 ;
        RECT -270.625 90.865 -270.295 91.845 ;
        RECT -267.935 91.685 -267.600 91.935 ;
        RECT -267.430 91.495 -267.260 92.095 ;
        RECT -267.955 90.865 -267.260 91.495 ;
        RECT -265.600 91.495 -265.430 92.095 ;
        RECT -262.975 92.005 -262.640 92.255 ;
        RECT -265.260 91.685 -264.925 91.935 ;
        RECT -262.470 91.845 -262.300 92.445 ;
        RECT -260.640 92.445 -259.945 93.075 ;
        RECT -260.640 91.845 -260.470 92.445 ;
        RECT -260.300 92.005 -259.965 92.255 ;
        RECT -257.605 92.095 -257.275 93.075 ;
        RECT -255.745 92.095 -255.415 93.075 ;
        RECT -253.075 92.445 -252.380 93.075 ;
        RECT -265.600 90.865 -264.905 91.495 ;
        RECT -262.565 90.865 -262.235 91.845 ;
        RECT -260.705 90.865 -260.375 91.845 ;
        RECT -258.015 91.685 -257.680 91.935 ;
        RECT -257.510 91.495 -257.340 92.095 ;
        RECT -258.035 90.865 -257.340 91.495 ;
        RECT -255.680 91.495 -255.510 92.095 ;
        RECT -253.055 92.005 -252.720 92.255 ;
        RECT -255.340 91.685 -255.005 91.935 ;
        RECT -252.550 91.845 -252.380 92.445 ;
        RECT -250.720 92.445 -250.025 93.075 ;
        RECT -250.720 91.845 -250.550 92.445 ;
        RECT -250.380 92.005 -250.045 92.255 ;
        RECT -247.685 92.095 -247.355 93.075 ;
        RECT -245.825 92.095 -245.495 93.075 ;
        RECT -243.155 92.445 -242.460 93.075 ;
        RECT -255.680 90.865 -254.985 91.495 ;
        RECT -252.645 90.865 -252.315 91.845 ;
        RECT -250.785 90.865 -250.455 91.845 ;
        RECT -248.095 91.685 -247.760 91.935 ;
        RECT -247.590 91.495 -247.420 92.095 ;
        RECT -248.115 90.865 -247.420 91.495 ;
        RECT -245.760 91.495 -245.590 92.095 ;
        RECT -243.135 92.005 -242.800 92.255 ;
        RECT -245.420 91.685 -245.085 91.935 ;
        RECT -242.630 91.845 -242.460 92.445 ;
        RECT -240.800 92.445 -240.105 93.075 ;
        RECT -240.800 91.845 -240.630 92.445 ;
        RECT -240.460 92.005 -240.125 92.255 ;
        RECT -237.765 92.095 -237.435 93.075 ;
        RECT -235.905 92.095 -235.575 93.075 ;
        RECT -233.235 92.445 -232.540 93.075 ;
        RECT -245.760 90.865 -245.065 91.495 ;
        RECT -242.725 90.865 -242.395 91.845 ;
        RECT -240.865 90.865 -240.535 91.845 ;
        RECT -238.175 91.685 -237.840 91.935 ;
        RECT -237.670 91.495 -237.500 92.095 ;
        RECT -238.195 90.865 -237.500 91.495 ;
        RECT -235.840 91.495 -235.670 92.095 ;
        RECT -233.215 92.005 -232.880 92.255 ;
        RECT -235.500 91.685 -235.165 91.935 ;
        RECT -232.710 91.845 -232.540 92.445 ;
        RECT -230.880 92.445 -230.185 93.075 ;
        RECT -230.880 91.845 -230.710 92.445 ;
        RECT -230.540 92.005 -230.205 92.255 ;
        RECT -227.845 92.095 -227.515 93.075 ;
        RECT -225.985 92.095 -225.655 93.075 ;
        RECT -223.315 92.445 -222.620 93.075 ;
        RECT -235.840 90.865 -235.145 91.495 ;
        RECT -232.805 90.865 -232.475 91.845 ;
        RECT -230.945 90.865 -230.615 91.845 ;
        RECT -228.255 91.685 -227.920 91.935 ;
        RECT -227.750 91.495 -227.580 92.095 ;
        RECT -228.275 90.865 -227.580 91.495 ;
        RECT -225.920 91.495 -225.750 92.095 ;
        RECT -223.295 92.005 -222.960 92.255 ;
        RECT -225.580 91.685 -225.245 91.935 ;
        RECT -222.790 91.845 -222.620 92.445 ;
        RECT -220.960 92.445 -220.265 93.075 ;
        RECT -220.960 91.845 -220.790 92.445 ;
        RECT -220.620 92.005 -220.285 92.255 ;
        RECT -217.925 92.095 -217.595 93.075 ;
        RECT -216.065 92.095 -215.735 93.075 ;
        RECT -213.395 92.445 -212.700 93.075 ;
        RECT -225.920 90.865 -225.225 91.495 ;
        RECT -222.885 90.865 -222.555 91.845 ;
        RECT -221.025 90.865 -220.695 91.845 ;
        RECT -218.335 91.685 -218.000 91.935 ;
        RECT -217.830 91.495 -217.660 92.095 ;
        RECT -218.355 90.865 -217.660 91.495 ;
        RECT -216.000 91.495 -215.830 92.095 ;
        RECT -213.375 92.005 -213.040 92.255 ;
        RECT -215.660 91.685 -215.325 91.935 ;
        RECT -212.870 91.845 -212.700 92.445 ;
        RECT -211.040 92.445 -210.345 93.075 ;
        RECT -211.040 91.845 -210.870 92.445 ;
        RECT -210.700 92.005 -210.365 92.255 ;
        RECT -208.005 92.095 -207.675 93.075 ;
        RECT -206.145 92.095 -205.815 93.075 ;
        RECT -203.475 92.445 -202.780 93.075 ;
        RECT -216.000 90.865 -215.305 91.495 ;
        RECT -212.965 90.865 -212.635 91.845 ;
        RECT -211.105 90.865 -210.775 91.845 ;
        RECT -208.415 91.685 -208.080 91.935 ;
        RECT -207.910 91.495 -207.740 92.095 ;
        RECT -208.435 90.865 -207.740 91.495 ;
        RECT -206.080 91.495 -205.910 92.095 ;
        RECT -203.455 92.005 -203.120 92.255 ;
        RECT -205.740 91.685 -205.405 91.935 ;
        RECT -202.950 91.845 -202.780 92.445 ;
        RECT -201.120 92.445 -200.425 93.075 ;
        RECT -201.120 91.845 -200.950 92.445 ;
        RECT -200.780 92.005 -200.445 92.255 ;
        RECT -198.085 92.095 -197.755 93.075 ;
        RECT -196.225 92.095 -195.895 93.075 ;
        RECT -193.555 92.445 -192.860 93.075 ;
        RECT -206.080 90.865 -205.385 91.495 ;
        RECT -203.045 90.865 -202.715 91.845 ;
        RECT -201.185 90.865 -200.855 91.845 ;
        RECT -198.495 91.685 -198.160 91.935 ;
        RECT -197.990 91.495 -197.820 92.095 ;
        RECT -198.515 90.865 -197.820 91.495 ;
        RECT -196.160 91.495 -195.990 92.095 ;
        RECT -193.535 92.005 -193.200 92.255 ;
        RECT -195.820 91.685 -195.485 91.935 ;
        RECT -193.030 91.845 -192.860 92.445 ;
        RECT -191.200 92.445 -190.505 93.075 ;
        RECT -191.200 91.845 -191.030 92.445 ;
        RECT -190.860 92.005 -190.525 92.255 ;
        RECT -188.165 92.095 -187.835 93.075 ;
        RECT -186.305 92.095 -185.975 93.075 ;
        RECT -183.635 92.445 -182.940 93.075 ;
        RECT -196.160 90.865 -195.465 91.495 ;
        RECT -193.125 90.865 -192.795 91.845 ;
        RECT -191.265 90.865 -190.935 91.845 ;
        RECT -188.575 91.685 -188.240 91.935 ;
        RECT -188.070 91.495 -187.900 92.095 ;
        RECT -188.595 90.865 -187.900 91.495 ;
        RECT -186.240 91.495 -186.070 92.095 ;
        RECT -183.615 92.005 -183.280 92.255 ;
        RECT -185.900 91.685 -185.565 91.935 ;
        RECT -183.110 91.845 -182.940 92.445 ;
        RECT -181.280 92.445 -180.585 93.075 ;
        RECT -181.280 91.845 -181.110 92.445 ;
        RECT -180.940 92.005 -180.605 92.255 ;
        RECT -178.245 92.095 -177.915 93.075 ;
        RECT -176.385 92.095 -176.055 93.075 ;
        RECT -173.715 92.445 -173.020 93.075 ;
        RECT -186.240 90.865 -185.545 91.495 ;
        RECT -183.205 90.865 -182.875 91.845 ;
        RECT -181.345 90.865 -181.015 91.845 ;
        RECT -178.655 91.685 -178.320 91.935 ;
        RECT -178.150 91.495 -177.980 92.095 ;
        RECT -178.675 90.865 -177.980 91.495 ;
        RECT -176.320 91.495 -176.150 92.095 ;
        RECT -173.695 92.005 -173.360 92.255 ;
        RECT -175.980 91.685 -175.645 91.935 ;
        RECT -173.190 91.845 -173.020 92.445 ;
        RECT -171.360 92.445 -170.665 93.075 ;
        RECT -171.360 91.845 -171.190 92.445 ;
        RECT -171.020 92.005 -170.685 92.255 ;
        RECT -168.325 92.095 -167.995 93.075 ;
        RECT -166.465 92.095 -166.135 93.075 ;
        RECT -163.795 92.445 -163.100 93.075 ;
        RECT -176.320 90.865 -175.625 91.495 ;
        RECT -173.285 90.865 -172.955 91.845 ;
        RECT -171.425 90.865 -171.095 91.845 ;
        RECT -168.735 91.685 -168.400 91.935 ;
        RECT -168.230 91.495 -168.060 92.095 ;
        RECT -168.755 90.865 -168.060 91.495 ;
        RECT -166.400 91.495 -166.230 92.095 ;
        RECT -163.775 92.005 -163.440 92.255 ;
        RECT -166.060 91.685 -165.725 91.935 ;
        RECT -163.270 91.845 -163.100 92.445 ;
        RECT -161.440 92.445 -160.745 93.075 ;
        RECT -161.440 91.845 -161.270 92.445 ;
        RECT -161.100 92.005 -160.765 92.255 ;
        RECT -158.405 92.095 -158.075 93.075 ;
        RECT -156.545 92.095 -156.215 93.075 ;
        RECT -153.875 92.445 -153.180 93.075 ;
        RECT -166.400 90.865 -165.705 91.495 ;
        RECT -163.365 90.865 -163.035 91.845 ;
        RECT -161.505 90.865 -161.175 91.845 ;
        RECT -158.815 91.685 -158.480 91.935 ;
        RECT -158.310 91.495 -158.140 92.095 ;
        RECT -158.835 90.865 -158.140 91.495 ;
        RECT -156.480 91.495 -156.310 92.095 ;
        RECT -153.855 92.005 -153.520 92.255 ;
        RECT -156.140 91.685 -155.805 91.935 ;
        RECT -153.350 91.845 -153.180 92.445 ;
        RECT -151.520 92.445 -150.825 93.075 ;
        RECT -151.520 91.845 -151.350 92.445 ;
        RECT -151.180 92.005 -150.845 92.255 ;
        RECT -148.485 92.095 -148.155 93.075 ;
        RECT -146.625 92.095 -146.295 93.075 ;
        RECT -143.955 92.445 -143.260 93.075 ;
        RECT -156.480 90.865 -155.785 91.495 ;
        RECT -153.445 90.865 -153.115 91.845 ;
        RECT -151.585 90.865 -151.255 91.845 ;
        RECT -148.895 91.685 -148.560 91.935 ;
        RECT -148.390 91.495 -148.220 92.095 ;
        RECT -148.915 90.865 -148.220 91.495 ;
        RECT -146.560 91.495 -146.390 92.095 ;
        RECT -143.935 92.005 -143.600 92.255 ;
        RECT -146.220 91.685 -145.885 91.935 ;
        RECT -143.430 91.845 -143.260 92.445 ;
        RECT -141.600 92.445 -140.905 93.075 ;
        RECT -141.600 91.845 -141.430 92.445 ;
        RECT -141.260 92.005 -140.925 92.255 ;
        RECT -138.565 92.095 -138.235 93.075 ;
        RECT -136.705 92.095 -136.375 93.075 ;
        RECT -134.035 92.445 -133.340 93.075 ;
        RECT -146.560 90.865 -145.865 91.495 ;
        RECT -143.525 90.865 -143.195 91.845 ;
        RECT -141.665 90.865 -141.335 91.845 ;
        RECT -138.975 91.685 -138.640 91.935 ;
        RECT -138.470 91.495 -138.300 92.095 ;
        RECT -138.995 90.865 -138.300 91.495 ;
        RECT -136.640 91.495 -136.470 92.095 ;
        RECT -134.015 92.005 -133.680 92.255 ;
        RECT -136.300 91.685 -135.965 91.935 ;
        RECT -133.510 91.845 -133.340 92.445 ;
        RECT -131.680 92.445 -130.985 93.075 ;
        RECT -131.680 91.845 -131.510 92.445 ;
        RECT -131.340 92.005 -131.005 92.255 ;
        RECT -128.645 92.095 -128.315 93.075 ;
        RECT -126.785 92.095 -126.455 93.075 ;
        RECT -124.115 92.445 -123.420 93.075 ;
        RECT -136.640 90.865 -135.945 91.495 ;
        RECT -133.605 90.865 -133.275 91.845 ;
        RECT -131.745 90.865 -131.415 91.845 ;
        RECT -129.055 91.685 -128.720 91.935 ;
        RECT -128.550 91.495 -128.380 92.095 ;
        RECT -129.075 90.865 -128.380 91.495 ;
        RECT -126.720 91.495 -126.550 92.095 ;
        RECT -124.095 92.005 -123.760 92.255 ;
        RECT -126.380 91.685 -126.045 91.935 ;
        RECT -123.590 91.845 -123.420 92.445 ;
        RECT -121.760 92.445 -121.065 93.075 ;
        RECT -121.760 91.845 -121.590 92.445 ;
        RECT -121.420 92.005 -121.085 92.255 ;
        RECT -118.725 92.095 -118.395 93.075 ;
        RECT -116.865 92.095 -116.535 93.075 ;
        RECT -114.195 92.445 -113.500 93.075 ;
        RECT -126.720 90.865 -126.025 91.495 ;
        RECT -123.685 90.865 -123.355 91.845 ;
        RECT -121.825 90.865 -121.495 91.845 ;
        RECT -119.135 91.685 -118.800 91.935 ;
        RECT -118.630 91.495 -118.460 92.095 ;
        RECT -119.155 90.865 -118.460 91.495 ;
        RECT -116.800 91.495 -116.630 92.095 ;
        RECT -114.175 92.005 -113.840 92.255 ;
        RECT -116.460 91.685 -116.125 91.935 ;
        RECT -113.670 91.845 -113.500 92.445 ;
        RECT -111.840 92.445 -111.145 93.075 ;
        RECT -111.840 91.845 -111.670 92.445 ;
        RECT -111.500 92.005 -111.165 92.255 ;
        RECT -108.805 92.095 -108.475 93.075 ;
        RECT -106.945 92.095 -106.615 93.075 ;
        RECT -104.275 92.445 -103.580 93.075 ;
        RECT -116.800 90.865 -116.105 91.495 ;
        RECT -113.765 90.865 -113.435 91.845 ;
        RECT -111.905 90.865 -111.575 91.845 ;
        RECT -109.215 91.685 -108.880 91.935 ;
        RECT -108.710 91.495 -108.540 92.095 ;
        RECT -109.235 90.865 -108.540 91.495 ;
        RECT -106.880 91.495 -106.710 92.095 ;
        RECT -104.255 92.005 -103.920 92.255 ;
        RECT -106.540 91.685 -106.205 91.935 ;
        RECT -103.750 91.845 -103.580 92.445 ;
        RECT -101.920 92.445 -101.225 93.075 ;
        RECT -101.920 91.845 -101.750 92.445 ;
        RECT -101.580 92.005 -101.245 92.255 ;
        RECT -98.885 92.095 -98.555 93.075 ;
        RECT -97.025 92.095 -96.695 93.075 ;
        RECT -94.355 92.445 -93.660 93.075 ;
        RECT -106.880 90.865 -106.185 91.495 ;
        RECT -103.845 90.865 -103.515 91.845 ;
        RECT -101.985 90.865 -101.655 91.845 ;
        RECT -99.295 91.685 -98.960 91.935 ;
        RECT -98.790 91.495 -98.620 92.095 ;
        RECT -99.315 90.865 -98.620 91.495 ;
        RECT -96.960 91.495 -96.790 92.095 ;
        RECT -94.335 92.005 -94.000 92.255 ;
        RECT -96.620 91.685 -96.285 91.935 ;
        RECT -93.830 91.845 -93.660 92.445 ;
        RECT -92.000 92.445 -91.305 93.075 ;
        RECT -92.000 91.845 -91.830 92.445 ;
        RECT -91.660 92.005 -91.325 92.255 ;
        RECT -88.965 92.095 -88.635 93.075 ;
        RECT -87.105 92.095 -86.775 93.075 ;
        RECT -84.435 92.445 -83.740 93.075 ;
        RECT -96.960 90.865 -96.265 91.495 ;
        RECT -93.925 90.865 -93.595 91.845 ;
        RECT -92.065 90.865 -91.735 91.845 ;
        RECT -89.375 91.685 -89.040 91.935 ;
        RECT -88.870 91.495 -88.700 92.095 ;
        RECT -89.395 90.865 -88.700 91.495 ;
        RECT -87.040 91.495 -86.870 92.095 ;
        RECT -84.415 92.005 -84.080 92.255 ;
        RECT -86.700 91.685 -86.365 91.935 ;
        RECT -83.910 91.845 -83.740 92.445 ;
        RECT -82.080 92.445 -81.385 93.075 ;
        RECT -82.080 91.845 -81.910 92.445 ;
        RECT -81.740 92.005 -81.405 92.255 ;
        RECT -79.045 92.095 -78.715 93.075 ;
        RECT -77.185 92.095 -76.855 93.075 ;
        RECT -74.515 92.445 -73.820 93.075 ;
        RECT -87.040 90.865 -86.345 91.495 ;
        RECT -84.005 90.865 -83.675 91.845 ;
        RECT -82.145 90.865 -81.815 91.845 ;
        RECT -79.455 91.685 -79.120 91.935 ;
        RECT -78.950 91.495 -78.780 92.095 ;
        RECT -79.475 90.865 -78.780 91.495 ;
        RECT -77.120 91.495 -76.950 92.095 ;
        RECT -74.495 92.005 -74.160 92.255 ;
        RECT -76.780 91.685 -76.445 91.935 ;
        RECT -73.990 91.845 -73.820 92.445 ;
        RECT -72.160 92.445 -71.465 93.075 ;
        RECT -72.160 91.845 -71.990 92.445 ;
        RECT -71.820 92.005 -71.485 92.255 ;
        RECT -69.125 92.095 -68.795 93.075 ;
        RECT -67.265 92.095 -66.935 93.075 ;
        RECT -64.595 92.445 -63.900 93.075 ;
        RECT -77.120 90.865 -76.425 91.495 ;
        RECT -74.085 90.865 -73.755 91.845 ;
        RECT -72.225 90.865 -71.895 91.845 ;
        RECT -69.535 91.685 -69.200 91.935 ;
        RECT -69.030 91.495 -68.860 92.095 ;
        RECT -69.555 90.865 -68.860 91.495 ;
        RECT -67.200 91.495 -67.030 92.095 ;
        RECT -64.575 92.005 -64.240 92.255 ;
        RECT -66.860 91.685 -66.525 91.935 ;
        RECT -64.070 91.845 -63.900 92.445 ;
        RECT -62.240 92.445 -61.545 93.075 ;
        RECT -62.240 91.845 -62.070 92.445 ;
        RECT -61.900 92.005 -61.565 92.255 ;
        RECT -59.205 92.095 -58.875 93.075 ;
        RECT -57.345 92.095 -57.015 93.075 ;
        RECT -54.675 92.445 -53.980 93.075 ;
        RECT -67.200 90.865 -66.505 91.495 ;
        RECT -64.165 90.865 -63.835 91.845 ;
        RECT -62.305 90.865 -61.975 91.845 ;
        RECT -59.615 91.685 -59.280 91.935 ;
        RECT -59.110 91.495 -58.940 92.095 ;
        RECT -59.635 90.865 -58.940 91.495 ;
        RECT -57.280 91.495 -57.110 92.095 ;
        RECT -54.655 92.005 -54.320 92.255 ;
        RECT -56.940 91.685 -56.605 91.935 ;
        RECT -54.150 91.845 -53.980 92.445 ;
        RECT -52.320 92.445 -51.625 93.075 ;
        RECT -52.320 91.845 -52.150 92.445 ;
        RECT -51.980 92.005 -51.645 92.255 ;
        RECT -49.285 92.095 -48.955 93.075 ;
        RECT -47.425 92.095 -47.095 93.075 ;
        RECT -44.755 92.445 -44.060 93.075 ;
        RECT -57.280 90.865 -56.585 91.495 ;
        RECT -54.245 90.865 -53.915 91.845 ;
        RECT -52.385 90.865 -52.055 91.845 ;
        RECT -49.695 91.685 -49.360 91.935 ;
        RECT -49.190 91.495 -49.020 92.095 ;
        RECT -49.715 90.865 -49.020 91.495 ;
        RECT -47.360 91.495 -47.190 92.095 ;
        RECT -44.735 92.005 -44.400 92.255 ;
        RECT -47.020 91.685 -46.685 91.935 ;
        RECT -44.230 91.845 -44.060 92.445 ;
        RECT -42.400 92.445 -41.705 93.075 ;
        RECT -42.400 91.845 -42.230 92.445 ;
        RECT -42.060 92.005 -41.725 92.255 ;
        RECT -39.365 92.095 -39.035 93.075 ;
        RECT -37.505 92.095 -37.175 93.075 ;
        RECT -34.835 92.445 -34.140 93.075 ;
        RECT -47.360 90.865 -46.665 91.495 ;
        RECT -44.325 90.865 -43.995 91.845 ;
        RECT -42.465 90.865 -42.135 91.845 ;
        RECT -39.775 91.685 -39.440 91.935 ;
        RECT -39.270 91.495 -39.100 92.095 ;
        RECT -39.795 90.865 -39.100 91.495 ;
        RECT -37.440 91.495 -37.270 92.095 ;
        RECT -34.815 92.005 -34.480 92.255 ;
        RECT -37.100 91.685 -36.765 91.935 ;
        RECT -34.310 91.845 -34.140 92.445 ;
        RECT -32.480 92.445 -31.785 93.075 ;
        RECT -32.480 91.845 -32.310 92.445 ;
        RECT -32.140 92.005 -31.805 92.255 ;
        RECT -29.445 92.095 -29.115 93.075 ;
        RECT -27.585 92.095 -27.255 93.075 ;
        RECT -24.915 92.445 -24.220 93.075 ;
        RECT -37.440 90.865 -36.745 91.495 ;
        RECT -34.405 90.865 -34.075 91.845 ;
        RECT -32.545 90.865 -32.215 91.845 ;
        RECT -29.855 91.685 -29.520 91.935 ;
        RECT -29.350 91.495 -29.180 92.095 ;
        RECT -29.875 90.865 -29.180 91.495 ;
        RECT -27.520 91.495 -27.350 92.095 ;
        RECT -24.895 92.005 -24.560 92.255 ;
        RECT -27.180 91.685 -26.845 91.935 ;
        RECT -24.390 91.845 -24.220 92.445 ;
        RECT -22.560 92.445 -21.865 93.075 ;
        RECT -22.560 91.845 -22.390 92.445 ;
        RECT -22.220 92.005 -21.885 92.255 ;
        RECT -19.525 92.095 -19.195 93.075 ;
        RECT -17.665 92.095 -17.335 93.075 ;
        RECT -14.995 92.445 -14.300 93.075 ;
        RECT -27.520 90.865 -26.825 91.495 ;
        RECT -24.485 90.865 -24.155 91.845 ;
        RECT -22.625 90.865 -22.295 91.845 ;
        RECT -19.935 91.685 -19.600 91.935 ;
        RECT -19.430 91.495 -19.260 92.095 ;
        RECT -19.955 90.865 -19.260 91.495 ;
        RECT -17.600 91.495 -17.430 92.095 ;
        RECT -14.975 92.005 -14.640 92.255 ;
        RECT -17.260 91.685 -16.925 91.935 ;
        RECT -14.470 91.845 -14.300 92.445 ;
        RECT -12.640 92.445 -11.945 93.075 ;
        RECT -12.640 91.845 -12.470 92.445 ;
        RECT -12.300 92.005 -11.965 92.255 ;
        RECT -9.605 92.095 -9.275 93.075 ;
        RECT -7.745 92.095 -7.415 93.075 ;
        RECT -5.075 92.445 -4.380 93.075 ;
        RECT -17.600 90.865 -16.905 91.495 ;
        RECT -14.565 90.865 -14.235 91.845 ;
        RECT -12.705 90.865 -12.375 91.845 ;
        RECT -10.015 91.685 -9.680 91.935 ;
        RECT -9.510 91.495 -9.340 92.095 ;
        RECT -10.035 90.865 -9.340 91.495 ;
        RECT -7.680 91.495 -7.510 92.095 ;
        RECT -5.055 92.005 -4.720 92.255 ;
        RECT -7.340 91.685 -7.005 91.935 ;
        RECT -4.550 91.845 -4.380 92.445 ;
        RECT -2.720 92.445 -2.025 93.075 ;
        RECT -2.720 91.845 -2.550 92.445 ;
        RECT -2.380 92.005 -2.045 92.255 ;
        RECT 0.315 92.095 0.645 93.075 ;
        RECT 2.175 92.095 2.505 93.075 ;
        RECT 4.845 92.445 5.540 93.075 ;
        RECT -7.680 90.865 -6.985 91.495 ;
        RECT -4.645 90.865 -4.315 91.845 ;
        RECT -2.785 90.865 -2.455 91.845 ;
        RECT -0.095 91.685 0.240 91.935 ;
        RECT 0.410 91.495 0.580 92.095 ;
        RECT -0.115 90.865 0.580 91.495 ;
        RECT 2.240 91.495 2.410 92.095 ;
        RECT 4.865 92.005 5.200 92.255 ;
        RECT 2.580 91.685 2.915 91.935 ;
        RECT 5.370 91.845 5.540 92.445 ;
        RECT 7.200 92.445 7.895 93.075 ;
        RECT 7.200 91.845 7.370 92.445 ;
        RECT 7.540 92.005 7.875 92.255 ;
        RECT 10.235 92.095 10.565 93.075 ;
        RECT 12.095 92.095 12.425 93.075 ;
        RECT 14.765 92.445 15.460 93.075 ;
        RECT 2.240 90.865 2.935 91.495 ;
        RECT 5.275 90.865 5.605 91.845 ;
        RECT 7.135 90.865 7.465 91.845 ;
        RECT 9.825 91.685 10.160 91.935 ;
        RECT 10.330 91.495 10.500 92.095 ;
        RECT 9.805 90.865 10.500 91.495 ;
        RECT 12.160 91.495 12.330 92.095 ;
        RECT 14.785 92.005 15.120 92.255 ;
        RECT 12.500 91.685 12.835 91.935 ;
        RECT 15.290 91.845 15.460 92.445 ;
        RECT 17.120 92.445 17.815 93.075 ;
        RECT 17.120 91.845 17.290 92.445 ;
        RECT 17.460 92.005 17.795 92.255 ;
        RECT 20.155 92.095 20.485 93.075 ;
        RECT 22.015 92.095 22.345 93.075 ;
        RECT 24.685 92.445 25.380 93.075 ;
        RECT 25.585 92.445 25.895 93.245 ;
        RECT 26.065 92.520 26.355 93.245 ;
        RECT 12.160 90.865 12.855 91.495 ;
        RECT 15.195 90.865 15.525 91.845 ;
        RECT 17.055 90.865 17.385 91.845 ;
        RECT 19.745 91.685 20.080 91.935 ;
        RECT 20.250 91.495 20.420 92.095 ;
        RECT 19.725 90.865 20.420 91.495 ;
        RECT 22.080 91.495 22.250 92.095 ;
        RECT 24.705 92.005 25.040 92.255 ;
        RECT 22.420 91.685 22.755 91.935 ;
        RECT 25.210 91.845 25.380 92.445 ;
        RECT 22.080 90.865 22.775 91.495 ;
        RECT 25.115 90.865 25.445 91.845 ;
        RECT -291.460 90.525 -289.620 90.695 ;
        RECT -290.075 89.140 -289.785 89.850 ;
        RECT -289.545 89.655 -289.375 90.180 ;
        RECT -289.205 89.835 -288.655 90.005 ;
        RECT -289.545 89.325 -288.995 89.655 ;
        RECT -288.825 89.510 -288.655 89.835 ;
        RECT -288.475 89.735 -288.105 90.075 ;
        RECT -287.925 89.835 -286.995 90.015 ;
        RECT -285.545 89.835 -284.615 90.015 ;
        RECT -287.925 89.510 -287.755 89.835 ;
        RECT -288.825 89.340 -287.755 89.510 ;
        RECT -284.785 89.510 -284.615 89.835 ;
        RECT -284.435 89.735 -284.065 90.075 ;
        RECT -283.885 89.835 -283.335 90.005 ;
        RECT -279.285 89.835 -278.735 90.005 ;
        RECT -283.885 89.510 -283.715 89.835 ;
        RECT -284.785 89.340 -283.715 89.510 ;
        RECT -278.905 89.510 -278.735 89.835 ;
        RECT -278.555 89.735 -278.185 90.075 ;
        RECT -278.005 89.835 -277.075 90.015 ;
        RECT -275.625 89.835 -274.695 90.015 ;
        RECT -278.005 89.510 -277.835 89.835 ;
        RECT -278.905 89.340 -277.835 89.510 ;
        RECT -274.865 89.510 -274.695 89.835 ;
        RECT -274.515 89.735 -274.145 90.075 ;
        RECT -273.965 89.835 -273.415 90.005 ;
        RECT -269.365 89.835 -268.815 90.005 ;
        RECT -273.965 89.510 -273.795 89.835 ;
        RECT -274.865 89.340 -273.795 89.510 ;
        RECT -268.985 89.510 -268.815 89.835 ;
        RECT -268.635 89.735 -268.265 90.075 ;
        RECT -268.085 89.835 -267.155 90.015 ;
        RECT -265.705 89.835 -264.775 90.015 ;
        RECT -268.085 89.510 -267.915 89.835 ;
        RECT -268.985 89.340 -267.915 89.510 ;
        RECT -264.945 89.510 -264.775 89.835 ;
        RECT -264.595 89.735 -264.225 90.075 ;
        RECT -264.045 89.835 -263.495 90.005 ;
        RECT -259.445 89.835 -258.895 90.005 ;
        RECT -264.045 89.510 -263.875 89.835 ;
        RECT -264.945 89.340 -263.875 89.510 ;
        RECT -259.065 89.510 -258.895 89.835 ;
        RECT -258.715 89.735 -258.345 90.075 ;
        RECT -258.165 89.835 -257.235 90.015 ;
        RECT -255.785 89.835 -254.855 90.015 ;
        RECT -258.165 89.510 -257.995 89.835 ;
        RECT -259.065 89.340 -257.995 89.510 ;
        RECT -255.025 89.510 -254.855 89.835 ;
        RECT -254.675 89.735 -254.305 90.075 ;
        RECT -254.125 89.835 -253.575 90.005 ;
        RECT -249.525 89.835 -248.975 90.005 ;
        RECT -254.125 89.510 -253.955 89.835 ;
        RECT -255.025 89.340 -253.955 89.510 ;
        RECT -249.145 89.510 -248.975 89.835 ;
        RECT -248.795 89.735 -248.425 90.075 ;
        RECT -248.245 89.835 -247.315 90.015 ;
        RECT -245.865 89.835 -244.935 90.015 ;
        RECT -248.245 89.510 -248.075 89.835 ;
        RECT -249.145 89.340 -248.075 89.510 ;
        RECT -245.105 89.510 -244.935 89.835 ;
        RECT -244.755 89.735 -244.385 90.075 ;
        RECT -244.205 89.835 -243.655 90.005 ;
        RECT -239.605 89.835 -239.055 90.005 ;
        RECT -244.205 89.510 -244.035 89.835 ;
        RECT -245.105 89.340 -244.035 89.510 ;
        RECT -239.225 89.510 -239.055 89.835 ;
        RECT -238.875 89.735 -238.505 90.075 ;
        RECT -238.325 89.835 -237.395 90.015 ;
        RECT -235.945 89.835 -235.015 90.015 ;
        RECT -238.325 89.510 -238.155 89.835 ;
        RECT -239.225 89.340 -238.155 89.510 ;
        RECT -235.185 89.510 -235.015 89.835 ;
        RECT -234.835 89.735 -234.465 90.075 ;
        RECT -234.285 89.835 -233.735 90.005 ;
        RECT -229.685 89.835 -229.135 90.005 ;
        RECT -234.285 89.510 -234.115 89.835 ;
        RECT -235.185 89.340 -234.115 89.510 ;
        RECT -229.305 89.510 -229.135 89.835 ;
        RECT -228.955 89.735 -228.585 90.075 ;
        RECT -228.405 89.835 -227.475 90.015 ;
        RECT -226.025 89.835 -225.095 90.015 ;
        RECT -228.405 89.510 -228.235 89.835 ;
        RECT -229.305 89.340 -228.235 89.510 ;
        RECT -225.265 89.510 -225.095 89.835 ;
        RECT -224.915 89.735 -224.545 90.075 ;
        RECT -224.365 89.835 -223.815 90.005 ;
        RECT -219.765 89.835 -219.215 90.005 ;
        RECT -224.365 89.510 -224.195 89.835 ;
        RECT -225.265 89.340 -224.195 89.510 ;
        RECT -219.385 89.510 -219.215 89.835 ;
        RECT -219.035 89.735 -218.665 90.075 ;
        RECT -218.485 89.835 -217.555 90.015 ;
        RECT -216.105 89.835 -215.175 90.015 ;
        RECT -218.485 89.510 -218.315 89.835 ;
        RECT -219.385 89.340 -218.315 89.510 ;
        RECT -215.345 89.510 -215.175 89.835 ;
        RECT -214.995 89.735 -214.625 90.075 ;
        RECT -214.445 89.835 -213.895 90.005 ;
        RECT -209.845 89.835 -209.295 90.005 ;
        RECT -214.445 89.510 -214.275 89.835 ;
        RECT -215.345 89.340 -214.275 89.510 ;
        RECT -209.465 89.510 -209.295 89.835 ;
        RECT -209.115 89.735 -208.745 90.075 ;
        RECT -208.565 89.835 -207.635 90.015 ;
        RECT -206.185 89.835 -205.255 90.015 ;
        RECT -208.565 89.510 -208.395 89.835 ;
        RECT -209.465 89.340 -208.395 89.510 ;
        RECT -205.425 89.510 -205.255 89.835 ;
        RECT -205.075 89.735 -204.705 90.075 ;
        RECT -204.525 89.835 -203.975 90.005 ;
        RECT -199.925 89.835 -199.375 90.005 ;
        RECT -204.525 89.510 -204.355 89.835 ;
        RECT -205.425 89.340 -204.355 89.510 ;
        RECT -199.545 89.510 -199.375 89.835 ;
        RECT -199.195 89.735 -198.825 90.075 ;
        RECT -198.645 89.835 -197.715 90.015 ;
        RECT -196.265 89.835 -195.335 90.015 ;
        RECT -198.645 89.510 -198.475 89.835 ;
        RECT -199.545 89.340 -198.475 89.510 ;
        RECT -195.505 89.510 -195.335 89.835 ;
        RECT -195.155 89.735 -194.785 90.075 ;
        RECT -194.605 89.835 -194.055 90.005 ;
        RECT -190.005 89.835 -189.455 90.005 ;
        RECT -194.605 89.510 -194.435 89.835 ;
        RECT -195.505 89.340 -194.435 89.510 ;
        RECT -189.625 89.510 -189.455 89.835 ;
        RECT -189.275 89.735 -188.905 90.075 ;
        RECT -188.725 89.835 -187.795 90.015 ;
        RECT -186.345 89.835 -185.415 90.015 ;
        RECT -188.725 89.510 -188.555 89.835 ;
        RECT -189.625 89.340 -188.555 89.510 ;
        RECT -185.585 89.510 -185.415 89.835 ;
        RECT -185.235 89.735 -184.865 90.075 ;
        RECT -184.685 89.835 -184.135 90.005 ;
        RECT -180.085 89.835 -179.535 90.005 ;
        RECT -184.685 89.510 -184.515 89.835 ;
        RECT -185.585 89.340 -184.515 89.510 ;
        RECT -179.705 89.510 -179.535 89.835 ;
        RECT -179.355 89.735 -178.985 90.075 ;
        RECT -178.805 89.835 -177.875 90.015 ;
        RECT -176.425 89.835 -175.495 90.015 ;
        RECT -178.805 89.510 -178.635 89.835 ;
        RECT -179.705 89.340 -178.635 89.510 ;
        RECT -175.665 89.510 -175.495 89.835 ;
        RECT -175.315 89.735 -174.945 90.075 ;
        RECT -174.765 89.835 -174.215 90.005 ;
        RECT -170.165 89.835 -169.615 90.005 ;
        RECT -174.765 89.510 -174.595 89.835 ;
        RECT -175.665 89.340 -174.595 89.510 ;
        RECT -169.785 89.510 -169.615 89.835 ;
        RECT -169.435 89.735 -169.065 90.075 ;
        RECT -168.885 89.835 -167.955 90.015 ;
        RECT -166.505 89.835 -165.575 90.015 ;
        RECT -168.885 89.510 -168.715 89.835 ;
        RECT -169.785 89.340 -168.715 89.510 ;
        RECT -165.745 89.510 -165.575 89.835 ;
        RECT -165.395 89.735 -165.025 90.075 ;
        RECT -164.845 89.835 -164.295 90.005 ;
        RECT -160.245 89.835 -159.695 90.005 ;
        RECT -164.845 89.510 -164.675 89.835 ;
        RECT -165.745 89.340 -164.675 89.510 ;
        RECT -159.865 89.510 -159.695 89.835 ;
        RECT -159.515 89.735 -159.145 90.075 ;
        RECT -158.965 89.835 -158.035 90.015 ;
        RECT -156.585 89.835 -155.655 90.015 ;
        RECT -158.965 89.510 -158.795 89.835 ;
        RECT -159.865 89.340 -158.795 89.510 ;
        RECT -155.825 89.510 -155.655 89.835 ;
        RECT -155.475 89.735 -155.105 90.075 ;
        RECT -154.925 89.835 -154.375 90.005 ;
        RECT -150.325 89.835 -149.775 90.005 ;
        RECT -154.925 89.510 -154.755 89.835 ;
        RECT -155.825 89.340 -154.755 89.510 ;
        RECT -149.945 89.510 -149.775 89.835 ;
        RECT -149.595 89.735 -149.225 90.075 ;
        RECT -149.045 89.835 -148.115 90.015 ;
        RECT -146.665 89.835 -145.735 90.015 ;
        RECT -149.045 89.510 -148.875 89.835 ;
        RECT -149.945 89.340 -148.875 89.510 ;
        RECT -145.905 89.510 -145.735 89.835 ;
        RECT -145.555 89.735 -145.185 90.075 ;
        RECT -145.005 89.835 -144.455 90.005 ;
        RECT -140.405 89.835 -139.855 90.005 ;
        RECT -145.005 89.510 -144.835 89.835 ;
        RECT -145.905 89.340 -144.835 89.510 ;
        RECT -140.025 89.510 -139.855 89.835 ;
        RECT -139.675 89.735 -139.305 90.075 ;
        RECT -139.125 89.835 -138.195 90.015 ;
        RECT -136.745 89.835 -135.815 90.015 ;
        RECT -139.125 89.510 -138.955 89.835 ;
        RECT -140.025 89.340 -138.955 89.510 ;
        RECT -135.985 89.510 -135.815 89.835 ;
        RECT -135.635 89.735 -135.265 90.075 ;
        RECT -135.085 89.835 -134.535 90.005 ;
        RECT -130.485 89.835 -129.935 90.005 ;
        RECT -135.085 89.510 -134.915 89.835 ;
        RECT -135.985 89.340 -134.915 89.510 ;
        RECT -130.105 89.510 -129.935 89.835 ;
        RECT -129.755 89.735 -129.385 90.075 ;
        RECT -129.205 89.835 -128.275 90.015 ;
        RECT -126.825 89.835 -125.895 90.015 ;
        RECT -129.205 89.510 -129.035 89.835 ;
        RECT -130.105 89.340 -129.035 89.510 ;
        RECT -126.065 89.510 -125.895 89.835 ;
        RECT -125.715 89.735 -125.345 90.075 ;
        RECT -125.165 89.835 -124.615 90.005 ;
        RECT -120.565 89.835 -120.015 90.005 ;
        RECT -125.165 89.510 -124.995 89.835 ;
        RECT -126.065 89.340 -124.995 89.510 ;
        RECT -120.185 89.510 -120.015 89.835 ;
        RECT -119.835 89.735 -119.465 90.075 ;
        RECT -119.285 89.835 -118.355 90.015 ;
        RECT -116.905 89.835 -115.975 90.015 ;
        RECT -119.285 89.510 -119.115 89.835 ;
        RECT -120.185 89.340 -119.115 89.510 ;
        RECT -116.145 89.510 -115.975 89.835 ;
        RECT -115.795 89.735 -115.425 90.075 ;
        RECT -115.245 89.835 -114.695 90.005 ;
        RECT -110.645 89.835 -110.095 90.005 ;
        RECT -115.245 89.510 -115.075 89.835 ;
        RECT -116.145 89.340 -115.075 89.510 ;
        RECT -110.265 89.510 -110.095 89.835 ;
        RECT -109.915 89.735 -109.545 90.075 ;
        RECT -109.365 89.835 -108.435 90.015 ;
        RECT -106.985 89.835 -106.055 90.015 ;
        RECT -109.365 89.510 -109.195 89.835 ;
        RECT -110.265 89.340 -109.195 89.510 ;
        RECT -106.225 89.510 -106.055 89.835 ;
        RECT -105.875 89.735 -105.505 90.075 ;
        RECT -105.325 89.835 -104.775 90.005 ;
        RECT -100.725 89.835 -100.175 90.005 ;
        RECT -105.325 89.510 -105.155 89.835 ;
        RECT -106.225 89.340 -105.155 89.510 ;
        RECT -100.345 89.510 -100.175 89.835 ;
        RECT -99.995 89.735 -99.625 90.075 ;
        RECT -99.445 89.835 -98.515 90.015 ;
        RECT -97.065 89.835 -96.135 90.015 ;
        RECT -99.445 89.510 -99.275 89.835 ;
        RECT -100.345 89.340 -99.275 89.510 ;
        RECT -96.305 89.510 -96.135 89.835 ;
        RECT -95.955 89.735 -95.585 90.075 ;
        RECT -95.405 89.835 -94.855 90.005 ;
        RECT -90.805 89.835 -90.255 90.005 ;
        RECT -95.405 89.510 -95.235 89.835 ;
        RECT -96.305 89.340 -95.235 89.510 ;
        RECT -90.425 89.510 -90.255 89.835 ;
        RECT -90.075 89.735 -89.705 90.075 ;
        RECT -89.525 89.835 -88.595 90.015 ;
        RECT -87.145 89.835 -86.215 90.015 ;
        RECT -89.525 89.510 -89.355 89.835 ;
        RECT -90.425 89.340 -89.355 89.510 ;
        RECT -86.385 89.510 -86.215 89.835 ;
        RECT -86.035 89.735 -85.665 90.075 ;
        RECT -85.485 89.835 -84.935 90.005 ;
        RECT -80.885 89.835 -80.335 90.005 ;
        RECT -85.485 89.510 -85.315 89.835 ;
        RECT -86.385 89.340 -85.315 89.510 ;
        RECT -80.505 89.510 -80.335 89.835 ;
        RECT -80.155 89.735 -79.785 90.075 ;
        RECT -79.605 89.835 -78.675 90.015 ;
        RECT -77.225 89.835 -76.295 90.015 ;
        RECT -79.605 89.510 -79.435 89.835 ;
        RECT -80.505 89.340 -79.435 89.510 ;
        RECT -76.465 89.510 -76.295 89.835 ;
        RECT -76.115 89.735 -75.745 90.075 ;
        RECT -75.565 89.835 -75.015 90.005 ;
        RECT -70.965 89.835 -70.415 90.005 ;
        RECT -75.565 89.510 -75.395 89.835 ;
        RECT -76.465 89.340 -75.395 89.510 ;
        RECT -70.585 89.510 -70.415 89.835 ;
        RECT -70.235 89.735 -69.865 90.075 ;
        RECT -69.685 89.835 -68.755 90.015 ;
        RECT -67.305 89.835 -66.375 90.015 ;
        RECT -69.685 89.510 -69.515 89.835 ;
        RECT -70.585 89.340 -69.515 89.510 ;
        RECT -66.545 89.510 -66.375 89.835 ;
        RECT -66.195 89.735 -65.825 90.075 ;
        RECT -65.645 89.835 -65.095 90.005 ;
        RECT -61.045 89.835 -60.495 90.005 ;
        RECT -65.645 89.510 -65.475 89.835 ;
        RECT -66.545 89.340 -65.475 89.510 ;
        RECT -60.665 89.510 -60.495 89.835 ;
        RECT -60.315 89.735 -59.945 90.075 ;
        RECT -59.765 89.835 -58.835 90.015 ;
        RECT -57.385 89.835 -56.455 90.015 ;
        RECT -59.765 89.510 -59.595 89.835 ;
        RECT -60.665 89.340 -59.595 89.510 ;
        RECT -56.625 89.510 -56.455 89.835 ;
        RECT -56.275 89.735 -55.905 90.075 ;
        RECT -55.725 89.835 -55.175 90.005 ;
        RECT -51.125 89.835 -50.575 90.005 ;
        RECT -55.725 89.510 -55.555 89.835 ;
        RECT -56.625 89.340 -55.555 89.510 ;
        RECT -50.745 89.510 -50.575 89.835 ;
        RECT -50.395 89.735 -50.025 90.075 ;
        RECT -49.845 89.835 -48.915 90.015 ;
        RECT -47.465 89.835 -46.535 90.015 ;
        RECT -49.845 89.510 -49.675 89.835 ;
        RECT -50.745 89.340 -49.675 89.510 ;
        RECT -46.705 89.510 -46.535 89.835 ;
        RECT -46.355 89.735 -45.985 90.075 ;
        RECT -45.805 89.835 -45.255 90.005 ;
        RECT -41.205 89.835 -40.655 90.005 ;
        RECT -45.805 89.510 -45.635 89.835 ;
        RECT -46.705 89.340 -45.635 89.510 ;
        RECT -40.825 89.510 -40.655 89.835 ;
        RECT -40.475 89.735 -40.105 90.075 ;
        RECT -39.925 89.835 -38.995 90.015 ;
        RECT -37.545 89.835 -36.615 90.015 ;
        RECT -39.925 89.510 -39.755 89.835 ;
        RECT -40.825 89.340 -39.755 89.510 ;
        RECT -36.785 89.510 -36.615 89.835 ;
        RECT -36.435 89.735 -36.065 90.075 ;
        RECT -35.885 89.835 -35.335 90.005 ;
        RECT -31.285 89.835 -30.735 90.005 ;
        RECT -35.885 89.510 -35.715 89.835 ;
        RECT -36.785 89.340 -35.715 89.510 ;
        RECT -30.905 89.510 -30.735 89.835 ;
        RECT -30.555 89.735 -30.185 90.075 ;
        RECT -30.005 89.835 -29.075 90.015 ;
        RECT -27.625 89.835 -26.695 90.015 ;
        RECT -30.005 89.510 -29.835 89.835 ;
        RECT -30.905 89.340 -29.835 89.510 ;
        RECT -26.865 89.510 -26.695 89.835 ;
        RECT -26.515 89.735 -26.145 90.075 ;
        RECT -25.965 89.835 -25.415 90.005 ;
        RECT -21.365 89.835 -20.815 90.005 ;
        RECT -25.965 89.510 -25.795 89.835 ;
        RECT -26.865 89.340 -25.795 89.510 ;
        RECT -20.985 89.510 -20.815 89.835 ;
        RECT -20.635 89.735 -20.265 90.075 ;
        RECT -20.085 89.835 -19.155 90.015 ;
        RECT -17.705 89.835 -16.775 90.015 ;
        RECT -20.085 89.510 -19.915 89.835 ;
        RECT -20.985 89.340 -19.915 89.510 ;
        RECT -16.945 89.510 -16.775 89.835 ;
        RECT -16.595 89.735 -16.225 90.075 ;
        RECT -16.045 89.835 -15.495 90.005 ;
        RECT -11.445 89.835 -10.895 90.005 ;
        RECT -16.045 89.510 -15.875 89.835 ;
        RECT -16.945 89.340 -15.875 89.510 ;
        RECT -11.065 89.510 -10.895 89.835 ;
        RECT -10.715 89.735 -10.345 90.075 ;
        RECT -10.165 89.835 -9.235 90.015 ;
        RECT -7.785 89.835 -6.855 90.015 ;
        RECT -10.165 89.510 -9.995 89.835 ;
        RECT -11.065 89.340 -9.995 89.510 ;
        RECT -7.025 89.510 -6.855 89.835 ;
        RECT -6.675 89.735 -6.305 90.075 ;
        RECT -6.125 89.835 -5.575 90.005 ;
        RECT -1.525 89.835 -0.975 90.005 ;
        RECT -6.125 89.510 -5.955 89.835 ;
        RECT -7.025 89.340 -5.955 89.510 ;
        RECT -1.145 89.510 -0.975 89.835 ;
        RECT -0.795 89.735 -0.425 90.075 ;
        RECT -0.245 89.835 0.685 90.015 ;
        RECT 2.135 89.835 3.065 90.015 ;
        RECT -0.245 89.510 -0.075 89.835 ;
        RECT -1.145 89.340 -0.075 89.510 ;
        RECT 2.895 89.510 3.065 89.835 ;
        RECT 3.245 89.735 3.615 90.075 ;
        RECT 3.795 89.835 4.345 90.005 ;
        RECT 8.395 89.835 8.945 90.005 ;
        RECT 3.795 89.510 3.965 89.835 ;
        RECT 2.895 89.340 3.965 89.510 ;
        RECT 8.775 89.510 8.945 89.835 ;
        RECT 9.125 89.735 9.495 90.075 ;
        RECT 9.675 89.835 10.605 90.015 ;
        RECT 12.055 89.835 12.985 90.015 ;
        RECT 9.675 89.510 9.845 89.835 ;
        RECT 8.775 89.340 9.845 89.510 ;
        RECT 12.815 89.510 12.985 89.835 ;
        RECT 13.165 89.735 13.535 90.075 ;
        RECT 13.715 89.835 14.265 90.005 ;
        RECT 18.315 89.835 18.865 90.005 ;
        RECT 13.715 89.510 13.885 89.835 ;
        RECT 12.815 89.340 13.885 89.510 ;
        RECT 18.695 89.510 18.865 89.835 ;
        RECT 19.045 89.735 19.415 90.075 ;
        RECT 19.595 89.835 20.525 90.015 ;
        RECT 21.975 89.835 22.905 90.015 ;
        RECT 19.595 89.510 19.765 89.835 ;
        RECT 18.695 89.340 19.765 89.510 ;
        RECT 22.735 89.510 22.905 89.835 ;
        RECT 23.085 89.735 23.455 90.075 ;
        RECT 23.635 89.835 24.185 90.005 ;
        RECT 23.635 89.510 23.805 89.835 ;
        RECT 24.355 89.655 24.525 90.180 ;
        RECT 22.735 89.340 23.805 89.510 ;
        RECT -289.545 89.140 -289.375 89.325 ;
        RECT -288.400 89.235 -288.070 89.340 ;
        RECT -284.470 89.235 -284.140 89.340 ;
        RECT -278.480 89.235 -278.150 89.340 ;
        RECT -274.550 89.235 -274.220 89.340 ;
        RECT -268.560 89.235 -268.230 89.340 ;
        RECT -264.630 89.235 -264.300 89.340 ;
        RECT -258.640 89.235 -258.310 89.340 ;
        RECT -254.710 89.235 -254.380 89.340 ;
        RECT -248.720 89.235 -248.390 89.340 ;
        RECT -244.790 89.235 -244.460 89.340 ;
        RECT -238.800 89.235 -238.470 89.340 ;
        RECT -234.870 89.235 -234.540 89.340 ;
        RECT -228.880 89.235 -228.550 89.340 ;
        RECT -224.950 89.235 -224.620 89.340 ;
        RECT -218.960 89.235 -218.630 89.340 ;
        RECT -215.030 89.235 -214.700 89.340 ;
        RECT -209.040 89.235 -208.710 89.340 ;
        RECT -205.110 89.235 -204.780 89.340 ;
        RECT -199.120 89.235 -198.790 89.340 ;
        RECT -195.190 89.235 -194.860 89.340 ;
        RECT -189.200 89.235 -188.870 89.340 ;
        RECT -185.270 89.235 -184.940 89.340 ;
        RECT -179.280 89.235 -178.950 89.340 ;
        RECT -175.350 89.235 -175.020 89.340 ;
        RECT -169.360 89.235 -169.030 89.340 ;
        RECT -165.430 89.235 -165.100 89.340 ;
        RECT -159.440 89.235 -159.110 89.340 ;
        RECT -155.510 89.235 -155.180 89.340 ;
        RECT -149.520 89.235 -149.190 89.340 ;
        RECT -145.590 89.235 -145.260 89.340 ;
        RECT -139.600 89.235 -139.270 89.340 ;
        RECT -135.670 89.235 -135.340 89.340 ;
        RECT -129.680 89.235 -129.350 89.340 ;
        RECT -125.750 89.235 -125.420 89.340 ;
        RECT -119.760 89.235 -119.430 89.340 ;
        RECT -115.830 89.235 -115.500 89.340 ;
        RECT -109.840 89.235 -109.510 89.340 ;
        RECT -105.910 89.235 -105.580 89.340 ;
        RECT -99.920 89.235 -99.590 89.340 ;
        RECT -95.990 89.235 -95.660 89.340 ;
        RECT -90.000 89.235 -89.670 89.340 ;
        RECT -86.070 89.235 -85.740 89.340 ;
        RECT -80.080 89.235 -79.750 89.340 ;
        RECT -76.150 89.235 -75.820 89.340 ;
        RECT -70.160 89.235 -69.830 89.340 ;
        RECT -66.230 89.235 -65.900 89.340 ;
        RECT -60.240 89.235 -59.910 89.340 ;
        RECT -56.310 89.235 -55.980 89.340 ;
        RECT -50.320 89.235 -49.990 89.340 ;
        RECT -46.390 89.235 -46.060 89.340 ;
        RECT -40.400 89.235 -40.070 89.340 ;
        RECT -36.470 89.235 -36.140 89.340 ;
        RECT -30.480 89.235 -30.150 89.340 ;
        RECT -26.550 89.235 -26.220 89.340 ;
        RECT -20.560 89.235 -20.230 89.340 ;
        RECT -16.630 89.235 -16.300 89.340 ;
        RECT -10.640 89.235 -10.310 89.340 ;
        RECT -6.710 89.235 -6.380 89.340 ;
        RECT -0.720 89.235 -0.390 89.340 ;
        RECT 3.210 89.235 3.540 89.340 ;
        RECT 9.200 89.235 9.530 89.340 ;
        RECT 13.130 89.235 13.460 89.340 ;
        RECT 19.120 89.235 19.450 89.340 ;
        RECT 23.050 89.235 23.380 89.340 ;
        RECT 23.975 89.325 24.525 89.655 ;
        RECT -290.075 89.125 -289.375 89.140 ;
        RECT -290.160 88.955 -289.375 89.125 ;
        RECT -289.840 88.950 -289.375 88.955 ;
        RECT -289.545 88.800 -289.375 88.950 ;
        RECT -285.545 89.065 -284.640 89.155 ;
        RECT -283.840 89.065 -283.335 89.145 ;
        RECT -285.545 88.885 -283.335 89.065 ;
        RECT -275.625 89.065 -274.720 89.155 ;
        RECT -273.920 89.065 -273.415 89.145 ;
        RECT -275.625 88.885 -273.415 89.065 ;
        RECT -265.705 89.065 -264.800 89.155 ;
        RECT -264.000 89.065 -263.495 89.145 ;
        RECT -265.705 88.885 -263.495 89.065 ;
        RECT -255.785 89.065 -254.880 89.155 ;
        RECT -254.080 89.065 -253.575 89.145 ;
        RECT -255.785 88.885 -253.575 89.065 ;
        RECT -245.865 89.065 -244.960 89.155 ;
        RECT -244.160 89.065 -243.655 89.145 ;
        RECT -245.865 88.885 -243.655 89.065 ;
        RECT -235.945 89.065 -235.040 89.155 ;
        RECT -234.240 89.065 -233.735 89.145 ;
        RECT -235.945 88.885 -233.735 89.065 ;
        RECT -226.025 89.065 -225.120 89.155 ;
        RECT -224.320 89.065 -223.815 89.145 ;
        RECT -226.025 88.885 -223.815 89.065 ;
        RECT -216.105 89.065 -215.200 89.155 ;
        RECT -214.400 89.065 -213.895 89.145 ;
        RECT -216.105 88.885 -213.895 89.065 ;
        RECT -206.185 89.065 -205.280 89.155 ;
        RECT -204.480 89.065 -203.975 89.145 ;
        RECT -206.185 88.885 -203.975 89.065 ;
        RECT -196.265 89.065 -195.360 89.155 ;
        RECT -194.560 89.065 -194.055 89.145 ;
        RECT -196.265 88.885 -194.055 89.065 ;
        RECT -186.345 89.065 -185.440 89.155 ;
        RECT -184.640 89.065 -184.135 89.145 ;
        RECT -186.345 88.885 -184.135 89.065 ;
        RECT -176.425 89.065 -175.520 89.155 ;
        RECT -174.720 89.065 -174.215 89.145 ;
        RECT -176.425 88.885 -174.215 89.065 ;
        RECT -166.505 89.065 -165.600 89.155 ;
        RECT -164.800 89.065 -164.295 89.145 ;
        RECT -166.505 88.885 -164.295 89.065 ;
        RECT -156.585 89.065 -155.680 89.155 ;
        RECT -154.880 89.065 -154.375 89.145 ;
        RECT -156.585 88.885 -154.375 89.065 ;
        RECT -146.665 89.065 -145.760 89.155 ;
        RECT -144.960 89.065 -144.455 89.145 ;
        RECT -146.665 88.885 -144.455 89.065 ;
        RECT -136.745 89.065 -135.840 89.155 ;
        RECT -135.040 89.065 -134.535 89.145 ;
        RECT -136.745 88.885 -134.535 89.065 ;
        RECT -126.825 89.065 -125.920 89.155 ;
        RECT -125.120 89.065 -124.615 89.145 ;
        RECT -126.825 88.885 -124.615 89.065 ;
        RECT -116.905 89.065 -116.000 89.155 ;
        RECT -115.200 89.065 -114.695 89.145 ;
        RECT -116.905 88.885 -114.695 89.065 ;
        RECT -106.985 89.065 -106.080 89.155 ;
        RECT -105.280 89.065 -104.775 89.145 ;
        RECT -106.985 88.885 -104.775 89.065 ;
        RECT -97.065 89.065 -96.160 89.155 ;
        RECT -95.360 89.065 -94.855 89.145 ;
        RECT -97.065 88.885 -94.855 89.065 ;
        RECT -87.145 89.065 -86.240 89.155 ;
        RECT -85.440 89.065 -84.935 89.145 ;
        RECT -87.145 88.885 -84.935 89.065 ;
        RECT -77.225 89.065 -76.320 89.155 ;
        RECT -75.520 89.065 -75.015 89.145 ;
        RECT -77.225 88.885 -75.015 89.065 ;
        RECT -67.305 89.065 -66.400 89.155 ;
        RECT -65.600 89.065 -65.095 89.145 ;
        RECT -67.305 88.885 -65.095 89.065 ;
        RECT -57.385 89.065 -56.480 89.155 ;
        RECT -55.680 89.065 -55.175 89.145 ;
        RECT -57.385 88.885 -55.175 89.065 ;
        RECT -47.465 89.065 -46.560 89.155 ;
        RECT -45.760 89.065 -45.255 89.145 ;
        RECT -47.465 88.885 -45.255 89.065 ;
        RECT -37.545 89.065 -36.640 89.155 ;
        RECT -35.840 89.065 -35.335 89.145 ;
        RECT -37.545 88.885 -35.335 89.065 ;
        RECT -27.625 89.065 -26.720 89.155 ;
        RECT -25.920 89.065 -25.415 89.145 ;
        RECT -27.625 88.885 -25.415 89.065 ;
        RECT -17.705 89.065 -16.800 89.155 ;
        RECT -16.000 89.065 -15.495 89.145 ;
        RECT -17.705 88.885 -15.495 89.065 ;
        RECT -7.785 89.065 -6.880 89.155 ;
        RECT -6.080 89.065 -5.575 89.145 ;
        RECT -7.785 88.885 -5.575 89.065 ;
        RECT 2.135 89.065 3.040 89.155 ;
        RECT 3.840 89.065 4.345 89.145 ;
        RECT 2.135 88.885 4.345 89.065 ;
        RECT 12.055 89.065 12.960 89.155 ;
        RECT 13.760 89.065 14.265 89.145 ;
        RECT 12.055 88.885 14.265 89.065 ;
        RECT 21.975 89.065 22.880 89.155 ;
        RECT 23.680 89.065 24.185 89.145 ;
        RECT 21.975 88.885 24.185 89.065 ;
        RECT 24.355 89.130 24.525 89.325 ;
        RECT 24.765 89.130 25.055 89.850 ;
        RECT 24.355 89.125 25.055 89.130 ;
        RECT 24.355 88.955 25.140 89.125 ;
        RECT 24.355 88.950 24.820 88.955 ;
        RECT 24.355 88.800 24.525 88.950 ;
        RECT -290.595 7.280 -290.425 7.430 ;
        RECT -291.210 7.110 -290.425 7.280 ;
        RECT -291.125 5.945 -290.835 7.110 ;
        RECT -290.595 6.905 -290.425 7.110 ;
        RECT -290.255 7.165 -288.045 7.345 ;
        RECT -290.255 7.075 -289.350 7.165 ;
        RECT -288.550 7.085 -288.045 7.165 ;
        RECT -280.335 7.165 -278.125 7.345 ;
        RECT -280.335 7.075 -279.430 7.165 ;
        RECT -278.630 7.085 -278.125 7.165 ;
        RECT -270.415 7.165 -268.205 7.345 ;
        RECT -270.415 7.075 -269.510 7.165 ;
        RECT -268.710 7.085 -268.205 7.165 ;
        RECT -260.495 7.165 -258.285 7.345 ;
        RECT -260.495 7.075 -259.590 7.165 ;
        RECT -258.790 7.085 -258.285 7.165 ;
        RECT -250.575 7.165 -248.365 7.345 ;
        RECT -250.575 7.075 -249.670 7.165 ;
        RECT -248.870 7.085 -248.365 7.165 ;
        RECT -240.655 7.165 -238.445 7.345 ;
        RECT -240.655 7.075 -239.750 7.165 ;
        RECT -238.950 7.085 -238.445 7.165 ;
        RECT -230.735 7.165 -228.525 7.345 ;
        RECT -230.735 7.075 -229.830 7.165 ;
        RECT -229.030 7.085 -228.525 7.165 ;
        RECT -220.815 7.165 -218.605 7.345 ;
        RECT -220.815 7.075 -219.910 7.165 ;
        RECT -219.110 7.085 -218.605 7.165 ;
        RECT -210.895 7.165 -208.685 7.345 ;
        RECT -210.895 7.075 -209.990 7.165 ;
        RECT -209.190 7.085 -208.685 7.165 ;
        RECT -200.975 7.165 -198.765 7.345 ;
        RECT -200.975 7.075 -200.070 7.165 ;
        RECT -199.270 7.085 -198.765 7.165 ;
        RECT -191.055 7.165 -188.845 7.345 ;
        RECT -191.055 7.075 -190.150 7.165 ;
        RECT -189.350 7.085 -188.845 7.165 ;
        RECT -181.135 7.165 -178.925 7.345 ;
        RECT -181.135 7.075 -180.230 7.165 ;
        RECT -179.430 7.085 -178.925 7.165 ;
        RECT -171.215 7.165 -169.005 7.345 ;
        RECT -171.215 7.075 -170.310 7.165 ;
        RECT -169.510 7.085 -169.005 7.165 ;
        RECT -161.295 7.165 -159.085 7.345 ;
        RECT -161.295 7.075 -160.390 7.165 ;
        RECT -159.590 7.085 -159.085 7.165 ;
        RECT -151.375 7.165 -149.165 7.345 ;
        RECT -151.375 7.075 -150.470 7.165 ;
        RECT -149.670 7.085 -149.165 7.165 ;
        RECT -141.455 7.165 -139.245 7.345 ;
        RECT -141.455 7.075 -140.550 7.165 ;
        RECT -139.750 7.085 -139.245 7.165 ;
        RECT -131.535 7.165 -129.325 7.345 ;
        RECT -131.535 7.075 -130.630 7.165 ;
        RECT -129.830 7.085 -129.325 7.165 ;
        RECT -121.615 7.165 -119.405 7.345 ;
        RECT -121.615 7.075 -120.710 7.165 ;
        RECT -119.910 7.085 -119.405 7.165 ;
        RECT -111.695 7.165 -109.485 7.345 ;
        RECT -111.695 7.075 -110.790 7.165 ;
        RECT -109.990 7.085 -109.485 7.165 ;
        RECT -101.775 7.165 -99.565 7.345 ;
        RECT -101.775 7.075 -100.870 7.165 ;
        RECT -100.070 7.085 -99.565 7.165 ;
        RECT -91.855 7.165 -89.645 7.345 ;
        RECT -91.855 7.075 -90.950 7.165 ;
        RECT -90.150 7.085 -89.645 7.165 ;
        RECT -81.935 7.165 -79.725 7.345 ;
        RECT -81.935 7.075 -81.030 7.165 ;
        RECT -80.230 7.085 -79.725 7.165 ;
        RECT -72.015 7.165 -69.805 7.345 ;
        RECT -72.015 7.075 -71.110 7.165 ;
        RECT -70.310 7.085 -69.805 7.165 ;
        RECT -62.095 7.165 -59.885 7.345 ;
        RECT -62.095 7.075 -61.190 7.165 ;
        RECT -60.390 7.085 -59.885 7.165 ;
        RECT -52.175 7.165 -49.965 7.345 ;
        RECT -52.175 7.075 -51.270 7.165 ;
        RECT -50.470 7.085 -49.965 7.165 ;
        RECT -42.255 7.165 -40.045 7.345 ;
        RECT -42.255 7.075 -41.350 7.165 ;
        RECT -40.550 7.085 -40.045 7.165 ;
        RECT -32.335 7.165 -30.125 7.345 ;
        RECT -32.335 7.075 -31.430 7.165 ;
        RECT -30.630 7.085 -30.125 7.165 ;
        RECT -22.415 7.165 -20.205 7.345 ;
        RECT -22.415 7.075 -21.510 7.165 ;
        RECT -20.710 7.085 -20.205 7.165 ;
        RECT -12.495 7.165 -10.285 7.345 ;
        RECT -12.495 7.075 -11.590 7.165 ;
        RECT -10.790 7.085 -10.285 7.165 ;
        RECT -2.575 7.165 -0.365 7.345 ;
        RECT -2.575 7.075 -1.670 7.165 ;
        RECT -0.870 7.085 -0.365 7.165 ;
        RECT 7.345 7.165 9.555 7.345 ;
        RECT 7.345 7.075 8.250 7.165 ;
        RECT 9.050 7.085 9.555 7.165 ;
        RECT 17.265 7.165 19.475 7.345 ;
        RECT 17.265 7.075 18.170 7.165 ;
        RECT 18.970 7.085 19.475 7.165 ;
        RECT -290.595 6.575 -289.665 6.905 ;
        RECT -289.180 6.890 -288.850 6.995 ;
        RECT -283.190 6.890 -282.860 6.995 ;
        RECT -279.260 6.890 -278.930 6.995 ;
        RECT -273.270 6.890 -272.940 6.995 ;
        RECT -269.340 6.890 -269.010 6.995 ;
        RECT -263.350 6.890 -263.020 6.995 ;
        RECT -259.420 6.890 -259.090 6.995 ;
        RECT -253.430 6.890 -253.100 6.995 ;
        RECT -249.500 6.890 -249.170 6.995 ;
        RECT -243.510 6.890 -243.180 6.995 ;
        RECT -239.580 6.890 -239.250 6.995 ;
        RECT -233.590 6.890 -233.260 6.995 ;
        RECT -229.660 6.890 -229.330 6.995 ;
        RECT -223.670 6.890 -223.340 6.995 ;
        RECT -219.740 6.890 -219.410 6.995 ;
        RECT -213.750 6.890 -213.420 6.995 ;
        RECT -209.820 6.890 -209.490 6.995 ;
        RECT -203.830 6.890 -203.500 6.995 ;
        RECT -199.900 6.890 -199.570 6.995 ;
        RECT -193.910 6.890 -193.580 6.995 ;
        RECT -189.980 6.890 -189.650 6.995 ;
        RECT -183.990 6.890 -183.660 6.995 ;
        RECT -180.060 6.890 -179.730 6.995 ;
        RECT -174.070 6.890 -173.740 6.995 ;
        RECT -170.140 6.890 -169.810 6.995 ;
        RECT -164.150 6.890 -163.820 6.995 ;
        RECT -160.220 6.890 -159.890 6.995 ;
        RECT -154.230 6.890 -153.900 6.995 ;
        RECT -150.300 6.890 -149.970 6.995 ;
        RECT -144.310 6.890 -143.980 6.995 ;
        RECT -140.380 6.890 -140.050 6.995 ;
        RECT -134.390 6.890 -134.060 6.995 ;
        RECT -130.460 6.890 -130.130 6.995 ;
        RECT -124.470 6.890 -124.140 6.995 ;
        RECT -120.540 6.890 -120.210 6.995 ;
        RECT -114.550 6.890 -114.220 6.995 ;
        RECT -110.620 6.890 -110.290 6.995 ;
        RECT -104.630 6.890 -104.300 6.995 ;
        RECT -100.700 6.890 -100.370 6.995 ;
        RECT -94.710 6.890 -94.380 6.995 ;
        RECT -90.780 6.890 -90.450 6.995 ;
        RECT -84.790 6.890 -84.460 6.995 ;
        RECT -80.860 6.890 -80.530 6.995 ;
        RECT -74.870 6.890 -74.540 6.995 ;
        RECT -70.940 6.890 -70.610 6.995 ;
        RECT -64.950 6.890 -64.620 6.995 ;
        RECT -61.020 6.890 -60.690 6.995 ;
        RECT -55.030 6.890 -54.700 6.995 ;
        RECT -51.100 6.890 -50.770 6.995 ;
        RECT -45.110 6.890 -44.780 6.995 ;
        RECT -41.180 6.890 -40.850 6.995 ;
        RECT -35.190 6.890 -34.860 6.995 ;
        RECT -31.260 6.890 -30.930 6.995 ;
        RECT -25.270 6.890 -24.940 6.995 ;
        RECT -21.340 6.890 -21.010 6.995 ;
        RECT -15.350 6.890 -15.020 6.995 ;
        RECT -11.420 6.890 -11.090 6.995 ;
        RECT -5.430 6.890 -5.100 6.995 ;
        RECT -1.500 6.890 -1.170 6.995 ;
        RECT 4.490 6.890 4.820 6.995 ;
        RECT 8.420 6.890 8.750 6.995 ;
        RECT 14.410 6.890 14.740 6.995 ;
        RECT 18.340 6.890 18.670 6.995 ;
        RECT 24.330 6.890 24.660 6.995 ;
        RECT -289.495 6.720 -288.425 6.890 ;
        RECT -290.595 6.050 -290.425 6.575 ;
        RECT -289.495 6.395 -289.325 6.720 ;
        RECT -290.255 6.215 -289.325 6.395 ;
        RECT -289.145 6.155 -288.775 6.495 ;
        RECT -288.595 6.395 -288.425 6.720 ;
        RECT -283.615 6.720 -282.545 6.890 ;
        RECT -283.615 6.395 -283.445 6.720 ;
        RECT -288.595 6.225 -288.045 6.395 ;
        RECT -283.995 6.225 -283.445 6.395 ;
        RECT -283.265 6.155 -282.895 6.495 ;
        RECT -282.715 6.395 -282.545 6.720 ;
        RECT -279.575 6.720 -278.505 6.890 ;
        RECT -279.575 6.395 -279.405 6.720 ;
        RECT -282.715 6.215 -281.785 6.395 ;
        RECT -280.335 6.215 -279.405 6.395 ;
        RECT -279.225 6.155 -278.855 6.495 ;
        RECT -278.675 6.395 -278.505 6.720 ;
        RECT -273.695 6.720 -272.625 6.890 ;
        RECT -273.695 6.395 -273.525 6.720 ;
        RECT -278.675 6.225 -278.125 6.395 ;
        RECT -274.075 6.225 -273.525 6.395 ;
        RECT -273.345 6.155 -272.975 6.495 ;
        RECT -272.795 6.395 -272.625 6.720 ;
        RECT -269.655 6.720 -268.585 6.890 ;
        RECT -269.655 6.395 -269.485 6.720 ;
        RECT -272.795 6.215 -271.865 6.395 ;
        RECT -270.415 6.215 -269.485 6.395 ;
        RECT -269.305 6.155 -268.935 6.495 ;
        RECT -268.755 6.395 -268.585 6.720 ;
        RECT -263.775 6.720 -262.705 6.890 ;
        RECT -263.775 6.395 -263.605 6.720 ;
        RECT -268.755 6.225 -268.205 6.395 ;
        RECT -264.155 6.225 -263.605 6.395 ;
        RECT -263.425 6.155 -263.055 6.495 ;
        RECT -262.875 6.395 -262.705 6.720 ;
        RECT -259.735 6.720 -258.665 6.890 ;
        RECT -259.735 6.395 -259.565 6.720 ;
        RECT -262.875 6.215 -261.945 6.395 ;
        RECT -260.495 6.215 -259.565 6.395 ;
        RECT -259.385 6.155 -259.015 6.495 ;
        RECT -258.835 6.395 -258.665 6.720 ;
        RECT -253.855 6.720 -252.785 6.890 ;
        RECT -253.855 6.395 -253.685 6.720 ;
        RECT -258.835 6.225 -258.285 6.395 ;
        RECT -254.235 6.225 -253.685 6.395 ;
        RECT -253.505 6.155 -253.135 6.495 ;
        RECT -252.955 6.395 -252.785 6.720 ;
        RECT -249.815 6.720 -248.745 6.890 ;
        RECT -249.815 6.395 -249.645 6.720 ;
        RECT -252.955 6.215 -252.025 6.395 ;
        RECT -250.575 6.215 -249.645 6.395 ;
        RECT -249.465 6.155 -249.095 6.495 ;
        RECT -248.915 6.395 -248.745 6.720 ;
        RECT -243.935 6.720 -242.865 6.890 ;
        RECT -243.935 6.395 -243.765 6.720 ;
        RECT -248.915 6.225 -248.365 6.395 ;
        RECT -244.315 6.225 -243.765 6.395 ;
        RECT -243.585 6.155 -243.215 6.495 ;
        RECT -243.035 6.395 -242.865 6.720 ;
        RECT -239.895 6.720 -238.825 6.890 ;
        RECT -239.895 6.395 -239.725 6.720 ;
        RECT -243.035 6.215 -242.105 6.395 ;
        RECT -240.655 6.215 -239.725 6.395 ;
        RECT -239.545 6.155 -239.175 6.495 ;
        RECT -238.995 6.395 -238.825 6.720 ;
        RECT -234.015 6.720 -232.945 6.890 ;
        RECT -234.015 6.395 -233.845 6.720 ;
        RECT -238.995 6.225 -238.445 6.395 ;
        RECT -234.395 6.225 -233.845 6.395 ;
        RECT -233.665 6.155 -233.295 6.495 ;
        RECT -233.115 6.395 -232.945 6.720 ;
        RECT -229.975 6.720 -228.905 6.890 ;
        RECT -229.975 6.395 -229.805 6.720 ;
        RECT -233.115 6.215 -232.185 6.395 ;
        RECT -230.735 6.215 -229.805 6.395 ;
        RECT -229.625 6.155 -229.255 6.495 ;
        RECT -229.075 6.395 -228.905 6.720 ;
        RECT -224.095 6.720 -223.025 6.890 ;
        RECT -224.095 6.395 -223.925 6.720 ;
        RECT -229.075 6.225 -228.525 6.395 ;
        RECT -224.475 6.225 -223.925 6.395 ;
        RECT -223.745 6.155 -223.375 6.495 ;
        RECT -223.195 6.395 -223.025 6.720 ;
        RECT -220.055 6.720 -218.985 6.890 ;
        RECT -220.055 6.395 -219.885 6.720 ;
        RECT -223.195 6.215 -222.265 6.395 ;
        RECT -220.815 6.215 -219.885 6.395 ;
        RECT -219.705 6.155 -219.335 6.495 ;
        RECT -219.155 6.395 -218.985 6.720 ;
        RECT -214.175 6.720 -213.105 6.890 ;
        RECT -214.175 6.395 -214.005 6.720 ;
        RECT -219.155 6.225 -218.605 6.395 ;
        RECT -214.555 6.225 -214.005 6.395 ;
        RECT -213.825 6.155 -213.455 6.495 ;
        RECT -213.275 6.395 -213.105 6.720 ;
        RECT -210.135 6.720 -209.065 6.890 ;
        RECT -210.135 6.395 -209.965 6.720 ;
        RECT -213.275 6.215 -212.345 6.395 ;
        RECT -210.895 6.215 -209.965 6.395 ;
        RECT -209.785 6.155 -209.415 6.495 ;
        RECT -209.235 6.395 -209.065 6.720 ;
        RECT -204.255 6.720 -203.185 6.890 ;
        RECT -204.255 6.395 -204.085 6.720 ;
        RECT -209.235 6.225 -208.685 6.395 ;
        RECT -204.635 6.225 -204.085 6.395 ;
        RECT -203.905 6.155 -203.535 6.495 ;
        RECT -203.355 6.395 -203.185 6.720 ;
        RECT -200.215 6.720 -199.145 6.890 ;
        RECT -200.215 6.395 -200.045 6.720 ;
        RECT -203.355 6.215 -202.425 6.395 ;
        RECT -200.975 6.215 -200.045 6.395 ;
        RECT -199.865 6.155 -199.495 6.495 ;
        RECT -199.315 6.395 -199.145 6.720 ;
        RECT -194.335 6.720 -193.265 6.890 ;
        RECT -194.335 6.395 -194.165 6.720 ;
        RECT -199.315 6.225 -198.765 6.395 ;
        RECT -194.715 6.225 -194.165 6.395 ;
        RECT -193.985 6.155 -193.615 6.495 ;
        RECT -193.435 6.395 -193.265 6.720 ;
        RECT -190.295 6.720 -189.225 6.890 ;
        RECT -190.295 6.395 -190.125 6.720 ;
        RECT -193.435 6.215 -192.505 6.395 ;
        RECT -191.055 6.215 -190.125 6.395 ;
        RECT -189.945 6.155 -189.575 6.495 ;
        RECT -189.395 6.395 -189.225 6.720 ;
        RECT -184.415 6.720 -183.345 6.890 ;
        RECT -184.415 6.395 -184.245 6.720 ;
        RECT -189.395 6.225 -188.845 6.395 ;
        RECT -184.795 6.225 -184.245 6.395 ;
        RECT -184.065 6.155 -183.695 6.495 ;
        RECT -183.515 6.395 -183.345 6.720 ;
        RECT -180.375 6.720 -179.305 6.890 ;
        RECT -180.375 6.395 -180.205 6.720 ;
        RECT -183.515 6.215 -182.585 6.395 ;
        RECT -181.135 6.215 -180.205 6.395 ;
        RECT -180.025 6.155 -179.655 6.495 ;
        RECT -179.475 6.395 -179.305 6.720 ;
        RECT -174.495 6.720 -173.425 6.890 ;
        RECT -174.495 6.395 -174.325 6.720 ;
        RECT -179.475 6.225 -178.925 6.395 ;
        RECT -174.875 6.225 -174.325 6.395 ;
        RECT -174.145 6.155 -173.775 6.495 ;
        RECT -173.595 6.395 -173.425 6.720 ;
        RECT -170.455 6.720 -169.385 6.890 ;
        RECT -170.455 6.395 -170.285 6.720 ;
        RECT -173.595 6.215 -172.665 6.395 ;
        RECT -171.215 6.215 -170.285 6.395 ;
        RECT -170.105 6.155 -169.735 6.495 ;
        RECT -169.555 6.395 -169.385 6.720 ;
        RECT -164.575 6.720 -163.505 6.890 ;
        RECT -164.575 6.395 -164.405 6.720 ;
        RECT -169.555 6.225 -169.005 6.395 ;
        RECT -164.955 6.225 -164.405 6.395 ;
        RECT -164.225 6.155 -163.855 6.495 ;
        RECT -163.675 6.395 -163.505 6.720 ;
        RECT -160.535 6.720 -159.465 6.890 ;
        RECT -160.535 6.395 -160.365 6.720 ;
        RECT -163.675 6.215 -162.745 6.395 ;
        RECT -161.295 6.215 -160.365 6.395 ;
        RECT -160.185 6.155 -159.815 6.495 ;
        RECT -159.635 6.395 -159.465 6.720 ;
        RECT -154.655 6.720 -153.585 6.890 ;
        RECT -154.655 6.395 -154.485 6.720 ;
        RECT -159.635 6.225 -159.085 6.395 ;
        RECT -155.035 6.225 -154.485 6.395 ;
        RECT -154.305 6.155 -153.935 6.495 ;
        RECT -153.755 6.395 -153.585 6.720 ;
        RECT -150.615 6.720 -149.545 6.890 ;
        RECT -150.615 6.395 -150.445 6.720 ;
        RECT -153.755 6.215 -152.825 6.395 ;
        RECT -151.375 6.215 -150.445 6.395 ;
        RECT -150.265 6.155 -149.895 6.495 ;
        RECT -149.715 6.395 -149.545 6.720 ;
        RECT -144.735 6.720 -143.665 6.890 ;
        RECT -144.735 6.395 -144.565 6.720 ;
        RECT -149.715 6.225 -149.165 6.395 ;
        RECT -145.115 6.225 -144.565 6.395 ;
        RECT -144.385 6.155 -144.015 6.495 ;
        RECT -143.835 6.395 -143.665 6.720 ;
        RECT -140.695 6.720 -139.625 6.890 ;
        RECT -140.695 6.395 -140.525 6.720 ;
        RECT -143.835 6.215 -142.905 6.395 ;
        RECT -141.455 6.215 -140.525 6.395 ;
        RECT -140.345 6.155 -139.975 6.495 ;
        RECT -139.795 6.395 -139.625 6.720 ;
        RECT -134.815 6.720 -133.745 6.890 ;
        RECT -134.815 6.395 -134.645 6.720 ;
        RECT -139.795 6.225 -139.245 6.395 ;
        RECT -135.195 6.225 -134.645 6.395 ;
        RECT -134.465 6.155 -134.095 6.495 ;
        RECT -133.915 6.395 -133.745 6.720 ;
        RECT -130.775 6.720 -129.705 6.890 ;
        RECT -130.775 6.395 -130.605 6.720 ;
        RECT -133.915 6.215 -132.985 6.395 ;
        RECT -131.535 6.215 -130.605 6.395 ;
        RECT -130.425 6.155 -130.055 6.495 ;
        RECT -129.875 6.395 -129.705 6.720 ;
        RECT -124.895 6.720 -123.825 6.890 ;
        RECT -124.895 6.395 -124.725 6.720 ;
        RECT -129.875 6.225 -129.325 6.395 ;
        RECT -125.275 6.225 -124.725 6.395 ;
        RECT -124.545 6.155 -124.175 6.495 ;
        RECT -123.995 6.395 -123.825 6.720 ;
        RECT -120.855 6.720 -119.785 6.890 ;
        RECT -120.855 6.395 -120.685 6.720 ;
        RECT -123.995 6.215 -123.065 6.395 ;
        RECT -121.615 6.215 -120.685 6.395 ;
        RECT -120.505 6.155 -120.135 6.495 ;
        RECT -119.955 6.395 -119.785 6.720 ;
        RECT -114.975 6.720 -113.905 6.890 ;
        RECT -114.975 6.395 -114.805 6.720 ;
        RECT -119.955 6.225 -119.405 6.395 ;
        RECT -115.355 6.225 -114.805 6.395 ;
        RECT -114.625 6.155 -114.255 6.495 ;
        RECT -114.075 6.395 -113.905 6.720 ;
        RECT -110.935 6.720 -109.865 6.890 ;
        RECT -110.935 6.395 -110.765 6.720 ;
        RECT -114.075 6.215 -113.145 6.395 ;
        RECT -111.695 6.215 -110.765 6.395 ;
        RECT -110.585 6.155 -110.215 6.495 ;
        RECT -110.035 6.395 -109.865 6.720 ;
        RECT -105.055 6.720 -103.985 6.890 ;
        RECT -105.055 6.395 -104.885 6.720 ;
        RECT -110.035 6.225 -109.485 6.395 ;
        RECT -105.435 6.225 -104.885 6.395 ;
        RECT -104.705 6.155 -104.335 6.495 ;
        RECT -104.155 6.395 -103.985 6.720 ;
        RECT -101.015 6.720 -99.945 6.890 ;
        RECT -101.015 6.395 -100.845 6.720 ;
        RECT -104.155 6.215 -103.225 6.395 ;
        RECT -101.775 6.215 -100.845 6.395 ;
        RECT -100.665 6.155 -100.295 6.495 ;
        RECT -100.115 6.395 -99.945 6.720 ;
        RECT -95.135 6.720 -94.065 6.890 ;
        RECT -95.135 6.395 -94.965 6.720 ;
        RECT -100.115 6.225 -99.565 6.395 ;
        RECT -95.515 6.225 -94.965 6.395 ;
        RECT -94.785 6.155 -94.415 6.495 ;
        RECT -94.235 6.395 -94.065 6.720 ;
        RECT -91.095 6.720 -90.025 6.890 ;
        RECT -91.095 6.395 -90.925 6.720 ;
        RECT -94.235 6.215 -93.305 6.395 ;
        RECT -91.855 6.215 -90.925 6.395 ;
        RECT -90.745 6.155 -90.375 6.495 ;
        RECT -90.195 6.395 -90.025 6.720 ;
        RECT -85.215 6.720 -84.145 6.890 ;
        RECT -85.215 6.395 -85.045 6.720 ;
        RECT -90.195 6.225 -89.645 6.395 ;
        RECT -85.595 6.225 -85.045 6.395 ;
        RECT -84.865 6.155 -84.495 6.495 ;
        RECT -84.315 6.395 -84.145 6.720 ;
        RECT -81.175 6.720 -80.105 6.890 ;
        RECT -81.175 6.395 -81.005 6.720 ;
        RECT -84.315 6.215 -83.385 6.395 ;
        RECT -81.935 6.215 -81.005 6.395 ;
        RECT -80.825 6.155 -80.455 6.495 ;
        RECT -80.275 6.395 -80.105 6.720 ;
        RECT -75.295 6.720 -74.225 6.890 ;
        RECT -75.295 6.395 -75.125 6.720 ;
        RECT -80.275 6.225 -79.725 6.395 ;
        RECT -75.675 6.225 -75.125 6.395 ;
        RECT -74.945 6.155 -74.575 6.495 ;
        RECT -74.395 6.395 -74.225 6.720 ;
        RECT -71.255 6.720 -70.185 6.890 ;
        RECT -71.255 6.395 -71.085 6.720 ;
        RECT -74.395 6.215 -73.465 6.395 ;
        RECT -72.015 6.215 -71.085 6.395 ;
        RECT -70.905 6.155 -70.535 6.495 ;
        RECT -70.355 6.395 -70.185 6.720 ;
        RECT -65.375 6.720 -64.305 6.890 ;
        RECT -65.375 6.395 -65.205 6.720 ;
        RECT -70.355 6.225 -69.805 6.395 ;
        RECT -65.755 6.225 -65.205 6.395 ;
        RECT -65.025 6.155 -64.655 6.495 ;
        RECT -64.475 6.395 -64.305 6.720 ;
        RECT -61.335 6.720 -60.265 6.890 ;
        RECT -61.335 6.395 -61.165 6.720 ;
        RECT -64.475 6.215 -63.545 6.395 ;
        RECT -62.095 6.215 -61.165 6.395 ;
        RECT -60.985 6.155 -60.615 6.495 ;
        RECT -60.435 6.395 -60.265 6.720 ;
        RECT -55.455 6.720 -54.385 6.890 ;
        RECT -55.455 6.395 -55.285 6.720 ;
        RECT -60.435 6.225 -59.885 6.395 ;
        RECT -55.835 6.225 -55.285 6.395 ;
        RECT -55.105 6.155 -54.735 6.495 ;
        RECT -54.555 6.395 -54.385 6.720 ;
        RECT -51.415 6.720 -50.345 6.890 ;
        RECT -51.415 6.395 -51.245 6.720 ;
        RECT -54.555 6.215 -53.625 6.395 ;
        RECT -52.175 6.215 -51.245 6.395 ;
        RECT -51.065 6.155 -50.695 6.495 ;
        RECT -50.515 6.395 -50.345 6.720 ;
        RECT -45.535 6.720 -44.465 6.890 ;
        RECT -45.535 6.395 -45.365 6.720 ;
        RECT -50.515 6.225 -49.965 6.395 ;
        RECT -45.915 6.225 -45.365 6.395 ;
        RECT -45.185 6.155 -44.815 6.495 ;
        RECT -44.635 6.395 -44.465 6.720 ;
        RECT -41.495 6.720 -40.425 6.890 ;
        RECT -41.495 6.395 -41.325 6.720 ;
        RECT -44.635 6.215 -43.705 6.395 ;
        RECT -42.255 6.215 -41.325 6.395 ;
        RECT -41.145 6.155 -40.775 6.495 ;
        RECT -40.595 6.395 -40.425 6.720 ;
        RECT -35.615 6.720 -34.545 6.890 ;
        RECT -35.615 6.395 -35.445 6.720 ;
        RECT -40.595 6.225 -40.045 6.395 ;
        RECT -35.995 6.225 -35.445 6.395 ;
        RECT -35.265 6.155 -34.895 6.495 ;
        RECT -34.715 6.395 -34.545 6.720 ;
        RECT -31.575 6.720 -30.505 6.890 ;
        RECT -31.575 6.395 -31.405 6.720 ;
        RECT -34.715 6.215 -33.785 6.395 ;
        RECT -32.335 6.215 -31.405 6.395 ;
        RECT -31.225 6.155 -30.855 6.495 ;
        RECT -30.675 6.395 -30.505 6.720 ;
        RECT -25.695 6.720 -24.625 6.890 ;
        RECT -25.695 6.395 -25.525 6.720 ;
        RECT -30.675 6.225 -30.125 6.395 ;
        RECT -26.075 6.225 -25.525 6.395 ;
        RECT -25.345 6.155 -24.975 6.495 ;
        RECT -24.795 6.395 -24.625 6.720 ;
        RECT -21.655 6.720 -20.585 6.890 ;
        RECT -21.655 6.395 -21.485 6.720 ;
        RECT -24.795 6.215 -23.865 6.395 ;
        RECT -22.415 6.215 -21.485 6.395 ;
        RECT -21.305 6.155 -20.935 6.495 ;
        RECT -20.755 6.395 -20.585 6.720 ;
        RECT -15.775 6.720 -14.705 6.890 ;
        RECT -15.775 6.395 -15.605 6.720 ;
        RECT -20.755 6.225 -20.205 6.395 ;
        RECT -16.155 6.225 -15.605 6.395 ;
        RECT -15.425 6.155 -15.055 6.495 ;
        RECT -14.875 6.395 -14.705 6.720 ;
        RECT -11.735 6.720 -10.665 6.890 ;
        RECT -11.735 6.395 -11.565 6.720 ;
        RECT -14.875 6.215 -13.945 6.395 ;
        RECT -12.495 6.215 -11.565 6.395 ;
        RECT -11.385 6.155 -11.015 6.495 ;
        RECT -10.835 6.395 -10.665 6.720 ;
        RECT -5.855 6.720 -4.785 6.890 ;
        RECT -5.855 6.395 -5.685 6.720 ;
        RECT -10.835 6.225 -10.285 6.395 ;
        RECT -6.235 6.225 -5.685 6.395 ;
        RECT -5.505 6.155 -5.135 6.495 ;
        RECT -4.955 6.395 -4.785 6.720 ;
        RECT -1.815 6.720 -0.745 6.890 ;
        RECT -1.815 6.395 -1.645 6.720 ;
        RECT -4.955 6.215 -4.025 6.395 ;
        RECT -2.575 6.215 -1.645 6.395 ;
        RECT -1.465 6.155 -1.095 6.495 ;
        RECT -0.915 6.395 -0.745 6.720 ;
        RECT 4.065 6.720 5.135 6.890 ;
        RECT 4.065 6.395 4.235 6.720 ;
        RECT -0.915 6.225 -0.365 6.395 ;
        RECT 3.685 6.225 4.235 6.395 ;
        RECT 4.415 6.155 4.785 6.495 ;
        RECT 4.965 6.395 5.135 6.720 ;
        RECT 8.105 6.720 9.175 6.890 ;
        RECT 8.105 6.395 8.275 6.720 ;
        RECT 4.965 6.215 5.895 6.395 ;
        RECT 7.345 6.215 8.275 6.395 ;
        RECT 8.455 6.155 8.825 6.495 ;
        RECT 9.005 6.395 9.175 6.720 ;
        RECT 13.985 6.720 15.055 6.890 ;
        RECT 13.985 6.395 14.155 6.720 ;
        RECT 9.005 6.225 9.555 6.395 ;
        RECT 13.605 6.225 14.155 6.395 ;
        RECT 14.335 6.155 14.705 6.495 ;
        RECT 14.885 6.395 15.055 6.720 ;
        RECT 18.025 6.720 19.095 6.890 ;
        RECT 18.025 6.395 18.195 6.720 ;
        RECT 14.885 6.215 15.815 6.395 ;
        RECT 17.265 6.215 18.195 6.395 ;
        RECT 18.375 6.155 18.745 6.495 ;
        RECT 18.925 6.395 19.095 6.720 ;
        RECT 23.905 6.720 24.975 6.890 ;
        RECT 23.905 6.395 24.075 6.720 ;
        RECT 18.925 6.225 19.475 6.395 ;
        RECT 23.525 6.225 24.075 6.395 ;
        RECT 24.255 6.155 24.625 6.495 ;
        RECT 24.805 6.395 24.975 6.720 ;
        RECT 24.805 6.215 25.735 6.395 ;
        RECT -291.210 5.535 -289.370 5.705 ;
        RECT 24.850 5.535 26.690 5.705 ;
        RECT -291.125 4.810 -290.835 5.535 ;
        RECT -290.665 4.735 -290.355 5.535 ;
        RECT -290.150 4.735 -289.455 5.365 ;
        RECT -291.125 2.985 -290.835 4.150 ;
        RECT -290.150 4.135 -289.980 4.735 ;
        RECT -289.810 4.295 -289.475 4.545 ;
        RECT -287.115 4.385 -286.785 5.365 ;
        RECT -285.255 4.385 -284.925 5.365 ;
        RECT -282.585 4.735 -281.890 5.365 ;
        RECT -290.665 2.985 -290.385 4.125 ;
        RECT -290.215 3.155 -289.885 4.135 ;
        RECT -289.715 2.985 -289.455 4.125 ;
        RECT -287.525 3.975 -287.190 4.225 ;
        RECT -287.020 3.785 -286.850 4.385 ;
        RECT -287.545 3.155 -286.850 3.785 ;
        RECT -285.190 3.785 -285.020 4.385 ;
        RECT -282.565 4.295 -282.230 4.545 ;
        RECT -284.850 3.975 -284.515 4.225 ;
        RECT -282.060 4.135 -281.890 4.735 ;
        RECT -280.230 4.735 -279.535 5.365 ;
        RECT -280.230 4.135 -280.060 4.735 ;
        RECT -279.890 4.295 -279.555 4.545 ;
        RECT -277.195 4.385 -276.865 5.365 ;
        RECT -275.335 4.385 -275.005 5.365 ;
        RECT -272.665 4.735 -271.970 5.365 ;
        RECT -285.190 3.155 -284.495 3.785 ;
        RECT -282.155 3.155 -281.825 4.135 ;
        RECT -280.295 3.155 -279.965 4.135 ;
        RECT -277.605 3.975 -277.270 4.225 ;
        RECT -277.100 3.785 -276.930 4.385 ;
        RECT -277.625 3.155 -276.930 3.785 ;
        RECT -275.270 3.785 -275.100 4.385 ;
        RECT -272.645 4.295 -272.310 4.545 ;
        RECT -274.930 3.975 -274.595 4.225 ;
        RECT -272.140 4.135 -271.970 4.735 ;
        RECT -270.310 4.735 -269.615 5.365 ;
        RECT -270.310 4.135 -270.140 4.735 ;
        RECT -269.970 4.295 -269.635 4.545 ;
        RECT -267.275 4.385 -266.945 5.365 ;
        RECT -265.415 4.385 -265.085 5.365 ;
        RECT -262.745 4.735 -262.050 5.365 ;
        RECT -275.270 3.155 -274.575 3.785 ;
        RECT -272.235 3.155 -271.905 4.135 ;
        RECT -270.375 3.155 -270.045 4.135 ;
        RECT -267.685 3.975 -267.350 4.225 ;
        RECT -267.180 3.785 -267.010 4.385 ;
        RECT -267.705 3.155 -267.010 3.785 ;
        RECT -265.350 3.785 -265.180 4.385 ;
        RECT -262.725 4.295 -262.390 4.545 ;
        RECT -265.010 3.975 -264.675 4.225 ;
        RECT -262.220 4.135 -262.050 4.735 ;
        RECT -260.390 4.735 -259.695 5.365 ;
        RECT -260.390 4.135 -260.220 4.735 ;
        RECT -260.050 4.295 -259.715 4.545 ;
        RECT -257.355 4.385 -257.025 5.365 ;
        RECT -255.495 4.385 -255.165 5.365 ;
        RECT -252.825 4.735 -252.130 5.365 ;
        RECT -265.350 3.155 -264.655 3.785 ;
        RECT -262.315 3.155 -261.985 4.135 ;
        RECT -260.455 3.155 -260.125 4.135 ;
        RECT -257.765 3.975 -257.430 4.225 ;
        RECT -257.260 3.785 -257.090 4.385 ;
        RECT -257.785 3.155 -257.090 3.785 ;
        RECT -255.430 3.785 -255.260 4.385 ;
        RECT -252.805 4.295 -252.470 4.545 ;
        RECT -255.090 3.975 -254.755 4.225 ;
        RECT -252.300 4.135 -252.130 4.735 ;
        RECT -250.470 4.735 -249.775 5.365 ;
        RECT -250.470 4.135 -250.300 4.735 ;
        RECT -250.130 4.295 -249.795 4.545 ;
        RECT -247.435 4.385 -247.105 5.365 ;
        RECT -245.575 4.385 -245.245 5.365 ;
        RECT -242.905 4.735 -242.210 5.365 ;
        RECT -255.430 3.155 -254.735 3.785 ;
        RECT -252.395 3.155 -252.065 4.135 ;
        RECT -250.535 3.155 -250.205 4.135 ;
        RECT -247.845 3.975 -247.510 4.225 ;
        RECT -247.340 3.785 -247.170 4.385 ;
        RECT -247.865 3.155 -247.170 3.785 ;
        RECT -245.510 3.785 -245.340 4.385 ;
        RECT -242.885 4.295 -242.550 4.545 ;
        RECT -245.170 3.975 -244.835 4.225 ;
        RECT -242.380 4.135 -242.210 4.735 ;
        RECT -240.550 4.735 -239.855 5.365 ;
        RECT -240.550 4.135 -240.380 4.735 ;
        RECT -240.210 4.295 -239.875 4.545 ;
        RECT -237.515 4.385 -237.185 5.365 ;
        RECT -235.655 4.385 -235.325 5.365 ;
        RECT -232.985 4.735 -232.290 5.365 ;
        RECT -245.510 3.155 -244.815 3.785 ;
        RECT -242.475 3.155 -242.145 4.135 ;
        RECT -240.615 3.155 -240.285 4.135 ;
        RECT -237.925 3.975 -237.590 4.225 ;
        RECT -237.420 3.785 -237.250 4.385 ;
        RECT -237.945 3.155 -237.250 3.785 ;
        RECT -235.590 3.785 -235.420 4.385 ;
        RECT -232.965 4.295 -232.630 4.545 ;
        RECT -235.250 3.975 -234.915 4.225 ;
        RECT -232.460 4.135 -232.290 4.735 ;
        RECT -230.630 4.735 -229.935 5.365 ;
        RECT -230.630 4.135 -230.460 4.735 ;
        RECT -230.290 4.295 -229.955 4.545 ;
        RECT -227.595 4.385 -227.265 5.365 ;
        RECT -225.735 4.385 -225.405 5.365 ;
        RECT -223.065 4.735 -222.370 5.365 ;
        RECT -235.590 3.155 -234.895 3.785 ;
        RECT -232.555 3.155 -232.225 4.135 ;
        RECT -230.695 3.155 -230.365 4.135 ;
        RECT -228.005 3.975 -227.670 4.225 ;
        RECT -227.500 3.785 -227.330 4.385 ;
        RECT -228.025 3.155 -227.330 3.785 ;
        RECT -225.670 3.785 -225.500 4.385 ;
        RECT -223.045 4.295 -222.710 4.545 ;
        RECT -225.330 3.975 -224.995 4.225 ;
        RECT -222.540 4.135 -222.370 4.735 ;
        RECT -220.710 4.735 -220.015 5.365 ;
        RECT -220.710 4.135 -220.540 4.735 ;
        RECT -220.370 4.295 -220.035 4.545 ;
        RECT -217.675 4.385 -217.345 5.365 ;
        RECT -215.815 4.385 -215.485 5.365 ;
        RECT -213.145 4.735 -212.450 5.365 ;
        RECT -225.670 3.155 -224.975 3.785 ;
        RECT -222.635 3.155 -222.305 4.135 ;
        RECT -220.775 3.155 -220.445 4.135 ;
        RECT -218.085 3.975 -217.750 4.225 ;
        RECT -217.580 3.785 -217.410 4.385 ;
        RECT -218.105 3.155 -217.410 3.785 ;
        RECT -215.750 3.785 -215.580 4.385 ;
        RECT -213.125 4.295 -212.790 4.545 ;
        RECT -215.410 3.975 -215.075 4.225 ;
        RECT -212.620 4.135 -212.450 4.735 ;
        RECT -210.790 4.735 -210.095 5.365 ;
        RECT -210.790 4.135 -210.620 4.735 ;
        RECT -210.450 4.295 -210.115 4.545 ;
        RECT -207.755 4.385 -207.425 5.365 ;
        RECT -205.895 4.385 -205.565 5.365 ;
        RECT -203.225 4.735 -202.530 5.365 ;
        RECT -215.750 3.155 -215.055 3.785 ;
        RECT -212.715 3.155 -212.385 4.135 ;
        RECT -210.855 3.155 -210.525 4.135 ;
        RECT -208.165 3.975 -207.830 4.225 ;
        RECT -207.660 3.785 -207.490 4.385 ;
        RECT -208.185 3.155 -207.490 3.785 ;
        RECT -205.830 3.785 -205.660 4.385 ;
        RECT -203.205 4.295 -202.870 4.545 ;
        RECT -205.490 3.975 -205.155 4.225 ;
        RECT -202.700 4.135 -202.530 4.735 ;
        RECT -200.870 4.735 -200.175 5.365 ;
        RECT -200.870 4.135 -200.700 4.735 ;
        RECT -200.530 4.295 -200.195 4.545 ;
        RECT -197.835 4.385 -197.505 5.365 ;
        RECT -195.975 4.385 -195.645 5.365 ;
        RECT -193.305 4.735 -192.610 5.365 ;
        RECT -205.830 3.155 -205.135 3.785 ;
        RECT -202.795 3.155 -202.465 4.135 ;
        RECT -200.935 3.155 -200.605 4.135 ;
        RECT -198.245 3.975 -197.910 4.225 ;
        RECT -197.740 3.785 -197.570 4.385 ;
        RECT -198.265 3.155 -197.570 3.785 ;
        RECT -195.910 3.785 -195.740 4.385 ;
        RECT -193.285 4.295 -192.950 4.545 ;
        RECT -195.570 3.975 -195.235 4.225 ;
        RECT -192.780 4.135 -192.610 4.735 ;
        RECT -190.950 4.735 -190.255 5.365 ;
        RECT -190.950 4.135 -190.780 4.735 ;
        RECT -190.610 4.295 -190.275 4.545 ;
        RECT -187.915 4.385 -187.585 5.365 ;
        RECT -186.055 4.385 -185.725 5.365 ;
        RECT -183.385 4.735 -182.690 5.365 ;
        RECT -195.910 3.155 -195.215 3.785 ;
        RECT -192.875 3.155 -192.545 4.135 ;
        RECT -191.015 3.155 -190.685 4.135 ;
        RECT -188.325 3.975 -187.990 4.225 ;
        RECT -187.820 3.785 -187.650 4.385 ;
        RECT -188.345 3.155 -187.650 3.785 ;
        RECT -185.990 3.785 -185.820 4.385 ;
        RECT -183.365 4.295 -183.030 4.545 ;
        RECT -185.650 3.975 -185.315 4.225 ;
        RECT -182.860 4.135 -182.690 4.735 ;
        RECT -181.030 4.735 -180.335 5.365 ;
        RECT -181.030 4.135 -180.860 4.735 ;
        RECT -180.690 4.295 -180.355 4.545 ;
        RECT -177.995 4.385 -177.665 5.365 ;
        RECT -176.135 4.385 -175.805 5.365 ;
        RECT -173.465 4.735 -172.770 5.365 ;
        RECT -185.990 3.155 -185.295 3.785 ;
        RECT -182.955 3.155 -182.625 4.135 ;
        RECT -181.095 3.155 -180.765 4.135 ;
        RECT -178.405 3.975 -178.070 4.225 ;
        RECT -177.900 3.785 -177.730 4.385 ;
        RECT -178.425 3.155 -177.730 3.785 ;
        RECT -176.070 3.785 -175.900 4.385 ;
        RECT -173.445 4.295 -173.110 4.545 ;
        RECT -175.730 3.975 -175.395 4.225 ;
        RECT -172.940 4.135 -172.770 4.735 ;
        RECT -171.110 4.735 -170.415 5.365 ;
        RECT -171.110 4.135 -170.940 4.735 ;
        RECT -170.770 4.295 -170.435 4.545 ;
        RECT -168.075 4.385 -167.745 5.365 ;
        RECT -166.215 4.385 -165.885 5.365 ;
        RECT -163.545 4.735 -162.850 5.365 ;
        RECT -176.070 3.155 -175.375 3.785 ;
        RECT -173.035 3.155 -172.705 4.135 ;
        RECT -171.175 3.155 -170.845 4.135 ;
        RECT -168.485 3.975 -168.150 4.225 ;
        RECT -167.980 3.785 -167.810 4.385 ;
        RECT -168.505 3.155 -167.810 3.785 ;
        RECT -166.150 3.785 -165.980 4.385 ;
        RECT -163.525 4.295 -163.190 4.545 ;
        RECT -165.810 3.975 -165.475 4.225 ;
        RECT -163.020 4.135 -162.850 4.735 ;
        RECT -161.190 4.735 -160.495 5.365 ;
        RECT -161.190 4.135 -161.020 4.735 ;
        RECT -160.850 4.295 -160.515 4.545 ;
        RECT -158.155 4.385 -157.825 5.365 ;
        RECT -156.295 4.385 -155.965 5.365 ;
        RECT -153.625 4.735 -152.930 5.365 ;
        RECT -166.150 3.155 -165.455 3.785 ;
        RECT -163.115 3.155 -162.785 4.135 ;
        RECT -161.255 3.155 -160.925 4.135 ;
        RECT -158.565 3.975 -158.230 4.225 ;
        RECT -158.060 3.785 -157.890 4.385 ;
        RECT -158.585 3.155 -157.890 3.785 ;
        RECT -156.230 3.785 -156.060 4.385 ;
        RECT -153.605 4.295 -153.270 4.545 ;
        RECT -155.890 3.975 -155.555 4.225 ;
        RECT -153.100 4.135 -152.930 4.735 ;
        RECT -151.270 4.735 -150.575 5.365 ;
        RECT -151.270 4.135 -151.100 4.735 ;
        RECT -150.930 4.295 -150.595 4.545 ;
        RECT -148.235 4.385 -147.905 5.365 ;
        RECT -146.375 4.385 -146.045 5.365 ;
        RECT -143.705 4.735 -143.010 5.365 ;
        RECT -156.230 3.155 -155.535 3.785 ;
        RECT -153.195 3.155 -152.865 4.135 ;
        RECT -151.335 3.155 -151.005 4.135 ;
        RECT -148.645 3.975 -148.310 4.225 ;
        RECT -148.140 3.785 -147.970 4.385 ;
        RECT -148.665 3.155 -147.970 3.785 ;
        RECT -146.310 3.785 -146.140 4.385 ;
        RECT -143.685 4.295 -143.350 4.545 ;
        RECT -145.970 3.975 -145.635 4.225 ;
        RECT -143.180 4.135 -143.010 4.735 ;
        RECT -141.350 4.735 -140.655 5.365 ;
        RECT -141.350 4.135 -141.180 4.735 ;
        RECT -141.010 4.295 -140.675 4.545 ;
        RECT -138.315 4.385 -137.985 5.365 ;
        RECT -136.455 4.385 -136.125 5.365 ;
        RECT -133.785 4.735 -133.090 5.365 ;
        RECT -146.310 3.155 -145.615 3.785 ;
        RECT -143.275 3.155 -142.945 4.135 ;
        RECT -141.415 3.155 -141.085 4.135 ;
        RECT -138.725 3.975 -138.390 4.225 ;
        RECT -138.220 3.785 -138.050 4.385 ;
        RECT -138.745 3.155 -138.050 3.785 ;
        RECT -136.390 3.785 -136.220 4.385 ;
        RECT -133.765 4.295 -133.430 4.545 ;
        RECT -136.050 3.975 -135.715 4.225 ;
        RECT -133.260 4.135 -133.090 4.735 ;
        RECT -131.430 4.735 -130.735 5.365 ;
        RECT -131.430 4.135 -131.260 4.735 ;
        RECT -131.090 4.295 -130.755 4.545 ;
        RECT -128.395 4.385 -128.065 5.365 ;
        RECT -126.535 4.385 -126.205 5.365 ;
        RECT -123.865 4.735 -123.170 5.365 ;
        RECT -136.390 3.155 -135.695 3.785 ;
        RECT -133.355 3.155 -133.025 4.135 ;
        RECT -131.495 3.155 -131.165 4.135 ;
        RECT -128.805 3.975 -128.470 4.225 ;
        RECT -128.300 3.785 -128.130 4.385 ;
        RECT -128.825 3.155 -128.130 3.785 ;
        RECT -126.470 3.785 -126.300 4.385 ;
        RECT -123.845 4.295 -123.510 4.545 ;
        RECT -126.130 3.975 -125.795 4.225 ;
        RECT -123.340 4.135 -123.170 4.735 ;
        RECT -121.510 4.735 -120.815 5.365 ;
        RECT -121.510 4.135 -121.340 4.735 ;
        RECT -121.170 4.295 -120.835 4.545 ;
        RECT -118.475 4.385 -118.145 5.365 ;
        RECT -116.615 4.385 -116.285 5.365 ;
        RECT -113.945 4.735 -113.250 5.365 ;
        RECT -126.470 3.155 -125.775 3.785 ;
        RECT -123.435 3.155 -123.105 4.135 ;
        RECT -121.575 3.155 -121.245 4.135 ;
        RECT -118.885 3.975 -118.550 4.225 ;
        RECT -118.380 3.785 -118.210 4.385 ;
        RECT -118.905 3.155 -118.210 3.785 ;
        RECT -116.550 3.785 -116.380 4.385 ;
        RECT -113.925 4.295 -113.590 4.545 ;
        RECT -116.210 3.975 -115.875 4.225 ;
        RECT -113.420 4.135 -113.250 4.735 ;
        RECT -111.590 4.735 -110.895 5.365 ;
        RECT -111.590 4.135 -111.420 4.735 ;
        RECT -111.250 4.295 -110.915 4.545 ;
        RECT -108.555 4.385 -108.225 5.365 ;
        RECT -106.695 4.385 -106.365 5.365 ;
        RECT -104.025 4.735 -103.330 5.365 ;
        RECT -116.550 3.155 -115.855 3.785 ;
        RECT -113.515 3.155 -113.185 4.135 ;
        RECT -111.655 3.155 -111.325 4.135 ;
        RECT -108.965 3.975 -108.630 4.225 ;
        RECT -108.460 3.785 -108.290 4.385 ;
        RECT -108.985 3.155 -108.290 3.785 ;
        RECT -106.630 3.785 -106.460 4.385 ;
        RECT -104.005 4.295 -103.670 4.545 ;
        RECT -106.290 3.975 -105.955 4.225 ;
        RECT -103.500 4.135 -103.330 4.735 ;
        RECT -101.670 4.735 -100.975 5.365 ;
        RECT -101.670 4.135 -101.500 4.735 ;
        RECT -101.330 4.295 -100.995 4.545 ;
        RECT -98.635 4.385 -98.305 5.365 ;
        RECT -96.775 4.385 -96.445 5.365 ;
        RECT -94.105 4.735 -93.410 5.365 ;
        RECT -106.630 3.155 -105.935 3.785 ;
        RECT -103.595 3.155 -103.265 4.135 ;
        RECT -101.735 3.155 -101.405 4.135 ;
        RECT -99.045 3.975 -98.710 4.225 ;
        RECT -98.540 3.785 -98.370 4.385 ;
        RECT -99.065 3.155 -98.370 3.785 ;
        RECT -96.710 3.785 -96.540 4.385 ;
        RECT -94.085 4.295 -93.750 4.545 ;
        RECT -96.370 3.975 -96.035 4.225 ;
        RECT -93.580 4.135 -93.410 4.735 ;
        RECT -91.750 4.735 -91.055 5.365 ;
        RECT -91.750 4.135 -91.580 4.735 ;
        RECT -91.410 4.295 -91.075 4.545 ;
        RECT -88.715 4.385 -88.385 5.365 ;
        RECT -86.855 4.385 -86.525 5.365 ;
        RECT -84.185 4.735 -83.490 5.365 ;
        RECT -96.710 3.155 -96.015 3.785 ;
        RECT -93.675 3.155 -93.345 4.135 ;
        RECT -91.815 3.155 -91.485 4.135 ;
        RECT -89.125 3.975 -88.790 4.225 ;
        RECT -88.620 3.785 -88.450 4.385 ;
        RECT -89.145 3.155 -88.450 3.785 ;
        RECT -86.790 3.785 -86.620 4.385 ;
        RECT -84.165 4.295 -83.830 4.545 ;
        RECT -86.450 3.975 -86.115 4.225 ;
        RECT -83.660 4.135 -83.490 4.735 ;
        RECT -81.830 4.735 -81.135 5.365 ;
        RECT -81.830 4.135 -81.660 4.735 ;
        RECT -81.490 4.295 -81.155 4.545 ;
        RECT -78.795 4.385 -78.465 5.365 ;
        RECT -76.935 4.385 -76.605 5.365 ;
        RECT -74.265 4.735 -73.570 5.365 ;
        RECT -86.790 3.155 -86.095 3.785 ;
        RECT -83.755 3.155 -83.425 4.135 ;
        RECT -81.895 3.155 -81.565 4.135 ;
        RECT -79.205 3.975 -78.870 4.225 ;
        RECT -78.700 3.785 -78.530 4.385 ;
        RECT -79.225 3.155 -78.530 3.785 ;
        RECT -76.870 3.785 -76.700 4.385 ;
        RECT -74.245 4.295 -73.910 4.545 ;
        RECT -76.530 3.975 -76.195 4.225 ;
        RECT -73.740 4.135 -73.570 4.735 ;
        RECT -71.910 4.735 -71.215 5.365 ;
        RECT -71.910 4.135 -71.740 4.735 ;
        RECT -71.570 4.295 -71.235 4.545 ;
        RECT -68.875 4.385 -68.545 5.365 ;
        RECT -67.015 4.385 -66.685 5.365 ;
        RECT -64.345 4.735 -63.650 5.365 ;
        RECT -76.870 3.155 -76.175 3.785 ;
        RECT -73.835 3.155 -73.505 4.135 ;
        RECT -71.975 3.155 -71.645 4.135 ;
        RECT -69.285 3.975 -68.950 4.225 ;
        RECT -68.780 3.785 -68.610 4.385 ;
        RECT -69.305 3.155 -68.610 3.785 ;
        RECT -66.950 3.785 -66.780 4.385 ;
        RECT -64.325 4.295 -63.990 4.545 ;
        RECT -66.610 3.975 -66.275 4.225 ;
        RECT -63.820 4.135 -63.650 4.735 ;
        RECT -61.990 4.735 -61.295 5.365 ;
        RECT -61.990 4.135 -61.820 4.735 ;
        RECT -61.650 4.295 -61.315 4.545 ;
        RECT -58.955 4.385 -58.625 5.365 ;
        RECT -57.095 4.385 -56.765 5.365 ;
        RECT -54.425 4.735 -53.730 5.365 ;
        RECT -66.950 3.155 -66.255 3.785 ;
        RECT -63.915 3.155 -63.585 4.135 ;
        RECT -62.055 3.155 -61.725 4.135 ;
        RECT -59.365 3.975 -59.030 4.225 ;
        RECT -58.860 3.785 -58.690 4.385 ;
        RECT -59.385 3.155 -58.690 3.785 ;
        RECT -57.030 3.785 -56.860 4.385 ;
        RECT -54.405 4.295 -54.070 4.545 ;
        RECT -56.690 3.975 -56.355 4.225 ;
        RECT -53.900 4.135 -53.730 4.735 ;
        RECT -52.070 4.735 -51.375 5.365 ;
        RECT -52.070 4.135 -51.900 4.735 ;
        RECT -51.730 4.295 -51.395 4.545 ;
        RECT -49.035 4.385 -48.705 5.365 ;
        RECT -47.175 4.385 -46.845 5.365 ;
        RECT -44.505 4.735 -43.810 5.365 ;
        RECT -57.030 3.155 -56.335 3.785 ;
        RECT -53.995 3.155 -53.665 4.135 ;
        RECT -52.135 3.155 -51.805 4.135 ;
        RECT -49.445 3.975 -49.110 4.225 ;
        RECT -48.940 3.785 -48.770 4.385 ;
        RECT -49.465 3.155 -48.770 3.785 ;
        RECT -47.110 3.785 -46.940 4.385 ;
        RECT -44.485 4.295 -44.150 4.545 ;
        RECT -46.770 3.975 -46.435 4.225 ;
        RECT -43.980 4.135 -43.810 4.735 ;
        RECT -42.150 4.735 -41.455 5.365 ;
        RECT -42.150 4.135 -41.980 4.735 ;
        RECT -41.810 4.295 -41.475 4.545 ;
        RECT -39.115 4.385 -38.785 5.365 ;
        RECT -37.255 4.385 -36.925 5.365 ;
        RECT -34.585 4.735 -33.890 5.365 ;
        RECT -47.110 3.155 -46.415 3.785 ;
        RECT -44.075 3.155 -43.745 4.135 ;
        RECT -42.215 3.155 -41.885 4.135 ;
        RECT -39.525 3.975 -39.190 4.225 ;
        RECT -39.020 3.785 -38.850 4.385 ;
        RECT -39.545 3.155 -38.850 3.785 ;
        RECT -37.190 3.785 -37.020 4.385 ;
        RECT -34.565 4.295 -34.230 4.545 ;
        RECT -36.850 3.975 -36.515 4.225 ;
        RECT -34.060 4.135 -33.890 4.735 ;
        RECT -32.230 4.735 -31.535 5.365 ;
        RECT -32.230 4.135 -32.060 4.735 ;
        RECT -31.890 4.295 -31.555 4.545 ;
        RECT -29.195 4.385 -28.865 5.365 ;
        RECT -27.335 4.385 -27.005 5.365 ;
        RECT -24.665 4.735 -23.970 5.365 ;
        RECT -37.190 3.155 -36.495 3.785 ;
        RECT -34.155 3.155 -33.825 4.135 ;
        RECT -32.295 3.155 -31.965 4.135 ;
        RECT -29.605 3.975 -29.270 4.225 ;
        RECT -29.100 3.785 -28.930 4.385 ;
        RECT -29.625 3.155 -28.930 3.785 ;
        RECT -27.270 3.785 -27.100 4.385 ;
        RECT -24.645 4.295 -24.310 4.545 ;
        RECT -26.930 3.975 -26.595 4.225 ;
        RECT -24.140 4.135 -23.970 4.735 ;
        RECT -22.310 4.735 -21.615 5.365 ;
        RECT -22.310 4.135 -22.140 4.735 ;
        RECT -21.970 4.295 -21.635 4.545 ;
        RECT -19.275 4.385 -18.945 5.365 ;
        RECT -17.415 4.385 -17.085 5.365 ;
        RECT -14.745 4.735 -14.050 5.365 ;
        RECT -27.270 3.155 -26.575 3.785 ;
        RECT -24.235 3.155 -23.905 4.135 ;
        RECT -22.375 3.155 -22.045 4.135 ;
        RECT -19.685 3.975 -19.350 4.225 ;
        RECT -19.180 3.785 -19.010 4.385 ;
        RECT -19.705 3.155 -19.010 3.785 ;
        RECT -17.350 3.785 -17.180 4.385 ;
        RECT -14.725 4.295 -14.390 4.545 ;
        RECT -17.010 3.975 -16.675 4.225 ;
        RECT -14.220 4.135 -14.050 4.735 ;
        RECT -12.390 4.735 -11.695 5.365 ;
        RECT -12.390 4.135 -12.220 4.735 ;
        RECT -12.050 4.295 -11.715 4.545 ;
        RECT -9.355 4.385 -9.025 5.365 ;
        RECT -7.495 4.385 -7.165 5.365 ;
        RECT -4.825 4.735 -4.130 5.365 ;
        RECT -17.350 3.155 -16.655 3.785 ;
        RECT -14.315 3.155 -13.985 4.135 ;
        RECT -12.455 3.155 -12.125 4.135 ;
        RECT -9.765 3.975 -9.430 4.225 ;
        RECT -9.260 3.785 -9.090 4.385 ;
        RECT -9.785 3.155 -9.090 3.785 ;
        RECT -7.430 3.785 -7.260 4.385 ;
        RECT -4.805 4.295 -4.470 4.545 ;
        RECT -7.090 3.975 -6.755 4.225 ;
        RECT -4.300 4.135 -4.130 4.735 ;
        RECT -2.470 4.735 -1.775 5.365 ;
        RECT -2.470 4.135 -2.300 4.735 ;
        RECT -2.130 4.295 -1.795 4.545 ;
        RECT 0.565 4.385 0.895 5.365 ;
        RECT 2.425 4.385 2.755 5.365 ;
        RECT 5.095 4.735 5.790 5.365 ;
        RECT -7.430 3.155 -6.735 3.785 ;
        RECT -4.395 3.155 -4.065 4.135 ;
        RECT -2.535 3.155 -2.205 4.135 ;
        RECT 0.155 3.975 0.490 4.225 ;
        RECT 0.660 3.785 0.830 4.385 ;
        RECT 0.135 3.155 0.830 3.785 ;
        RECT 2.490 3.785 2.660 4.385 ;
        RECT 5.115 4.295 5.450 4.545 ;
        RECT 2.830 3.975 3.165 4.225 ;
        RECT 5.620 4.135 5.790 4.735 ;
        RECT 7.450 4.735 8.145 5.365 ;
        RECT 7.450 4.135 7.620 4.735 ;
        RECT 7.790 4.295 8.125 4.545 ;
        RECT 10.485 4.385 10.815 5.365 ;
        RECT 12.345 4.385 12.675 5.365 ;
        RECT 15.015 4.735 15.710 5.365 ;
        RECT 2.490 3.155 3.185 3.785 ;
        RECT 5.525 3.155 5.855 4.135 ;
        RECT 7.385 3.155 7.715 4.135 ;
        RECT 10.075 3.975 10.410 4.225 ;
        RECT 10.580 3.785 10.750 4.385 ;
        RECT 10.055 3.155 10.750 3.785 ;
        RECT 12.410 3.785 12.580 4.385 ;
        RECT 15.035 4.295 15.370 4.545 ;
        RECT 12.750 3.975 13.085 4.225 ;
        RECT 15.540 4.135 15.710 4.735 ;
        RECT 17.370 4.735 18.065 5.365 ;
        RECT 17.370 4.135 17.540 4.735 ;
        RECT 17.710 4.295 18.045 4.545 ;
        RECT 20.405 4.385 20.735 5.365 ;
        RECT 22.265 4.385 22.595 5.365 ;
        RECT 24.935 4.735 25.630 5.365 ;
        RECT 25.835 4.735 26.145 5.535 ;
        RECT 26.315 4.810 26.605 5.535 ;
        RECT 12.410 3.155 13.105 3.785 ;
        RECT 15.445 3.155 15.775 4.135 ;
        RECT 17.305 3.155 17.635 4.135 ;
        RECT 19.995 3.975 20.330 4.225 ;
        RECT 20.500 3.785 20.670 4.385 ;
        RECT 19.975 3.155 20.670 3.785 ;
        RECT 22.330 3.785 22.500 4.385 ;
        RECT 24.955 4.295 25.290 4.545 ;
        RECT 22.670 3.975 23.005 4.225 ;
        RECT 25.460 4.135 25.630 4.735 ;
        RECT 22.330 3.155 23.025 3.785 ;
        RECT 25.365 3.155 25.695 4.135 ;
        RECT -291.210 2.815 -289.370 2.985 ;
        RECT -289.825 1.430 -289.535 2.140 ;
        RECT -289.295 1.945 -289.125 2.470 ;
        RECT -288.955 2.125 -288.405 2.295 ;
        RECT -289.295 1.615 -288.745 1.945 ;
        RECT -288.575 1.800 -288.405 2.125 ;
        RECT -288.225 2.025 -287.855 2.365 ;
        RECT -287.675 2.125 -286.745 2.305 ;
        RECT -285.295 2.125 -284.365 2.305 ;
        RECT -287.675 1.800 -287.505 2.125 ;
        RECT -288.575 1.630 -287.505 1.800 ;
        RECT -284.535 1.800 -284.365 2.125 ;
        RECT -284.185 2.025 -283.815 2.365 ;
        RECT -283.635 2.125 -283.085 2.295 ;
        RECT -279.035 2.125 -278.485 2.295 ;
        RECT -283.635 1.800 -283.465 2.125 ;
        RECT -284.535 1.630 -283.465 1.800 ;
        RECT -278.655 1.800 -278.485 2.125 ;
        RECT -278.305 2.025 -277.935 2.365 ;
        RECT -277.755 2.125 -276.825 2.305 ;
        RECT -275.375 2.125 -274.445 2.305 ;
        RECT -277.755 1.800 -277.585 2.125 ;
        RECT -278.655 1.630 -277.585 1.800 ;
        RECT -274.615 1.800 -274.445 2.125 ;
        RECT -274.265 2.025 -273.895 2.365 ;
        RECT -273.715 2.125 -273.165 2.295 ;
        RECT -269.115 2.125 -268.565 2.295 ;
        RECT -273.715 1.800 -273.545 2.125 ;
        RECT -274.615 1.630 -273.545 1.800 ;
        RECT -268.735 1.800 -268.565 2.125 ;
        RECT -268.385 2.025 -268.015 2.365 ;
        RECT -267.835 2.125 -266.905 2.305 ;
        RECT -265.455 2.125 -264.525 2.305 ;
        RECT -267.835 1.800 -267.665 2.125 ;
        RECT -268.735 1.630 -267.665 1.800 ;
        RECT -264.695 1.800 -264.525 2.125 ;
        RECT -264.345 2.025 -263.975 2.365 ;
        RECT -263.795 2.125 -263.245 2.295 ;
        RECT -259.195 2.125 -258.645 2.295 ;
        RECT -263.795 1.800 -263.625 2.125 ;
        RECT -264.695 1.630 -263.625 1.800 ;
        RECT -258.815 1.800 -258.645 2.125 ;
        RECT -258.465 2.025 -258.095 2.365 ;
        RECT -257.915 2.125 -256.985 2.305 ;
        RECT -255.535 2.125 -254.605 2.305 ;
        RECT -257.915 1.800 -257.745 2.125 ;
        RECT -258.815 1.630 -257.745 1.800 ;
        RECT -254.775 1.800 -254.605 2.125 ;
        RECT -254.425 2.025 -254.055 2.365 ;
        RECT -253.875 2.125 -253.325 2.295 ;
        RECT -249.275 2.125 -248.725 2.295 ;
        RECT -253.875 1.800 -253.705 2.125 ;
        RECT -254.775 1.630 -253.705 1.800 ;
        RECT -248.895 1.800 -248.725 2.125 ;
        RECT -248.545 2.025 -248.175 2.365 ;
        RECT -247.995 2.125 -247.065 2.305 ;
        RECT -245.615 2.125 -244.685 2.305 ;
        RECT -247.995 1.800 -247.825 2.125 ;
        RECT -248.895 1.630 -247.825 1.800 ;
        RECT -244.855 1.800 -244.685 2.125 ;
        RECT -244.505 2.025 -244.135 2.365 ;
        RECT -243.955 2.125 -243.405 2.295 ;
        RECT -239.355 2.125 -238.805 2.295 ;
        RECT -243.955 1.800 -243.785 2.125 ;
        RECT -244.855 1.630 -243.785 1.800 ;
        RECT -238.975 1.800 -238.805 2.125 ;
        RECT -238.625 2.025 -238.255 2.365 ;
        RECT -238.075 2.125 -237.145 2.305 ;
        RECT -235.695 2.125 -234.765 2.305 ;
        RECT -238.075 1.800 -237.905 2.125 ;
        RECT -238.975 1.630 -237.905 1.800 ;
        RECT -234.935 1.800 -234.765 2.125 ;
        RECT -234.585 2.025 -234.215 2.365 ;
        RECT -234.035 2.125 -233.485 2.295 ;
        RECT -229.435 2.125 -228.885 2.295 ;
        RECT -234.035 1.800 -233.865 2.125 ;
        RECT -234.935 1.630 -233.865 1.800 ;
        RECT -229.055 1.800 -228.885 2.125 ;
        RECT -228.705 2.025 -228.335 2.365 ;
        RECT -228.155 2.125 -227.225 2.305 ;
        RECT -225.775 2.125 -224.845 2.305 ;
        RECT -228.155 1.800 -227.985 2.125 ;
        RECT -229.055 1.630 -227.985 1.800 ;
        RECT -225.015 1.800 -224.845 2.125 ;
        RECT -224.665 2.025 -224.295 2.365 ;
        RECT -224.115 2.125 -223.565 2.295 ;
        RECT -219.515 2.125 -218.965 2.295 ;
        RECT -224.115 1.800 -223.945 2.125 ;
        RECT -225.015 1.630 -223.945 1.800 ;
        RECT -219.135 1.800 -218.965 2.125 ;
        RECT -218.785 2.025 -218.415 2.365 ;
        RECT -218.235 2.125 -217.305 2.305 ;
        RECT -215.855 2.125 -214.925 2.305 ;
        RECT -218.235 1.800 -218.065 2.125 ;
        RECT -219.135 1.630 -218.065 1.800 ;
        RECT -215.095 1.800 -214.925 2.125 ;
        RECT -214.745 2.025 -214.375 2.365 ;
        RECT -214.195 2.125 -213.645 2.295 ;
        RECT -209.595 2.125 -209.045 2.295 ;
        RECT -214.195 1.800 -214.025 2.125 ;
        RECT -215.095 1.630 -214.025 1.800 ;
        RECT -209.215 1.800 -209.045 2.125 ;
        RECT -208.865 2.025 -208.495 2.365 ;
        RECT -208.315 2.125 -207.385 2.305 ;
        RECT -205.935 2.125 -205.005 2.305 ;
        RECT -208.315 1.800 -208.145 2.125 ;
        RECT -209.215 1.630 -208.145 1.800 ;
        RECT -205.175 1.800 -205.005 2.125 ;
        RECT -204.825 2.025 -204.455 2.365 ;
        RECT -204.275 2.125 -203.725 2.295 ;
        RECT -199.675 2.125 -199.125 2.295 ;
        RECT -204.275 1.800 -204.105 2.125 ;
        RECT -205.175 1.630 -204.105 1.800 ;
        RECT -199.295 1.800 -199.125 2.125 ;
        RECT -198.945 2.025 -198.575 2.365 ;
        RECT -198.395 2.125 -197.465 2.305 ;
        RECT -196.015 2.125 -195.085 2.305 ;
        RECT -198.395 1.800 -198.225 2.125 ;
        RECT -199.295 1.630 -198.225 1.800 ;
        RECT -195.255 1.800 -195.085 2.125 ;
        RECT -194.905 2.025 -194.535 2.365 ;
        RECT -194.355 2.125 -193.805 2.295 ;
        RECT -189.755 2.125 -189.205 2.295 ;
        RECT -194.355 1.800 -194.185 2.125 ;
        RECT -195.255 1.630 -194.185 1.800 ;
        RECT -189.375 1.800 -189.205 2.125 ;
        RECT -189.025 2.025 -188.655 2.365 ;
        RECT -188.475 2.125 -187.545 2.305 ;
        RECT -186.095 2.125 -185.165 2.305 ;
        RECT -188.475 1.800 -188.305 2.125 ;
        RECT -189.375 1.630 -188.305 1.800 ;
        RECT -185.335 1.800 -185.165 2.125 ;
        RECT -184.985 2.025 -184.615 2.365 ;
        RECT -184.435 2.125 -183.885 2.295 ;
        RECT -179.835 2.125 -179.285 2.295 ;
        RECT -184.435 1.800 -184.265 2.125 ;
        RECT -185.335 1.630 -184.265 1.800 ;
        RECT -179.455 1.800 -179.285 2.125 ;
        RECT -179.105 2.025 -178.735 2.365 ;
        RECT -178.555 2.125 -177.625 2.305 ;
        RECT -176.175 2.125 -175.245 2.305 ;
        RECT -178.555 1.800 -178.385 2.125 ;
        RECT -179.455 1.630 -178.385 1.800 ;
        RECT -175.415 1.800 -175.245 2.125 ;
        RECT -175.065 2.025 -174.695 2.365 ;
        RECT -174.515 2.125 -173.965 2.295 ;
        RECT -169.915 2.125 -169.365 2.295 ;
        RECT -174.515 1.800 -174.345 2.125 ;
        RECT -175.415 1.630 -174.345 1.800 ;
        RECT -169.535 1.800 -169.365 2.125 ;
        RECT -169.185 2.025 -168.815 2.365 ;
        RECT -168.635 2.125 -167.705 2.305 ;
        RECT -166.255 2.125 -165.325 2.305 ;
        RECT -168.635 1.800 -168.465 2.125 ;
        RECT -169.535 1.630 -168.465 1.800 ;
        RECT -165.495 1.800 -165.325 2.125 ;
        RECT -165.145 2.025 -164.775 2.365 ;
        RECT -164.595 2.125 -164.045 2.295 ;
        RECT -159.995 2.125 -159.445 2.295 ;
        RECT -164.595 1.800 -164.425 2.125 ;
        RECT -165.495 1.630 -164.425 1.800 ;
        RECT -159.615 1.800 -159.445 2.125 ;
        RECT -159.265 2.025 -158.895 2.365 ;
        RECT -158.715 2.125 -157.785 2.305 ;
        RECT -156.335 2.125 -155.405 2.305 ;
        RECT -158.715 1.800 -158.545 2.125 ;
        RECT -159.615 1.630 -158.545 1.800 ;
        RECT -155.575 1.800 -155.405 2.125 ;
        RECT -155.225 2.025 -154.855 2.365 ;
        RECT -154.675 2.125 -154.125 2.295 ;
        RECT -150.075 2.125 -149.525 2.295 ;
        RECT -154.675 1.800 -154.505 2.125 ;
        RECT -155.575 1.630 -154.505 1.800 ;
        RECT -149.695 1.800 -149.525 2.125 ;
        RECT -149.345 2.025 -148.975 2.365 ;
        RECT -148.795 2.125 -147.865 2.305 ;
        RECT -146.415 2.125 -145.485 2.305 ;
        RECT -148.795 1.800 -148.625 2.125 ;
        RECT -149.695 1.630 -148.625 1.800 ;
        RECT -145.655 1.800 -145.485 2.125 ;
        RECT -145.305 2.025 -144.935 2.365 ;
        RECT -144.755 2.125 -144.205 2.295 ;
        RECT -140.155 2.125 -139.605 2.295 ;
        RECT -144.755 1.800 -144.585 2.125 ;
        RECT -145.655 1.630 -144.585 1.800 ;
        RECT -139.775 1.800 -139.605 2.125 ;
        RECT -139.425 2.025 -139.055 2.365 ;
        RECT -138.875 2.125 -137.945 2.305 ;
        RECT -136.495 2.125 -135.565 2.305 ;
        RECT -138.875 1.800 -138.705 2.125 ;
        RECT -139.775 1.630 -138.705 1.800 ;
        RECT -135.735 1.800 -135.565 2.125 ;
        RECT -135.385 2.025 -135.015 2.365 ;
        RECT -134.835 2.125 -134.285 2.295 ;
        RECT -130.235 2.125 -129.685 2.295 ;
        RECT -134.835 1.800 -134.665 2.125 ;
        RECT -135.735 1.630 -134.665 1.800 ;
        RECT -129.855 1.800 -129.685 2.125 ;
        RECT -129.505 2.025 -129.135 2.365 ;
        RECT -128.955 2.125 -128.025 2.305 ;
        RECT -126.575 2.125 -125.645 2.305 ;
        RECT -128.955 1.800 -128.785 2.125 ;
        RECT -129.855 1.630 -128.785 1.800 ;
        RECT -125.815 1.800 -125.645 2.125 ;
        RECT -125.465 2.025 -125.095 2.365 ;
        RECT -124.915 2.125 -124.365 2.295 ;
        RECT -120.315 2.125 -119.765 2.295 ;
        RECT -124.915 1.800 -124.745 2.125 ;
        RECT -125.815 1.630 -124.745 1.800 ;
        RECT -119.935 1.800 -119.765 2.125 ;
        RECT -119.585 2.025 -119.215 2.365 ;
        RECT -119.035 2.125 -118.105 2.305 ;
        RECT -116.655 2.125 -115.725 2.305 ;
        RECT -119.035 1.800 -118.865 2.125 ;
        RECT -119.935 1.630 -118.865 1.800 ;
        RECT -115.895 1.800 -115.725 2.125 ;
        RECT -115.545 2.025 -115.175 2.365 ;
        RECT -114.995 2.125 -114.445 2.295 ;
        RECT -110.395 2.125 -109.845 2.295 ;
        RECT -114.995 1.800 -114.825 2.125 ;
        RECT -115.895 1.630 -114.825 1.800 ;
        RECT -110.015 1.800 -109.845 2.125 ;
        RECT -109.665 2.025 -109.295 2.365 ;
        RECT -109.115 2.125 -108.185 2.305 ;
        RECT -106.735 2.125 -105.805 2.305 ;
        RECT -109.115 1.800 -108.945 2.125 ;
        RECT -110.015 1.630 -108.945 1.800 ;
        RECT -105.975 1.800 -105.805 2.125 ;
        RECT -105.625 2.025 -105.255 2.365 ;
        RECT -105.075 2.125 -104.525 2.295 ;
        RECT -100.475 2.125 -99.925 2.295 ;
        RECT -105.075 1.800 -104.905 2.125 ;
        RECT -105.975 1.630 -104.905 1.800 ;
        RECT -100.095 1.800 -99.925 2.125 ;
        RECT -99.745 2.025 -99.375 2.365 ;
        RECT -99.195 2.125 -98.265 2.305 ;
        RECT -96.815 2.125 -95.885 2.305 ;
        RECT -99.195 1.800 -99.025 2.125 ;
        RECT -100.095 1.630 -99.025 1.800 ;
        RECT -96.055 1.800 -95.885 2.125 ;
        RECT -95.705 2.025 -95.335 2.365 ;
        RECT -95.155 2.125 -94.605 2.295 ;
        RECT -90.555 2.125 -90.005 2.295 ;
        RECT -95.155 1.800 -94.985 2.125 ;
        RECT -96.055 1.630 -94.985 1.800 ;
        RECT -90.175 1.800 -90.005 2.125 ;
        RECT -89.825 2.025 -89.455 2.365 ;
        RECT -89.275 2.125 -88.345 2.305 ;
        RECT -86.895 2.125 -85.965 2.305 ;
        RECT -89.275 1.800 -89.105 2.125 ;
        RECT -90.175 1.630 -89.105 1.800 ;
        RECT -86.135 1.800 -85.965 2.125 ;
        RECT -85.785 2.025 -85.415 2.365 ;
        RECT -85.235 2.125 -84.685 2.295 ;
        RECT -80.635 2.125 -80.085 2.295 ;
        RECT -85.235 1.800 -85.065 2.125 ;
        RECT -86.135 1.630 -85.065 1.800 ;
        RECT -80.255 1.800 -80.085 2.125 ;
        RECT -79.905 2.025 -79.535 2.365 ;
        RECT -79.355 2.125 -78.425 2.305 ;
        RECT -76.975 2.125 -76.045 2.305 ;
        RECT -79.355 1.800 -79.185 2.125 ;
        RECT -80.255 1.630 -79.185 1.800 ;
        RECT -76.215 1.800 -76.045 2.125 ;
        RECT -75.865 2.025 -75.495 2.365 ;
        RECT -75.315 2.125 -74.765 2.295 ;
        RECT -70.715 2.125 -70.165 2.295 ;
        RECT -75.315 1.800 -75.145 2.125 ;
        RECT -76.215 1.630 -75.145 1.800 ;
        RECT -70.335 1.800 -70.165 2.125 ;
        RECT -69.985 2.025 -69.615 2.365 ;
        RECT -69.435 2.125 -68.505 2.305 ;
        RECT -67.055 2.125 -66.125 2.305 ;
        RECT -69.435 1.800 -69.265 2.125 ;
        RECT -70.335 1.630 -69.265 1.800 ;
        RECT -66.295 1.800 -66.125 2.125 ;
        RECT -65.945 2.025 -65.575 2.365 ;
        RECT -65.395 2.125 -64.845 2.295 ;
        RECT -60.795 2.125 -60.245 2.295 ;
        RECT -65.395 1.800 -65.225 2.125 ;
        RECT -66.295 1.630 -65.225 1.800 ;
        RECT -60.415 1.800 -60.245 2.125 ;
        RECT -60.065 2.025 -59.695 2.365 ;
        RECT -59.515 2.125 -58.585 2.305 ;
        RECT -57.135 2.125 -56.205 2.305 ;
        RECT -59.515 1.800 -59.345 2.125 ;
        RECT -60.415 1.630 -59.345 1.800 ;
        RECT -56.375 1.800 -56.205 2.125 ;
        RECT -56.025 2.025 -55.655 2.365 ;
        RECT -55.475 2.125 -54.925 2.295 ;
        RECT -50.875 2.125 -50.325 2.295 ;
        RECT -55.475 1.800 -55.305 2.125 ;
        RECT -56.375 1.630 -55.305 1.800 ;
        RECT -50.495 1.800 -50.325 2.125 ;
        RECT -50.145 2.025 -49.775 2.365 ;
        RECT -49.595 2.125 -48.665 2.305 ;
        RECT -47.215 2.125 -46.285 2.305 ;
        RECT -49.595 1.800 -49.425 2.125 ;
        RECT -50.495 1.630 -49.425 1.800 ;
        RECT -46.455 1.800 -46.285 2.125 ;
        RECT -46.105 2.025 -45.735 2.365 ;
        RECT -45.555 2.125 -45.005 2.295 ;
        RECT -40.955 2.125 -40.405 2.295 ;
        RECT -45.555 1.800 -45.385 2.125 ;
        RECT -46.455 1.630 -45.385 1.800 ;
        RECT -40.575 1.800 -40.405 2.125 ;
        RECT -40.225 2.025 -39.855 2.365 ;
        RECT -39.675 2.125 -38.745 2.305 ;
        RECT -37.295 2.125 -36.365 2.305 ;
        RECT -39.675 1.800 -39.505 2.125 ;
        RECT -40.575 1.630 -39.505 1.800 ;
        RECT -36.535 1.800 -36.365 2.125 ;
        RECT -36.185 2.025 -35.815 2.365 ;
        RECT -35.635 2.125 -35.085 2.295 ;
        RECT -31.035 2.125 -30.485 2.295 ;
        RECT -35.635 1.800 -35.465 2.125 ;
        RECT -36.535 1.630 -35.465 1.800 ;
        RECT -30.655 1.800 -30.485 2.125 ;
        RECT -30.305 2.025 -29.935 2.365 ;
        RECT -29.755 2.125 -28.825 2.305 ;
        RECT -27.375 2.125 -26.445 2.305 ;
        RECT -29.755 1.800 -29.585 2.125 ;
        RECT -30.655 1.630 -29.585 1.800 ;
        RECT -26.615 1.800 -26.445 2.125 ;
        RECT -26.265 2.025 -25.895 2.365 ;
        RECT -25.715 2.125 -25.165 2.295 ;
        RECT -21.115 2.125 -20.565 2.295 ;
        RECT -25.715 1.800 -25.545 2.125 ;
        RECT -26.615 1.630 -25.545 1.800 ;
        RECT -20.735 1.800 -20.565 2.125 ;
        RECT -20.385 2.025 -20.015 2.365 ;
        RECT -19.835 2.125 -18.905 2.305 ;
        RECT -17.455 2.125 -16.525 2.305 ;
        RECT -19.835 1.800 -19.665 2.125 ;
        RECT -20.735 1.630 -19.665 1.800 ;
        RECT -16.695 1.800 -16.525 2.125 ;
        RECT -16.345 2.025 -15.975 2.365 ;
        RECT -15.795 2.125 -15.245 2.295 ;
        RECT -11.195 2.125 -10.645 2.295 ;
        RECT -15.795 1.800 -15.625 2.125 ;
        RECT -16.695 1.630 -15.625 1.800 ;
        RECT -10.815 1.800 -10.645 2.125 ;
        RECT -10.465 2.025 -10.095 2.365 ;
        RECT -9.915 2.125 -8.985 2.305 ;
        RECT -7.535 2.125 -6.605 2.305 ;
        RECT -9.915 1.800 -9.745 2.125 ;
        RECT -10.815 1.630 -9.745 1.800 ;
        RECT -6.775 1.800 -6.605 2.125 ;
        RECT -6.425 2.025 -6.055 2.365 ;
        RECT -5.875 2.125 -5.325 2.295 ;
        RECT -1.275 2.125 -0.725 2.295 ;
        RECT -5.875 1.800 -5.705 2.125 ;
        RECT -6.775 1.630 -5.705 1.800 ;
        RECT -0.895 1.800 -0.725 2.125 ;
        RECT -0.545 2.025 -0.175 2.365 ;
        RECT 0.005 2.125 0.935 2.305 ;
        RECT 2.385 2.125 3.315 2.305 ;
        RECT 0.005 1.800 0.175 2.125 ;
        RECT -0.895 1.630 0.175 1.800 ;
        RECT 3.145 1.800 3.315 2.125 ;
        RECT 3.495 2.025 3.865 2.365 ;
        RECT 4.045 2.125 4.595 2.295 ;
        RECT 8.645 2.125 9.195 2.295 ;
        RECT 4.045 1.800 4.215 2.125 ;
        RECT 3.145 1.630 4.215 1.800 ;
        RECT 9.025 1.800 9.195 2.125 ;
        RECT 9.375 2.025 9.745 2.365 ;
        RECT 9.925 2.125 10.855 2.305 ;
        RECT 12.305 2.125 13.235 2.305 ;
        RECT 9.925 1.800 10.095 2.125 ;
        RECT 9.025 1.630 10.095 1.800 ;
        RECT 13.065 1.800 13.235 2.125 ;
        RECT 13.415 2.025 13.785 2.365 ;
        RECT 13.965 2.125 14.515 2.295 ;
        RECT 18.565 2.125 19.115 2.295 ;
        RECT 13.965 1.800 14.135 2.125 ;
        RECT 13.065 1.630 14.135 1.800 ;
        RECT 18.945 1.800 19.115 2.125 ;
        RECT 19.295 2.025 19.665 2.365 ;
        RECT 19.845 2.125 20.775 2.305 ;
        RECT 22.225 2.125 23.155 2.305 ;
        RECT 19.845 1.800 20.015 2.125 ;
        RECT 18.945 1.630 20.015 1.800 ;
        RECT 22.985 1.800 23.155 2.125 ;
        RECT 23.335 2.025 23.705 2.365 ;
        RECT 23.885 2.125 24.435 2.295 ;
        RECT 23.885 1.800 24.055 2.125 ;
        RECT 24.605 1.945 24.775 2.470 ;
        RECT 22.985 1.630 24.055 1.800 ;
        RECT -289.295 1.430 -289.125 1.615 ;
        RECT -288.150 1.525 -287.820 1.630 ;
        RECT -284.220 1.525 -283.890 1.630 ;
        RECT -278.230 1.525 -277.900 1.630 ;
        RECT -274.300 1.525 -273.970 1.630 ;
        RECT -268.310 1.525 -267.980 1.630 ;
        RECT -264.380 1.525 -264.050 1.630 ;
        RECT -258.390 1.525 -258.060 1.630 ;
        RECT -254.460 1.525 -254.130 1.630 ;
        RECT -248.470 1.525 -248.140 1.630 ;
        RECT -244.540 1.525 -244.210 1.630 ;
        RECT -238.550 1.525 -238.220 1.630 ;
        RECT -234.620 1.525 -234.290 1.630 ;
        RECT -228.630 1.525 -228.300 1.630 ;
        RECT -224.700 1.525 -224.370 1.630 ;
        RECT -218.710 1.525 -218.380 1.630 ;
        RECT -214.780 1.525 -214.450 1.630 ;
        RECT -208.790 1.525 -208.460 1.630 ;
        RECT -204.860 1.525 -204.530 1.630 ;
        RECT -198.870 1.525 -198.540 1.630 ;
        RECT -194.940 1.525 -194.610 1.630 ;
        RECT -188.950 1.525 -188.620 1.630 ;
        RECT -185.020 1.525 -184.690 1.630 ;
        RECT -179.030 1.525 -178.700 1.630 ;
        RECT -175.100 1.525 -174.770 1.630 ;
        RECT -169.110 1.525 -168.780 1.630 ;
        RECT -165.180 1.525 -164.850 1.630 ;
        RECT -159.190 1.525 -158.860 1.630 ;
        RECT -155.260 1.525 -154.930 1.630 ;
        RECT -149.270 1.525 -148.940 1.630 ;
        RECT -145.340 1.525 -145.010 1.630 ;
        RECT -139.350 1.525 -139.020 1.630 ;
        RECT -135.420 1.525 -135.090 1.630 ;
        RECT -129.430 1.525 -129.100 1.630 ;
        RECT -125.500 1.525 -125.170 1.630 ;
        RECT -119.510 1.525 -119.180 1.630 ;
        RECT -115.580 1.525 -115.250 1.630 ;
        RECT -109.590 1.525 -109.260 1.630 ;
        RECT -105.660 1.525 -105.330 1.630 ;
        RECT -99.670 1.525 -99.340 1.630 ;
        RECT -95.740 1.525 -95.410 1.630 ;
        RECT -89.750 1.525 -89.420 1.630 ;
        RECT -85.820 1.525 -85.490 1.630 ;
        RECT -79.830 1.525 -79.500 1.630 ;
        RECT -75.900 1.525 -75.570 1.630 ;
        RECT -69.910 1.525 -69.580 1.630 ;
        RECT -65.980 1.525 -65.650 1.630 ;
        RECT -59.990 1.525 -59.660 1.630 ;
        RECT -56.060 1.525 -55.730 1.630 ;
        RECT -50.070 1.525 -49.740 1.630 ;
        RECT -46.140 1.525 -45.810 1.630 ;
        RECT -40.150 1.525 -39.820 1.630 ;
        RECT -36.220 1.525 -35.890 1.630 ;
        RECT -30.230 1.525 -29.900 1.630 ;
        RECT -26.300 1.525 -25.970 1.630 ;
        RECT -20.310 1.525 -19.980 1.630 ;
        RECT -16.380 1.525 -16.050 1.630 ;
        RECT -10.390 1.525 -10.060 1.630 ;
        RECT -6.460 1.525 -6.130 1.630 ;
        RECT -0.470 1.525 -0.140 1.630 ;
        RECT 3.460 1.525 3.790 1.630 ;
        RECT 9.450 1.525 9.780 1.630 ;
        RECT 13.380 1.525 13.710 1.630 ;
        RECT 19.370 1.525 19.700 1.630 ;
        RECT 23.300 1.525 23.630 1.630 ;
        RECT 24.225 1.615 24.775 1.945 ;
        RECT -289.825 1.415 -289.125 1.430 ;
        RECT -289.910 1.245 -289.125 1.415 ;
        RECT -289.590 1.240 -289.125 1.245 ;
        RECT -289.295 1.090 -289.125 1.240 ;
        RECT -285.295 1.355 -284.390 1.445 ;
        RECT -283.590 1.355 -283.085 1.435 ;
        RECT -285.295 1.175 -283.085 1.355 ;
        RECT -275.375 1.355 -274.470 1.445 ;
        RECT -273.670 1.355 -273.165 1.435 ;
        RECT -275.375 1.175 -273.165 1.355 ;
        RECT -265.455 1.355 -264.550 1.445 ;
        RECT -263.750 1.355 -263.245 1.435 ;
        RECT -265.455 1.175 -263.245 1.355 ;
        RECT -255.535 1.355 -254.630 1.445 ;
        RECT -253.830 1.355 -253.325 1.435 ;
        RECT -255.535 1.175 -253.325 1.355 ;
        RECT -245.615 1.355 -244.710 1.445 ;
        RECT -243.910 1.355 -243.405 1.435 ;
        RECT -245.615 1.175 -243.405 1.355 ;
        RECT -235.695 1.355 -234.790 1.445 ;
        RECT -233.990 1.355 -233.485 1.435 ;
        RECT -235.695 1.175 -233.485 1.355 ;
        RECT -225.775 1.355 -224.870 1.445 ;
        RECT -224.070 1.355 -223.565 1.435 ;
        RECT -225.775 1.175 -223.565 1.355 ;
        RECT -215.855 1.355 -214.950 1.445 ;
        RECT -214.150 1.355 -213.645 1.435 ;
        RECT -215.855 1.175 -213.645 1.355 ;
        RECT -205.935 1.355 -205.030 1.445 ;
        RECT -204.230 1.355 -203.725 1.435 ;
        RECT -205.935 1.175 -203.725 1.355 ;
        RECT -196.015 1.355 -195.110 1.445 ;
        RECT -194.310 1.355 -193.805 1.435 ;
        RECT -196.015 1.175 -193.805 1.355 ;
        RECT -186.095 1.355 -185.190 1.445 ;
        RECT -184.390 1.355 -183.885 1.435 ;
        RECT -186.095 1.175 -183.885 1.355 ;
        RECT -176.175 1.355 -175.270 1.445 ;
        RECT -174.470 1.355 -173.965 1.435 ;
        RECT -176.175 1.175 -173.965 1.355 ;
        RECT -166.255 1.355 -165.350 1.445 ;
        RECT -164.550 1.355 -164.045 1.435 ;
        RECT -166.255 1.175 -164.045 1.355 ;
        RECT -156.335 1.355 -155.430 1.445 ;
        RECT -154.630 1.355 -154.125 1.435 ;
        RECT -156.335 1.175 -154.125 1.355 ;
        RECT -146.415 1.355 -145.510 1.445 ;
        RECT -144.710 1.355 -144.205 1.435 ;
        RECT -146.415 1.175 -144.205 1.355 ;
        RECT -136.495 1.355 -135.590 1.445 ;
        RECT -134.790 1.355 -134.285 1.435 ;
        RECT -136.495 1.175 -134.285 1.355 ;
        RECT -126.575 1.355 -125.670 1.445 ;
        RECT -124.870 1.355 -124.365 1.435 ;
        RECT -126.575 1.175 -124.365 1.355 ;
        RECT -116.655 1.355 -115.750 1.445 ;
        RECT -114.950 1.355 -114.445 1.435 ;
        RECT -116.655 1.175 -114.445 1.355 ;
        RECT -106.735 1.355 -105.830 1.445 ;
        RECT -105.030 1.355 -104.525 1.435 ;
        RECT -106.735 1.175 -104.525 1.355 ;
        RECT -96.815 1.355 -95.910 1.445 ;
        RECT -95.110 1.355 -94.605 1.435 ;
        RECT -96.815 1.175 -94.605 1.355 ;
        RECT -86.895 1.355 -85.990 1.445 ;
        RECT -85.190 1.355 -84.685 1.435 ;
        RECT -86.895 1.175 -84.685 1.355 ;
        RECT -76.975 1.355 -76.070 1.445 ;
        RECT -75.270 1.355 -74.765 1.435 ;
        RECT -76.975 1.175 -74.765 1.355 ;
        RECT -67.055 1.355 -66.150 1.445 ;
        RECT -65.350 1.355 -64.845 1.435 ;
        RECT -67.055 1.175 -64.845 1.355 ;
        RECT -57.135 1.355 -56.230 1.445 ;
        RECT -55.430 1.355 -54.925 1.435 ;
        RECT -57.135 1.175 -54.925 1.355 ;
        RECT -47.215 1.355 -46.310 1.445 ;
        RECT -45.510 1.355 -45.005 1.435 ;
        RECT -47.215 1.175 -45.005 1.355 ;
        RECT -37.295 1.355 -36.390 1.445 ;
        RECT -35.590 1.355 -35.085 1.435 ;
        RECT -37.295 1.175 -35.085 1.355 ;
        RECT -27.375 1.355 -26.470 1.445 ;
        RECT -25.670 1.355 -25.165 1.435 ;
        RECT -27.375 1.175 -25.165 1.355 ;
        RECT -17.455 1.355 -16.550 1.445 ;
        RECT -15.750 1.355 -15.245 1.435 ;
        RECT -17.455 1.175 -15.245 1.355 ;
        RECT -7.535 1.355 -6.630 1.445 ;
        RECT -5.830 1.355 -5.325 1.435 ;
        RECT -7.535 1.175 -5.325 1.355 ;
        RECT 2.385 1.355 3.290 1.445 ;
        RECT 4.090 1.355 4.595 1.435 ;
        RECT 2.385 1.175 4.595 1.355 ;
        RECT 12.305 1.355 13.210 1.445 ;
        RECT 14.010 1.355 14.515 1.435 ;
        RECT 12.305 1.175 14.515 1.355 ;
        RECT 22.225 1.355 23.130 1.445 ;
        RECT 23.930 1.355 24.435 1.435 ;
        RECT 22.225 1.175 24.435 1.355 ;
        RECT 24.605 1.420 24.775 1.615 ;
        RECT 25.015 1.420 25.305 2.140 ;
        RECT 24.605 1.415 25.305 1.420 ;
        RECT 24.605 1.245 25.390 1.415 ;
        RECT 24.605 1.240 25.070 1.245 ;
        RECT 24.605 1.090 24.775 1.240 ;
        RECT -288.835 -86.070 -288.665 -85.920 ;
        RECT -289.450 -86.240 -288.665 -86.070 ;
        RECT -289.365 -87.405 -289.075 -86.240 ;
        RECT -288.835 -86.445 -288.665 -86.240 ;
        RECT -288.495 -86.185 -286.285 -86.005 ;
        RECT -288.495 -86.275 -287.590 -86.185 ;
        RECT -286.790 -86.265 -286.285 -86.185 ;
        RECT -278.575 -86.185 -276.365 -86.005 ;
        RECT -278.575 -86.275 -277.670 -86.185 ;
        RECT -276.870 -86.265 -276.365 -86.185 ;
        RECT -268.655 -86.185 -266.445 -86.005 ;
        RECT -268.655 -86.275 -267.750 -86.185 ;
        RECT -266.950 -86.265 -266.445 -86.185 ;
        RECT -258.735 -86.185 -256.525 -86.005 ;
        RECT -258.735 -86.275 -257.830 -86.185 ;
        RECT -257.030 -86.265 -256.525 -86.185 ;
        RECT -248.815 -86.185 -246.605 -86.005 ;
        RECT -248.815 -86.275 -247.910 -86.185 ;
        RECT -247.110 -86.265 -246.605 -86.185 ;
        RECT -238.895 -86.185 -236.685 -86.005 ;
        RECT -238.895 -86.275 -237.990 -86.185 ;
        RECT -237.190 -86.265 -236.685 -86.185 ;
        RECT -228.975 -86.185 -226.765 -86.005 ;
        RECT -228.975 -86.275 -228.070 -86.185 ;
        RECT -227.270 -86.265 -226.765 -86.185 ;
        RECT -219.055 -86.185 -216.845 -86.005 ;
        RECT -219.055 -86.275 -218.150 -86.185 ;
        RECT -217.350 -86.265 -216.845 -86.185 ;
        RECT -209.135 -86.185 -206.925 -86.005 ;
        RECT -209.135 -86.275 -208.230 -86.185 ;
        RECT -207.430 -86.265 -206.925 -86.185 ;
        RECT -199.215 -86.185 -197.005 -86.005 ;
        RECT -199.215 -86.275 -198.310 -86.185 ;
        RECT -197.510 -86.265 -197.005 -86.185 ;
        RECT -189.295 -86.185 -187.085 -86.005 ;
        RECT -189.295 -86.275 -188.390 -86.185 ;
        RECT -187.590 -86.265 -187.085 -86.185 ;
        RECT -179.375 -86.185 -177.165 -86.005 ;
        RECT -179.375 -86.275 -178.470 -86.185 ;
        RECT -177.670 -86.265 -177.165 -86.185 ;
        RECT -169.455 -86.185 -167.245 -86.005 ;
        RECT -169.455 -86.275 -168.550 -86.185 ;
        RECT -167.750 -86.265 -167.245 -86.185 ;
        RECT -159.535 -86.185 -157.325 -86.005 ;
        RECT -159.535 -86.275 -158.630 -86.185 ;
        RECT -157.830 -86.265 -157.325 -86.185 ;
        RECT -149.615 -86.185 -147.405 -86.005 ;
        RECT -149.615 -86.275 -148.710 -86.185 ;
        RECT -147.910 -86.265 -147.405 -86.185 ;
        RECT -139.695 -86.185 -137.485 -86.005 ;
        RECT -139.695 -86.275 -138.790 -86.185 ;
        RECT -137.990 -86.265 -137.485 -86.185 ;
        RECT -129.775 -86.185 -127.565 -86.005 ;
        RECT -129.775 -86.275 -128.870 -86.185 ;
        RECT -128.070 -86.265 -127.565 -86.185 ;
        RECT -119.855 -86.185 -117.645 -86.005 ;
        RECT -119.855 -86.275 -118.950 -86.185 ;
        RECT -118.150 -86.265 -117.645 -86.185 ;
        RECT -109.935 -86.185 -107.725 -86.005 ;
        RECT -109.935 -86.275 -109.030 -86.185 ;
        RECT -108.230 -86.265 -107.725 -86.185 ;
        RECT -100.015 -86.185 -97.805 -86.005 ;
        RECT -100.015 -86.275 -99.110 -86.185 ;
        RECT -98.310 -86.265 -97.805 -86.185 ;
        RECT -90.095 -86.185 -87.885 -86.005 ;
        RECT -90.095 -86.275 -89.190 -86.185 ;
        RECT -88.390 -86.265 -87.885 -86.185 ;
        RECT -80.175 -86.185 -77.965 -86.005 ;
        RECT -80.175 -86.275 -79.270 -86.185 ;
        RECT -78.470 -86.265 -77.965 -86.185 ;
        RECT -70.255 -86.185 -68.045 -86.005 ;
        RECT -70.255 -86.275 -69.350 -86.185 ;
        RECT -68.550 -86.265 -68.045 -86.185 ;
        RECT -60.335 -86.185 -58.125 -86.005 ;
        RECT -60.335 -86.275 -59.430 -86.185 ;
        RECT -58.630 -86.265 -58.125 -86.185 ;
        RECT -50.415 -86.185 -48.205 -86.005 ;
        RECT -50.415 -86.275 -49.510 -86.185 ;
        RECT -48.710 -86.265 -48.205 -86.185 ;
        RECT -40.495 -86.185 -38.285 -86.005 ;
        RECT -40.495 -86.275 -39.590 -86.185 ;
        RECT -38.790 -86.265 -38.285 -86.185 ;
        RECT -30.575 -86.185 -28.365 -86.005 ;
        RECT -30.575 -86.275 -29.670 -86.185 ;
        RECT -28.870 -86.265 -28.365 -86.185 ;
        RECT -20.655 -86.185 -18.445 -86.005 ;
        RECT -20.655 -86.275 -19.750 -86.185 ;
        RECT -18.950 -86.265 -18.445 -86.185 ;
        RECT -10.735 -86.185 -8.525 -86.005 ;
        RECT -10.735 -86.275 -9.830 -86.185 ;
        RECT -9.030 -86.265 -8.525 -86.185 ;
        RECT -0.815 -86.185 1.395 -86.005 ;
        RECT -0.815 -86.275 0.090 -86.185 ;
        RECT 0.890 -86.265 1.395 -86.185 ;
        RECT 9.105 -86.185 11.315 -86.005 ;
        RECT 9.105 -86.275 10.010 -86.185 ;
        RECT 10.810 -86.265 11.315 -86.185 ;
        RECT 19.025 -86.185 21.235 -86.005 ;
        RECT 19.025 -86.275 19.930 -86.185 ;
        RECT 20.730 -86.265 21.235 -86.185 ;
        RECT -288.835 -86.775 -287.905 -86.445 ;
        RECT -287.420 -86.460 -287.090 -86.355 ;
        RECT -281.430 -86.460 -281.100 -86.355 ;
        RECT -277.500 -86.460 -277.170 -86.355 ;
        RECT -271.510 -86.460 -271.180 -86.355 ;
        RECT -267.580 -86.460 -267.250 -86.355 ;
        RECT -261.590 -86.460 -261.260 -86.355 ;
        RECT -257.660 -86.460 -257.330 -86.355 ;
        RECT -251.670 -86.460 -251.340 -86.355 ;
        RECT -247.740 -86.460 -247.410 -86.355 ;
        RECT -241.750 -86.460 -241.420 -86.355 ;
        RECT -237.820 -86.460 -237.490 -86.355 ;
        RECT -231.830 -86.460 -231.500 -86.355 ;
        RECT -227.900 -86.460 -227.570 -86.355 ;
        RECT -221.910 -86.460 -221.580 -86.355 ;
        RECT -217.980 -86.460 -217.650 -86.355 ;
        RECT -211.990 -86.460 -211.660 -86.355 ;
        RECT -208.060 -86.460 -207.730 -86.355 ;
        RECT -202.070 -86.460 -201.740 -86.355 ;
        RECT -198.140 -86.460 -197.810 -86.355 ;
        RECT -192.150 -86.460 -191.820 -86.355 ;
        RECT -188.220 -86.460 -187.890 -86.355 ;
        RECT -182.230 -86.460 -181.900 -86.355 ;
        RECT -178.300 -86.460 -177.970 -86.355 ;
        RECT -172.310 -86.460 -171.980 -86.355 ;
        RECT -168.380 -86.460 -168.050 -86.355 ;
        RECT -162.390 -86.460 -162.060 -86.355 ;
        RECT -158.460 -86.460 -158.130 -86.355 ;
        RECT -152.470 -86.460 -152.140 -86.355 ;
        RECT -148.540 -86.460 -148.210 -86.355 ;
        RECT -142.550 -86.460 -142.220 -86.355 ;
        RECT -138.620 -86.460 -138.290 -86.355 ;
        RECT -132.630 -86.460 -132.300 -86.355 ;
        RECT -128.700 -86.460 -128.370 -86.355 ;
        RECT -122.710 -86.460 -122.380 -86.355 ;
        RECT -118.780 -86.460 -118.450 -86.355 ;
        RECT -112.790 -86.460 -112.460 -86.355 ;
        RECT -108.860 -86.460 -108.530 -86.355 ;
        RECT -102.870 -86.460 -102.540 -86.355 ;
        RECT -98.940 -86.460 -98.610 -86.355 ;
        RECT -92.950 -86.460 -92.620 -86.355 ;
        RECT -89.020 -86.460 -88.690 -86.355 ;
        RECT -83.030 -86.460 -82.700 -86.355 ;
        RECT -79.100 -86.460 -78.770 -86.355 ;
        RECT -73.110 -86.460 -72.780 -86.355 ;
        RECT -69.180 -86.460 -68.850 -86.355 ;
        RECT -63.190 -86.460 -62.860 -86.355 ;
        RECT -59.260 -86.460 -58.930 -86.355 ;
        RECT -53.270 -86.460 -52.940 -86.355 ;
        RECT -49.340 -86.460 -49.010 -86.355 ;
        RECT -43.350 -86.460 -43.020 -86.355 ;
        RECT -39.420 -86.460 -39.090 -86.355 ;
        RECT -33.430 -86.460 -33.100 -86.355 ;
        RECT -29.500 -86.460 -29.170 -86.355 ;
        RECT -23.510 -86.460 -23.180 -86.355 ;
        RECT -19.580 -86.460 -19.250 -86.355 ;
        RECT -13.590 -86.460 -13.260 -86.355 ;
        RECT -9.660 -86.460 -9.330 -86.355 ;
        RECT -3.670 -86.460 -3.340 -86.355 ;
        RECT 0.260 -86.460 0.590 -86.355 ;
        RECT 6.250 -86.460 6.580 -86.355 ;
        RECT 10.180 -86.460 10.510 -86.355 ;
        RECT 16.170 -86.460 16.500 -86.355 ;
        RECT 20.100 -86.460 20.430 -86.355 ;
        RECT 26.090 -86.460 26.420 -86.355 ;
        RECT -287.735 -86.630 -286.665 -86.460 ;
        RECT -288.835 -87.300 -288.665 -86.775 ;
        RECT -287.735 -86.955 -287.565 -86.630 ;
        RECT -288.495 -87.135 -287.565 -86.955 ;
        RECT -287.385 -87.195 -287.015 -86.855 ;
        RECT -286.835 -86.955 -286.665 -86.630 ;
        RECT -281.855 -86.630 -280.785 -86.460 ;
        RECT -281.855 -86.955 -281.685 -86.630 ;
        RECT -286.835 -87.125 -286.285 -86.955 ;
        RECT -282.235 -87.125 -281.685 -86.955 ;
        RECT -281.505 -87.195 -281.135 -86.855 ;
        RECT -280.955 -86.955 -280.785 -86.630 ;
        RECT -277.815 -86.630 -276.745 -86.460 ;
        RECT -277.815 -86.955 -277.645 -86.630 ;
        RECT -280.955 -87.135 -280.025 -86.955 ;
        RECT -278.575 -87.135 -277.645 -86.955 ;
        RECT -277.465 -87.195 -277.095 -86.855 ;
        RECT -276.915 -86.955 -276.745 -86.630 ;
        RECT -271.935 -86.630 -270.865 -86.460 ;
        RECT -271.935 -86.955 -271.765 -86.630 ;
        RECT -276.915 -87.125 -276.365 -86.955 ;
        RECT -272.315 -87.125 -271.765 -86.955 ;
        RECT -271.585 -87.195 -271.215 -86.855 ;
        RECT -271.035 -86.955 -270.865 -86.630 ;
        RECT -267.895 -86.630 -266.825 -86.460 ;
        RECT -267.895 -86.955 -267.725 -86.630 ;
        RECT -271.035 -87.135 -270.105 -86.955 ;
        RECT -268.655 -87.135 -267.725 -86.955 ;
        RECT -267.545 -87.195 -267.175 -86.855 ;
        RECT -266.995 -86.955 -266.825 -86.630 ;
        RECT -262.015 -86.630 -260.945 -86.460 ;
        RECT -262.015 -86.955 -261.845 -86.630 ;
        RECT -266.995 -87.125 -266.445 -86.955 ;
        RECT -262.395 -87.125 -261.845 -86.955 ;
        RECT -261.665 -87.195 -261.295 -86.855 ;
        RECT -261.115 -86.955 -260.945 -86.630 ;
        RECT -257.975 -86.630 -256.905 -86.460 ;
        RECT -257.975 -86.955 -257.805 -86.630 ;
        RECT -261.115 -87.135 -260.185 -86.955 ;
        RECT -258.735 -87.135 -257.805 -86.955 ;
        RECT -257.625 -87.195 -257.255 -86.855 ;
        RECT -257.075 -86.955 -256.905 -86.630 ;
        RECT -252.095 -86.630 -251.025 -86.460 ;
        RECT -252.095 -86.955 -251.925 -86.630 ;
        RECT -257.075 -87.125 -256.525 -86.955 ;
        RECT -252.475 -87.125 -251.925 -86.955 ;
        RECT -251.745 -87.195 -251.375 -86.855 ;
        RECT -251.195 -86.955 -251.025 -86.630 ;
        RECT -248.055 -86.630 -246.985 -86.460 ;
        RECT -248.055 -86.955 -247.885 -86.630 ;
        RECT -251.195 -87.135 -250.265 -86.955 ;
        RECT -248.815 -87.135 -247.885 -86.955 ;
        RECT -247.705 -87.195 -247.335 -86.855 ;
        RECT -247.155 -86.955 -246.985 -86.630 ;
        RECT -242.175 -86.630 -241.105 -86.460 ;
        RECT -242.175 -86.955 -242.005 -86.630 ;
        RECT -247.155 -87.125 -246.605 -86.955 ;
        RECT -242.555 -87.125 -242.005 -86.955 ;
        RECT -241.825 -87.195 -241.455 -86.855 ;
        RECT -241.275 -86.955 -241.105 -86.630 ;
        RECT -238.135 -86.630 -237.065 -86.460 ;
        RECT -238.135 -86.955 -237.965 -86.630 ;
        RECT -241.275 -87.135 -240.345 -86.955 ;
        RECT -238.895 -87.135 -237.965 -86.955 ;
        RECT -237.785 -87.195 -237.415 -86.855 ;
        RECT -237.235 -86.955 -237.065 -86.630 ;
        RECT -232.255 -86.630 -231.185 -86.460 ;
        RECT -232.255 -86.955 -232.085 -86.630 ;
        RECT -237.235 -87.125 -236.685 -86.955 ;
        RECT -232.635 -87.125 -232.085 -86.955 ;
        RECT -231.905 -87.195 -231.535 -86.855 ;
        RECT -231.355 -86.955 -231.185 -86.630 ;
        RECT -228.215 -86.630 -227.145 -86.460 ;
        RECT -228.215 -86.955 -228.045 -86.630 ;
        RECT -231.355 -87.135 -230.425 -86.955 ;
        RECT -228.975 -87.135 -228.045 -86.955 ;
        RECT -227.865 -87.195 -227.495 -86.855 ;
        RECT -227.315 -86.955 -227.145 -86.630 ;
        RECT -222.335 -86.630 -221.265 -86.460 ;
        RECT -222.335 -86.955 -222.165 -86.630 ;
        RECT -227.315 -87.125 -226.765 -86.955 ;
        RECT -222.715 -87.125 -222.165 -86.955 ;
        RECT -221.985 -87.195 -221.615 -86.855 ;
        RECT -221.435 -86.955 -221.265 -86.630 ;
        RECT -218.295 -86.630 -217.225 -86.460 ;
        RECT -218.295 -86.955 -218.125 -86.630 ;
        RECT -221.435 -87.135 -220.505 -86.955 ;
        RECT -219.055 -87.135 -218.125 -86.955 ;
        RECT -217.945 -87.195 -217.575 -86.855 ;
        RECT -217.395 -86.955 -217.225 -86.630 ;
        RECT -212.415 -86.630 -211.345 -86.460 ;
        RECT -212.415 -86.955 -212.245 -86.630 ;
        RECT -217.395 -87.125 -216.845 -86.955 ;
        RECT -212.795 -87.125 -212.245 -86.955 ;
        RECT -212.065 -87.195 -211.695 -86.855 ;
        RECT -211.515 -86.955 -211.345 -86.630 ;
        RECT -208.375 -86.630 -207.305 -86.460 ;
        RECT -208.375 -86.955 -208.205 -86.630 ;
        RECT -211.515 -87.135 -210.585 -86.955 ;
        RECT -209.135 -87.135 -208.205 -86.955 ;
        RECT -208.025 -87.195 -207.655 -86.855 ;
        RECT -207.475 -86.955 -207.305 -86.630 ;
        RECT -202.495 -86.630 -201.425 -86.460 ;
        RECT -202.495 -86.955 -202.325 -86.630 ;
        RECT -207.475 -87.125 -206.925 -86.955 ;
        RECT -202.875 -87.125 -202.325 -86.955 ;
        RECT -202.145 -87.195 -201.775 -86.855 ;
        RECT -201.595 -86.955 -201.425 -86.630 ;
        RECT -198.455 -86.630 -197.385 -86.460 ;
        RECT -198.455 -86.955 -198.285 -86.630 ;
        RECT -201.595 -87.135 -200.665 -86.955 ;
        RECT -199.215 -87.135 -198.285 -86.955 ;
        RECT -198.105 -87.195 -197.735 -86.855 ;
        RECT -197.555 -86.955 -197.385 -86.630 ;
        RECT -192.575 -86.630 -191.505 -86.460 ;
        RECT -192.575 -86.955 -192.405 -86.630 ;
        RECT -197.555 -87.125 -197.005 -86.955 ;
        RECT -192.955 -87.125 -192.405 -86.955 ;
        RECT -192.225 -87.195 -191.855 -86.855 ;
        RECT -191.675 -86.955 -191.505 -86.630 ;
        RECT -188.535 -86.630 -187.465 -86.460 ;
        RECT -188.535 -86.955 -188.365 -86.630 ;
        RECT -191.675 -87.135 -190.745 -86.955 ;
        RECT -189.295 -87.135 -188.365 -86.955 ;
        RECT -188.185 -87.195 -187.815 -86.855 ;
        RECT -187.635 -86.955 -187.465 -86.630 ;
        RECT -182.655 -86.630 -181.585 -86.460 ;
        RECT -182.655 -86.955 -182.485 -86.630 ;
        RECT -187.635 -87.125 -187.085 -86.955 ;
        RECT -183.035 -87.125 -182.485 -86.955 ;
        RECT -182.305 -87.195 -181.935 -86.855 ;
        RECT -181.755 -86.955 -181.585 -86.630 ;
        RECT -178.615 -86.630 -177.545 -86.460 ;
        RECT -178.615 -86.955 -178.445 -86.630 ;
        RECT -181.755 -87.135 -180.825 -86.955 ;
        RECT -179.375 -87.135 -178.445 -86.955 ;
        RECT -178.265 -87.195 -177.895 -86.855 ;
        RECT -177.715 -86.955 -177.545 -86.630 ;
        RECT -172.735 -86.630 -171.665 -86.460 ;
        RECT -172.735 -86.955 -172.565 -86.630 ;
        RECT -177.715 -87.125 -177.165 -86.955 ;
        RECT -173.115 -87.125 -172.565 -86.955 ;
        RECT -172.385 -87.195 -172.015 -86.855 ;
        RECT -171.835 -86.955 -171.665 -86.630 ;
        RECT -168.695 -86.630 -167.625 -86.460 ;
        RECT -168.695 -86.955 -168.525 -86.630 ;
        RECT -171.835 -87.135 -170.905 -86.955 ;
        RECT -169.455 -87.135 -168.525 -86.955 ;
        RECT -168.345 -87.195 -167.975 -86.855 ;
        RECT -167.795 -86.955 -167.625 -86.630 ;
        RECT -162.815 -86.630 -161.745 -86.460 ;
        RECT -162.815 -86.955 -162.645 -86.630 ;
        RECT -167.795 -87.125 -167.245 -86.955 ;
        RECT -163.195 -87.125 -162.645 -86.955 ;
        RECT -162.465 -87.195 -162.095 -86.855 ;
        RECT -161.915 -86.955 -161.745 -86.630 ;
        RECT -158.775 -86.630 -157.705 -86.460 ;
        RECT -158.775 -86.955 -158.605 -86.630 ;
        RECT -161.915 -87.135 -160.985 -86.955 ;
        RECT -159.535 -87.135 -158.605 -86.955 ;
        RECT -158.425 -87.195 -158.055 -86.855 ;
        RECT -157.875 -86.955 -157.705 -86.630 ;
        RECT -152.895 -86.630 -151.825 -86.460 ;
        RECT -152.895 -86.955 -152.725 -86.630 ;
        RECT -157.875 -87.125 -157.325 -86.955 ;
        RECT -153.275 -87.125 -152.725 -86.955 ;
        RECT -152.545 -87.195 -152.175 -86.855 ;
        RECT -151.995 -86.955 -151.825 -86.630 ;
        RECT -148.855 -86.630 -147.785 -86.460 ;
        RECT -148.855 -86.955 -148.685 -86.630 ;
        RECT -151.995 -87.135 -151.065 -86.955 ;
        RECT -149.615 -87.135 -148.685 -86.955 ;
        RECT -148.505 -87.195 -148.135 -86.855 ;
        RECT -147.955 -86.955 -147.785 -86.630 ;
        RECT -142.975 -86.630 -141.905 -86.460 ;
        RECT -142.975 -86.955 -142.805 -86.630 ;
        RECT -147.955 -87.125 -147.405 -86.955 ;
        RECT -143.355 -87.125 -142.805 -86.955 ;
        RECT -142.625 -87.195 -142.255 -86.855 ;
        RECT -142.075 -86.955 -141.905 -86.630 ;
        RECT -138.935 -86.630 -137.865 -86.460 ;
        RECT -138.935 -86.955 -138.765 -86.630 ;
        RECT -142.075 -87.135 -141.145 -86.955 ;
        RECT -139.695 -87.135 -138.765 -86.955 ;
        RECT -138.585 -87.195 -138.215 -86.855 ;
        RECT -138.035 -86.955 -137.865 -86.630 ;
        RECT -133.055 -86.630 -131.985 -86.460 ;
        RECT -133.055 -86.955 -132.885 -86.630 ;
        RECT -138.035 -87.125 -137.485 -86.955 ;
        RECT -133.435 -87.125 -132.885 -86.955 ;
        RECT -132.705 -87.195 -132.335 -86.855 ;
        RECT -132.155 -86.955 -131.985 -86.630 ;
        RECT -129.015 -86.630 -127.945 -86.460 ;
        RECT -129.015 -86.955 -128.845 -86.630 ;
        RECT -132.155 -87.135 -131.225 -86.955 ;
        RECT -129.775 -87.135 -128.845 -86.955 ;
        RECT -128.665 -87.195 -128.295 -86.855 ;
        RECT -128.115 -86.955 -127.945 -86.630 ;
        RECT -123.135 -86.630 -122.065 -86.460 ;
        RECT -123.135 -86.955 -122.965 -86.630 ;
        RECT -128.115 -87.125 -127.565 -86.955 ;
        RECT -123.515 -87.125 -122.965 -86.955 ;
        RECT -122.785 -87.195 -122.415 -86.855 ;
        RECT -122.235 -86.955 -122.065 -86.630 ;
        RECT -119.095 -86.630 -118.025 -86.460 ;
        RECT -119.095 -86.955 -118.925 -86.630 ;
        RECT -122.235 -87.135 -121.305 -86.955 ;
        RECT -119.855 -87.135 -118.925 -86.955 ;
        RECT -118.745 -87.195 -118.375 -86.855 ;
        RECT -118.195 -86.955 -118.025 -86.630 ;
        RECT -113.215 -86.630 -112.145 -86.460 ;
        RECT -113.215 -86.955 -113.045 -86.630 ;
        RECT -118.195 -87.125 -117.645 -86.955 ;
        RECT -113.595 -87.125 -113.045 -86.955 ;
        RECT -112.865 -87.195 -112.495 -86.855 ;
        RECT -112.315 -86.955 -112.145 -86.630 ;
        RECT -109.175 -86.630 -108.105 -86.460 ;
        RECT -109.175 -86.955 -109.005 -86.630 ;
        RECT -112.315 -87.135 -111.385 -86.955 ;
        RECT -109.935 -87.135 -109.005 -86.955 ;
        RECT -108.825 -87.195 -108.455 -86.855 ;
        RECT -108.275 -86.955 -108.105 -86.630 ;
        RECT -103.295 -86.630 -102.225 -86.460 ;
        RECT -103.295 -86.955 -103.125 -86.630 ;
        RECT -108.275 -87.125 -107.725 -86.955 ;
        RECT -103.675 -87.125 -103.125 -86.955 ;
        RECT -102.945 -87.195 -102.575 -86.855 ;
        RECT -102.395 -86.955 -102.225 -86.630 ;
        RECT -99.255 -86.630 -98.185 -86.460 ;
        RECT -99.255 -86.955 -99.085 -86.630 ;
        RECT -102.395 -87.135 -101.465 -86.955 ;
        RECT -100.015 -87.135 -99.085 -86.955 ;
        RECT -98.905 -87.195 -98.535 -86.855 ;
        RECT -98.355 -86.955 -98.185 -86.630 ;
        RECT -93.375 -86.630 -92.305 -86.460 ;
        RECT -93.375 -86.955 -93.205 -86.630 ;
        RECT -98.355 -87.125 -97.805 -86.955 ;
        RECT -93.755 -87.125 -93.205 -86.955 ;
        RECT -93.025 -87.195 -92.655 -86.855 ;
        RECT -92.475 -86.955 -92.305 -86.630 ;
        RECT -89.335 -86.630 -88.265 -86.460 ;
        RECT -89.335 -86.955 -89.165 -86.630 ;
        RECT -92.475 -87.135 -91.545 -86.955 ;
        RECT -90.095 -87.135 -89.165 -86.955 ;
        RECT -88.985 -87.195 -88.615 -86.855 ;
        RECT -88.435 -86.955 -88.265 -86.630 ;
        RECT -83.455 -86.630 -82.385 -86.460 ;
        RECT -83.455 -86.955 -83.285 -86.630 ;
        RECT -88.435 -87.125 -87.885 -86.955 ;
        RECT -83.835 -87.125 -83.285 -86.955 ;
        RECT -83.105 -87.195 -82.735 -86.855 ;
        RECT -82.555 -86.955 -82.385 -86.630 ;
        RECT -79.415 -86.630 -78.345 -86.460 ;
        RECT -79.415 -86.955 -79.245 -86.630 ;
        RECT -82.555 -87.135 -81.625 -86.955 ;
        RECT -80.175 -87.135 -79.245 -86.955 ;
        RECT -79.065 -87.195 -78.695 -86.855 ;
        RECT -78.515 -86.955 -78.345 -86.630 ;
        RECT -73.535 -86.630 -72.465 -86.460 ;
        RECT -73.535 -86.955 -73.365 -86.630 ;
        RECT -78.515 -87.125 -77.965 -86.955 ;
        RECT -73.915 -87.125 -73.365 -86.955 ;
        RECT -73.185 -87.195 -72.815 -86.855 ;
        RECT -72.635 -86.955 -72.465 -86.630 ;
        RECT -69.495 -86.630 -68.425 -86.460 ;
        RECT -69.495 -86.955 -69.325 -86.630 ;
        RECT -72.635 -87.135 -71.705 -86.955 ;
        RECT -70.255 -87.135 -69.325 -86.955 ;
        RECT -69.145 -87.195 -68.775 -86.855 ;
        RECT -68.595 -86.955 -68.425 -86.630 ;
        RECT -63.615 -86.630 -62.545 -86.460 ;
        RECT -63.615 -86.955 -63.445 -86.630 ;
        RECT -68.595 -87.125 -68.045 -86.955 ;
        RECT -63.995 -87.125 -63.445 -86.955 ;
        RECT -63.265 -87.195 -62.895 -86.855 ;
        RECT -62.715 -86.955 -62.545 -86.630 ;
        RECT -59.575 -86.630 -58.505 -86.460 ;
        RECT -59.575 -86.955 -59.405 -86.630 ;
        RECT -62.715 -87.135 -61.785 -86.955 ;
        RECT -60.335 -87.135 -59.405 -86.955 ;
        RECT -59.225 -87.195 -58.855 -86.855 ;
        RECT -58.675 -86.955 -58.505 -86.630 ;
        RECT -53.695 -86.630 -52.625 -86.460 ;
        RECT -53.695 -86.955 -53.525 -86.630 ;
        RECT -58.675 -87.125 -58.125 -86.955 ;
        RECT -54.075 -87.125 -53.525 -86.955 ;
        RECT -53.345 -87.195 -52.975 -86.855 ;
        RECT -52.795 -86.955 -52.625 -86.630 ;
        RECT -49.655 -86.630 -48.585 -86.460 ;
        RECT -49.655 -86.955 -49.485 -86.630 ;
        RECT -52.795 -87.135 -51.865 -86.955 ;
        RECT -50.415 -87.135 -49.485 -86.955 ;
        RECT -49.305 -87.195 -48.935 -86.855 ;
        RECT -48.755 -86.955 -48.585 -86.630 ;
        RECT -43.775 -86.630 -42.705 -86.460 ;
        RECT -43.775 -86.955 -43.605 -86.630 ;
        RECT -48.755 -87.125 -48.205 -86.955 ;
        RECT -44.155 -87.125 -43.605 -86.955 ;
        RECT -43.425 -87.195 -43.055 -86.855 ;
        RECT -42.875 -86.955 -42.705 -86.630 ;
        RECT -39.735 -86.630 -38.665 -86.460 ;
        RECT -39.735 -86.955 -39.565 -86.630 ;
        RECT -42.875 -87.135 -41.945 -86.955 ;
        RECT -40.495 -87.135 -39.565 -86.955 ;
        RECT -39.385 -87.195 -39.015 -86.855 ;
        RECT -38.835 -86.955 -38.665 -86.630 ;
        RECT -33.855 -86.630 -32.785 -86.460 ;
        RECT -33.855 -86.955 -33.685 -86.630 ;
        RECT -38.835 -87.125 -38.285 -86.955 ;
        RECT -34.235 -87.125 -33.685 -86.955 ;
        RECT -33.505 -87.195 -33.135 -86.855 ;
        RECT -32.955 -86.955 -32.785 -86.630 ;
        RECT -29.815 -86.630 -28.745 -86.460 ;
        RECT -29.815 -86.955 -29.645 -86.630 ;
        RECT -32.955 -87.135 -32.025 -86.955 ;
        RECT -30.575 -87.135 -29.645 -86.955 ;
        RECT -29.465 -87.195 -29.095 -86.855 ;
        RECT -28.915 -86.955 -28.745 -86.630 ;
        RECT -23.935 -86.630 -22.865 -86.460 ;
        RECT -23.935 -86.955 -23.765 -86.630 ;
        RECT -28.915 -87.125 -28.365 -86.955 ;
        RECT -24.315 -87.125 -23.765 -86.955 ;
        RECT -23.585 -87.195 -23.215 -86.855 ;
        RECT -23.035 -86.955 -22.865 -86.630 ;
        RECT -19.895 -86.630 -18.825 -86.460 ;
        RECT -19.895 -86.955 -19.725 -86.630 ;
        RECT -23.035 -87.135 -22.105 -86.955 ;
        RECT -20.655 -87.135 -19.725 -86.955 ;
        RECT -19.545 -87.195 -19.175 -86.855 ;
        RECT -18.995 -86.955 -18.825 -86.630 ;
        RECT -14.015 -86.630 -12.945 -86.460 ;
        RECT -14.015 -86.955 -13.845 -86.630 ;
        RECT -18.995 -87.125 -18.445 -86.955 ;
        RECT -14.395 -87.125 -13.845 -86.955 ;
        RECT -13.665 -87.195 -13.295 -86.855 ;
        RECT -13.115 -86.955 -12.945 -86.630 ;
        RECT -9.975 -86.630 -8.905 -86.460 ;
        RECT -9.975 -86.955 -9.805 -86.630 ;
        RECT -13.115 -87.135 -12.185 -86.955 ;
        RECT -10.735 -87.135 -9.805 -86.955 ;
        RECT -9.625 -87.195 -9.255 -86.855 ;
        RECT -9.075 -86.955 -8.905 -86.630 ;
        RECT -4.095 -86.630 -3.025 -86.460 ;
        RECT -4.095 -86.955 -3.925 -86.630 ;
        RECT -9.075 -87.125 -8.525 -86.955 ;
        RECT -4.475 -87.125 -3.925 -86.955 ;
        RECT -3.745 -87.195 -3.375 -86.855 ;
        RECT -3.195 -86.955 -3.025 -86.630 ;
        RECT -0.055 -86.630 1.015 -86.460 ;
        RECT -0.055 -86.955 0.115 -86.630 ;
        RECT -3.195 -87.135 -2.265 -86.955 ;
        RECT -0.815 -87.135 0.115 -86.955 ;
        RECT 0.295 -87.195 0.665 -86.855 ;
        RECT 0.845 -86.955 1.015 -86.630 ;
        RECT 5.825 -86.630 6.895 -86.460 ;
        RECT 5.825 -86.955 5.995 -86.630 ;
        RECT 0.845 -87.125 1.395 -86.955 ;
        RECT 5.445 -87.125 5.995 -86.955 ;
        RECT 6.175 -87.195 6.545 -86.855 ;
        RECT 6.725 -86.955 6.895 -86.630 ;
        RECT 9.865 -86.630 10.935 -86.460 ;
        RECT 9.865 -86.955 10.035 -86.630 ;
        RECT 6.725 -87.135 7.655 -86.955 ;
        RECT 9.105 -87.135 10.035 -86.955 ;
        RECT 10.215 -87.195 10.585 -86.855 ;
        RECT 10.765 -86.955 10.935 -86.630 ;
        RECT 15.745 -86.630 16.815 -86.460 ;
        RECT 15.745 -86.955 15.915 -86.630 ;
        RECT 10.765 -87.125 11.315 -86.955 ;
        RECT 15.365 -87.125 15.915 -86.955 ;
        RECT 16.095 -87.195 16.465 -86.855 ;
        RECT 16.645 -86.955 16.815 -86.630 ;
        RECT 19.785 -86.630 20.855 -86.460 ;
        RECT 19.785 -86.955 19.955 -86.630 ;
        RECT 16.645 -87.135 17.575 -86.955 ;
        RECT 19.025 -87.135 19.955 -86.955 ;
        RECT 20.135 -87.195 20.505 -86.855 ;
        RECT 20.685 -86.955 20.855 -86.630 ;
        RECT 25.665 -86.630 26.735 -86.460 ;
        RECT 25.665 -86.955 25.835 -86.630 ;
        RECT 20.685 -87.125 21.235 -86.955 ;
        RECT 25.285 -87.125 25.835 -86.955 ;
        RECT 26.015 -87.195 26.385 -86.855 ;
        RECT 26.565 -86.955 26.735 -86.630 ;
        RECT 26.565 -87.135 27.495 -86.955 ;
        RECT -289.450 -87.815 -287.610 -87.645 ;
        RECT 26.610 -87.815 28.450 -87.645 ;
        RECT -289.365 -88.540 -289.075 -87.815 ;
        RECT -288.905 -88.615 -288.595 -87.815 ;
        RECT -288.390 -88.615 -287.695 -87.985 ;
        RECT -289.365 -90.365 -289.075 -89.200 ;
        RECT -288.390 -89.215 -288.220 -88.615 ;
        RECT -288.050 -89.055 -287.715 -88.805 ;
        RECT -285.355 -88.965 -285.025 -87.985 ;
        RECT -283.495 -88.965 -283.165 -87.985 ;
        RECT -280.825 -88.615 -280.130 -87.985 ;
        RECT -288.905 -90.365 -288.625 -89.225 ;
        RECT -288.455 -90.195 -288.125 -89.215 ;
        RECT -287.955 -90.365 -287.695 -89.225 ;
        RECT -285.765 -89.375 -285.430 -89.125 ;
        RECT -285.260 -89.565 -285.090 -88.965 ;
        RECT -285.785 -90.195 -285.090 -89.565 ;
        RECT -283.430 -89.565 -283.260 -88.965 ;
        RECT -280.805 -89.055 -280.470 -88.805 ;
        RECT -283.090 -89.375 -282.755 -89.125 ;
        RECT -280.300 -89.215 -280.130 -88.615 ;
        RECT -278.470 -88.615 -277.775 -87.985 ;
        RECT -278.470 -89.215 -278.300 -88.615 ;
        RECT -278.130 -89.055 -277.795 -88.805 ;
        RECT -275.435 -88.965 -275.105 -87.985 ;
        RECT -273.575 -88.965 -273.245 -87.985 ;
        RECT -270.905 -88.615 -270.210 -87.985 ;
        RECT -283.430 -90.195 -282.735 -89.565 ;
        RECT -280.395 -90.195 -280.065 -89.215 ;
        RECT -278.535 -90.195 -278.205 -89.215 ;
        RECT -275.845 -89.375 -275.510 -89.125 ;
        RECT -275.340 -89.565 -275.170 -88.965 ;
        RECT -275.865 -90.195 -275.170 -89.565 ;
        RECT -273.510 -89.565 -273.340 -88.965 ;
        RECT -270.885 -89.055 -270.550 -88.805 ;
        RECT -273.170 -89.375 -272.835 -89.125 ;
        RECT -270.380 -89.215 -270.210 -88.615 ;
        RECT -268.550 -88.615 -267.855 -87.985 ;
        RECT -268.550 -89.215 -268.380 -88.615 ;
        RECT -268.210 -89.055 -267.875 -88.805 ;
        RECT -265.515 -88.965 -265.185 -87.985 ;
        RECT -263.655 -88.965 -263.325 -87.985 ;
        RECT -260.985 -88.615 -260.290 -87.985 ;
        RECT -273.510 -90.195 -272.815 -89.565 ;
        RECT -270.475 -90.195 -270.145 -89.215 ;
        RECT -268.615 -90.195 -268.285 -89.215 ;
        RECT -265.925 -89.375 -265.590 -89.125 ;
        RECT -265.420 -89.565 -265.250 -88.965 ;
        RECT -265.945 -90.195 -265.250 -89.565 ;
        RECT -263.590 -89.565 -263.420 -88.965 ;
        RECT -260.965 -89.055 -260.630 -88.805 ;
        RECT -263.250 -89.375 -262.915 -89.125 ;
        RECT -260.460 -89.215 -260.290 -88.615 ;
        RECT -258.630 -88.615 -257.935 -87.985 ;
        RECT -258.630 -89.215 -258.460 -88.615 ;
        RECT -258.290 -89.055 -257.955 -88.805 ;
        RECT -255.595 -88.965 -255.265 -87.985 ;
        RECT -253.735 -88.965 -253.405 -87.985 ;
        RECT -251.065 -88.615 -250.370 -87.985 ;
        RECT -263.590 -90.195 -262.895 -89.565 ;
        RECT -260.555 -90.195 -260.225 -89.215 ;
        RECT -258.695 -90.195 -258.365 -89.215 ;
        RECT -256.005 -89.375 -255.670 -89.125 ;
        RECT -255.500 -89.565 -255.330 -88.965 ;
        RECT -256.025 -90.195 -255.330 -89.565 ;
        RECT -253.670 -89.565 -253.500 -88.965 ;
        RECT -251.045 -89.055 -250.710 -88.805 ;
        RECT -253.330 -89.375 -252.995 -89.125 ;
        RECT -250.540 -89.215 -250.370 -88.615 ;
        RECT -248.710 -88.615 -248.015 -87.985 ;
        RECT -248.710 -89.215 -248.540 -88.615 ;
        RECT -248.370 -89.055 -248.035 -88.805 ;
        RECT -245.675 -88.965 -245.345 -87.985 ;
        RECT -243.815 -88.965 -243.485 -87.985 ;
        RECT -241.145 -88.615 -240.450 -87.985 ;
        RECT -253.670 -90.195 -252.975 -89.565 ;
        RECT -250.635 -90.195 -250.305 -89.215 ;
        RECT -248.775 -90.195 -248.445 -89.215 ;
        RECT -246.085 -89.375 -245.750 -89.125 ;
        RECT -245.580 -89.565 -245.410 -88.965 ;
        RECT -246.105 -90.195 -245.410 -89.565 ;
        RECT -243.750 -89.565 -243.580 -88.965 ;
        RECT -241.125 -89.055 -240.790 -88.805 ;
        RECT -243.410 -89.375 -243.075 -89.125 ;
        RECT -240.620 -89.215 -240.450 -88.615 ;
        RECT -238.790 -88.615 -238.095 -87.985 ;
        RECT -238.790 -89.215 -238.620 -88.615 ;
        RECT -238.450 -89.055 -238.115 -88.805 ;
        RECT -235.755 -88.965 -235.425 -87.985 ;
        RECT -233.895 -88.965 -233.565 -87.985 ;
        RECT -231.225 -88.615 -230.530 -87.985 ;
        RECT -243.750 -90.195 -243.055 -89.565 ;
        RECT -240.715 -90.195 -240.385 -89.215 ;
        RECT -238.855 -90.195 -238.525 -89.215 ;
        RECT -236.165 -89.375 -235.830 -89.125 ;
        RECT -235.660 -89.565 -235.490 -88.965 ;
        RECT -236.185 -90.195 -235.490 -89.565 ;
        RECT -233.830 -89.565 -233.660 -88.965 ;
        RECT -231.205 -89.055 -230.870 -88.805 ;
        RECT -233.490 -89.375 -233.155 -89.125 ;
        RECT -230.700 -89.215 -230.530 -88.615 ;
        RECT -228.870 -88.615 -228.175 -87.985 ;
        RECT -228.870 -89.215 -228.700 -88.615 ;
        RECT -228.530 -89.055 -228.195 -88.805 ;
        RECT -225.835 -88.965 -225.505 -87.985 ;
        RECT -223.975 -88.965 -223.645 -87.985 ;
        RECT -221.305 -88.615 -220.610 -87.985 ;
        RECT -233.830 -90.195 -233.135 -89.565 ;
        RECT -230.795 -90.195 -230.465 -89.215 ;
        RECT -228.935 -90.195 -228.605 -89.215 ;
        RECT -226.245 -89.375 -225.910 -89.125 ;
        RECT -225.740 -89.565 -225.570 -88.965 ;
        RECT -226.265 -90.195 -225.570 -89.565 ;
        RECT -223.910 -89.565 -223.740 -88.965 ;
        RECT -221.285 -89.055 -220.950 -88.805 ;
        RECT -223.570 -89.375 -223.235 -89.125 ;
        RECT -220.780 -89.215 -220.610 -88.615 ;
        RECT -218.950 -88.615 -218.255 -87.985 ;
        RECT -218.950 -89.215 -218.780 -88.615 ;
        RECT -218.610 -89.055 -218.275 -88.805 ;
        RECT -215.915 -88.965 -215.585 -87.985 ;
        RECT -214.055 -88.965 -213.725 -87.985 ;
        RECT -211.385 -88.615 -210.690 -87.985 ;
        RECT -223.910 -90.195 -223.215 -89.565 ;
        RECT -220.875 -90.195 -220.545 -89.215 ;
        RECT -219.015 -90.195 -218.685 -89.215 ;
        RECT -216.325 -89.375 -215.990 -89.125 ;
        RECT -215.820 -89.565 -215.650 -88.965 ;
        RECT -216.345 -90.195 -215.650 -89.565 ;
        RECT -213.990 -89.565 -213.820 -88.965 ;
        RECT -211.365 -89.055 -211.030 -88.805 ;
        RECT -213.650 -89.375 -213.315 -89.125 ;
        RECT -210.860 -89.215 -210.690 -88.615 ;
        RECT -209.030 -88.615 -208.335 -87.985 ;
        RECT -209.030 -89.215 -208.860 -88.615 ;
        RECT -208.690 -89.055 -208.355 -88.805 ;
        RECT -205.995 -88.965 -205.665 -87.985 ;
        RECT -204.135 -88.965 -203.805 -87.985 ;
        RECT -201.465 -88.615 -200.770 -87.985 ;
        RECT -213.990 -90.195 -213.295 -89.565 ;
        RECT -210.955 -90.195 -210.625 -89.215 ;
        RECT -209.095 -90.195 -208.765 -89.215 ;
        RECT -206.405 -89.375 -206.070 -89.125 ;
        RECT -205.900 -89.565 -205.730 -88.965 ;
        RECT -206.425 -90.195 -205.730 -89.565 ;
        RECT -204.070 -89.565 -203.900 -88.965 ;
        RECT -201.445 -89.055 -201.110 -88.805 ;
        RECT -203.730 -89.375 -203.395 -89.125 ;
        RECT -200.940 -89.215 -200.770 -88.615 ;
        RECT -199.110 -88.615 -198.415 -87.985 ;
        RECT -199.110 -89.215 -198.940 -88.615 ;
        RECT -198.770 -89.055 -198.435 -88.805 ;
        RECT -196.075 -88.965 -195.745 -87.985 ;
        RECT -194.215 -88.965 -193.885 -87.985 ;
        RECT -191.545 -88.615 -190.850 -87.985 ;
        RECT -204.070 -90.195 -203.375 -89.565 ;
        RECT -201.035 -90.195 -200.705 -89.215 ;
        RECT -199.175 -90.195 -198.845 -89.215 ;
        RECT -196.485 -89.375 -196.150 -89.125 ;
        RECT -195.980 -89.565 -195.810 -88.965 ;
        RECT -196.505 -90.195 -195.810 -89.565 ;
        RECT -194.150 -89.565 -193.980 -88.965 ;
        RECT -191.525 -89.055 -191.190 -88.805 ;
        RECT -193.810 -89.375 -193.475 -89.125 ;
        RECT -191.020 -89.215 -190.850 -88.615 ;
        RECT -189.190 -88.615 -188.495 -87.985 ;
        RECT -189.190 -89.215 -189.020 -88.615 ;
        RECT -188.850 -89.055 -188.515 -88.805 ;
        RECT -186.155 -88.965 -185.825 -87.985 ;
        RECT -184.295 -88.965 -183.965 -87.985 ;
        RECT -181.625 -88.615 -180.930 -87.985 ;
        RECT -194.150 -90.195 -193.455 -89.565 ;
        RECT -191.115 -90.195 -190.785 -89.215 ;
        RECT -189.255 -90.195 -188.925 -89.215 ;
        RECT -186.565 -89.375 -186.230 -89.125 ;
        RECT -186.060 -89.565 -185.890 -88.965 ;
        RECT -186.585 -90.195 -185.890 -89.565 ;
        RECT -184.230 -89.565 -184.060 -88.965 ;
        RECT -181.605 -89.055 -181.270 -88.805 ;
        RECT -183.890 -89.375 -183.555 -89.125 ;
        RECT -181.100 -89.215 -180.930 -88.615 ;
        RECT -179.270 -88.615 -178.575 -87.985 ;
        RECT -179.270 -89.215 -179.100 -88.615 ;
        RECT -178.930 -89.055 -178.595 -88.805 ;
        RECT -176.235 -88.965 -175.905 -87.985 ;
        RECT -174.375 -88.965 -174.045 -87.985 ;
        RECT -171.705 -88.615 -171.010 -87.985 ;
        RECT -184.230 -90.195 -183.535 -89.565 ;
        RECT -181.195 -90.195 -180.865 -89.215 ;
        RECT -179.335 -90.195 -179.005 -89.215 ;
        RECT -176.645 -89.375 -176.310 -89.125 ;
        RECT -176.140 -89.565 -175.970 -88.965 ;
        RECT -176.665 -90.195 -175.970 -89.565 ;
        RECT -174.310 -89.565 -174.140 -88.965 ;
        RECT -171.685 -89.055 -171.350 -88.805 ;
        RECT -173.970 -89.375 -173.635 -89.125 ;
        RECT -171.180 -89.215 -171.010 -88.615 ;
        RECT -169.350 -88.615 -168.655 -87.985 ;
        RECT -169.350 -89.215 -169.180 -88.615 ;
        RECT -169.010 -89.055 -168.675 -88.805 ;
        RECT -166.315 -88.965 -165.985 -87.985 ;
        RECT -164.455 -88.965 -164.125 -87.985 ;
        RECT -161.785 -88.615 -161.090 -87.985 ;
        RECT -174.310 -90.195 -173.615 -89.565 ;
        RECT -171.275 -90.195 -170.945 -89.215 ;
        RECT -169.415 -90.195 -169.085 -89.215 ;
        RECT -166.725 -89.375 -166.390 -89.125 ;
        RECT -166.220 -89.565 -166.050 -88.965 ;
        RECT -166.745 -90.195 -166.050 -89.565 ;
        RECT -164.390 -89.565 -164.220 -88.965 ;
        RECT -161.765 -89.055 -161.430 -88.805 ;
        RECT -164.050 -89.375 -163.715 -89.125 ;
        RECT -161.260 -89.215 -161.090 -88.615 ;
        RECT -159.430 -88.615 -158.735 -87.985 ;
        RECT -159.430 -89.215 -159.260 -88.615 ;
        RECT -159.090 -89.055 -158.755 -88.805 ;
        RECT -156.395 -88.965 -156.065 -87.985 ;
        RECT -154.535 -88.965 -154.205 -87.985 ;
        RECT -151.865 -88.615 -151.170 -87.985 ;
        RECT -164.390 -90.195 -163.695 -89.565 ;
        RECT -161.355 -90.195 -161.025 -89.215 ;
        RECT -159.495 -90.195 -159.165 -89.215 ;
        RECT -156.805 -89.375 -156.470 -89.125 ;
        RECT -156.300 -89.565 -156.130 -88.965 ;
        RECT -156.825 -90.195 -156.130 -89.565 ;
        RECT -154.470 -89.565 -154.300 -88.965 ;
        RECT -151.845 -89.055 -151.510 -88.805 ;
        RECT -154.130 -89.375 -153.795 -89.125 ;
        RECT -151.340 -89.215 -151.170 -88.615 ;
        RECT -149.510 -88.615 -148.815 -87.985 ;
        RECT -149.510 -89.215 -149.340 -88.615 ;
        RECT -149.170 -89.055 -148.835 -88.805 ;
        RECT -146.475 -88.965 -146.145 -87.985 ;
        RECT -144.615 -88.965 -144.285 -87.985 ;
        RECT -141.945 -88.615 -141.250 -87.985 ;
        RECT -154.470 -90.195 -153.775 -89.565 ;
        RECT -151.435 -90.195 -151.105 -89.215 ;
        RECT -149.575 -90.195 -149.245 -89.215 ;
        RECT -146.885 -89.375 -146.550 -89.125 ;
        RECT -146.380 -89.565 -146.210 -88.965 ;
        RECT -146.905 -90.195 -146.210 -89.565 ;
        RECT -144.550 -89.565 -144.380 -88.965 ;
        RECT -141.925 -89.055 -141.590 -88.805 ;
        RECT -144.210 -89.375 -143.875 -89.125 ;
        RECT -141.420 -89.215 -141.250 -88.615 ;
        RECT -139.590 -88.615 -138.895 -87.985 ;
        RECT -139.590 -89.215 -139.420 -88.615 ;
        RECT -139.250 -89.055 -138.915 -88.805 ;
        RECT -136.555 -88.965 -136.225 -87.985 ;
        RECT -134.695 -88.965 -134.365 -87.985 ;
        RECT -132.025 -88.615 -131.330 -87.985 ;
        RECT -144.550 -90.195 -143.855 -89.565 ;
        RECT -141.515 -90.195 -141.185 -89.215 ;
        RECT -139.655 -90.195 -139.325 -89.215 ;
        RECT -136.965 -89.375 -136.630 -89.125 ;
        RECT -136.460 -89.565 -136.290 -88.965 ;
        RECT -136.985 -90.195 -136.290 -89.565 ;
        RECT -134.630 -89.565 -134.460 -88.965 ;
        RECT -132.005 -89.055 -131.670 -88.805 ;
        RECT -134.290 -89.375 -133.955 -89.125 ;
        RECT -131.500 -89.215 -131.330 -88.615 ;
        RECT -129.670 -88.615 -128.975 -87.985 ;
        RECT -129.670 -89.215 -129.500 -88.615 ;
        RECT -129.330 -89.055 -128.995 -88.805 ;
        RECT -126.635 -88.965 -126.305 -87.985 ;
        RECT -124.775 -88.965 -124.445 -87.985 ;
        RECT -122.105 -88.615 -121.410 -87.985 ;
        RECT -134.630 -90.195 -133.935 -89.565 ;
        RECT -131.595 -90.195 -131.265 -89.215 ;
        RECT -129.735 -90.195 -129.405 -89.215 ;
        RECT -127.045 -89.375 -126.710 -89.125 ;
        RECT -126.540 -89.565 -126.370 -88.965 ;
        RECT -127.065 -90.195 -126.370 -89.565 ;
        RECT -124.710 -89.565 -124.540 -88.965 ;
        RECT -122.085 -89.055 -121.750 -88.805 ;
        RECT -124.370 -89.375 -124.035 -89.125 ;
        RECT -121.580 -89.215 -121.410 -88.615 ;
        RECT -119.750 -88.615 -119.055 -87.985 ;
        RECT -119.750 -89.215 -119.580 -88.615 ;
        RECT -119.410 -89.055 -119.075 -88.805 ;
        RECT -116.715 -88.965 -116.385 -87.985 ;
        RECT -114.855 -88.965 -114.525 -87.985 ;
        RECT -112.185 -88.615 -111.490 -87.985 ;
        RECT -124.710 -90.195 -124.015 -89.565 ;
        RECT -121.675 -90.195 -121.345 -89.215 ;
        RECT -119.815 -90.195 -119.485 -89.215 ;
        RECT -117.125 -89.375 -116.790 -89.125 ;
        RECT -116.620 -89.565 -116.450 -88.965 ;
        RECT -117.145 -90.195 -116.450 -89.565 ;
        RECT -114.790 -89.565 -114.620 -88.965 ;
        RECT -112.165 -89.055 -111.830 -88.805 ;
        RECT -114.450 -89.375 -114.115 -89.125 ;
        RECT -111.660 -89.215 -111.490 -88.615 ;
        RECT -109.830 -88.615 -109.135 -87.985 ;
        RECT -109.830 -89.215 -109.660 -88.615 ;
        RECT -109.490 -89.055 -109.155 -88.805 ;
        RECT -106.795 -88.965 -106.465 -87.985 ;
        RECT -104.935 -88.965 -104.605 -87.985 ;
        RECT -102.265 -88.615 -101.570 -87.985 ;
        RECT -114.790 -90.195 -114.095 -89.565 ;
        RECT -111.755 -90.195 -111.425 -89.215 ;
        RECT -109.895 -90.195 -109.565 -89.215 ;
        RECT -107.205 -89.375 -106.870 -89.125 ;
        RECT -106.700 -89.565 -106.530 -88.965 ;
        RECT -107.225 -90.195 -106.530 -89.565 ;
        RECT -104.870 -89.565 -104.700 -88.965 ;
        RECT -102.245 -89.055 -101.910 -88.805 ;
        RECT -104.530 -89.375 -104.195 -89.125 ;
        RECT -101.740 -89.215 -101.570 -88.615 ;
        RECT -99.910 -88.615 -99.215 -87.985 ;
        RECT -99.910 -89.215 -99.740 -88.615 ;
        RECT -99.570 -89.055 -99.235 -88.805 ;
        RECT -96.875 -88.965 -96.545 -87.985 ;
        RECT -95.015 -88.965 -94.685 -87.985 ;
        RECT -92.345 -88.615 -91.650 -87.985 ;
        RECT -104.870 -90.195 -104.175 -89.565 ;
        RECT -101.835 -90.195 -101.505 -89.215 ;
        RECT -99.975 -90.195 -99.645 -89.215 ;
        RECT -97.285 -89.375 -96.950 -89.125 ;
        RECT -96.780 -89.565 -96.610 -88.965 ;
        RECT -97.305 -90.195 -96.610 -89.565 ;
        RECT -94.950 -89.565 -94.780 -88.965 ;
        RECT -92.325 -89.055 -91.990 -88.805 ;
        RECT -94.610 -89.375 -94.275 -89.125 ;
        RECT -91.820 -89.215 -91.650 -88.615 ;
        RECT -89.990 -88.615 -89.295 -87.985 ;
        RECT -89.990 -89.215 -89.820 -88.615 ;
        RECT -89.650 -89.055 -89.315 -88.805 ;
        RECT -86.955 -88.965 -86.625 -87.985 ;
        RECT -85.095 -88.965 -84.765 -87.985 ;
        RECT -82.425 -88.615 -81.730 -87.985 ;
        RECT -94.950 -90.195 -94.255 -89.565 ;
        RECT -91.915 -90.195 -91.585 -89.215 ;
        RECT -90.055 -90.195 -89.725 -89.215 ;
        RECT -87.365 -89.375 -87.030 -89.125 ;
        RECT -86.860 -89.565 -86.690 -88.965 ;
        RECT -87.385 -90.195 -86.690 -89.565 ;
        RECT -85.030 -89.565 -84.860 -88.965 ;
        RECT -82.405 -89.055 -82.070 -88.805 ;
        RECT -84.690 -89.375 -84.355 -89.125 ;
        RECT -81.900 -89.215 -81.730 -88.615 ;
        RECT -80.070 -88.615 -79.375 -87.985 ;
        RECT -80.070 -89.215 -79.900 -88.615 ;
        RECT -79.730 -89.055 -79.395 -88.805 ;
        RECT -77.035 -88.965 -76.705 -87.985 ;
        RECT -75.175 -88.965 -74.845 -87.985 ;
        RECT -72.505 -88.615 -71.810 -87.985 ;
        RECT -85.030 -90.195 -84.335 -89.565 ;
        RECT -81.995 -90.195 -81.665 -89.215 ;
        RECT -80.135 -90.195 -79.805 -89.215 ;
        RECT -77.445 -89.375 -77.110 -89.125 ;
        RECT -76.940 -89.565 -76.770 -88.965 ;
        RECT -77.465 -90.195 -76.770 -89.565 ;
        RECT -75.110 -89.565 -74.940 -88.965 ;
        RECT -72.485 -89.055 -72.150 -88.805 ;
        RECT -74.770 -89.375 -74.435 -89.125 ;
        RECT -71.980 -89.215 -71.810 -88.615 ;
        RECT -70.150 -88.615 -69.455 -87.985 ;
        RECT -70.150 -89.215 -69.980 -88.615 ;
        RECT -69.810 -89.055 -69.475 -88.805 ;
        RECT -67.115 -88.965 -66.785 -87.985 ;
        RECT -65.255 -88.965 -64.925 -87.985 ;
        RECT -62.585 -88.615 -61.890 -87.985 ;
        RECT -75.110 -90.195 -74.415 -89.565 ;
        RECT -72.075 -90.195 -71.745 -89.215 ;
        RECT -70.215 -90.195 -69.885 -89.215 ;
        RECT -67.525 -89.375 -67.190 -89.125 ;
        RECT -67.020 -89.565 -66.850 -88.965 ;
        RECT -67.545 -90.195 -66.850 -89.565 ;
        RECT -65.190 -89.565 -65.020 -88.965 ;
        RECT -62.565 -89.055 -62.230 -88.805 ;
        RECT -64.850 -89.375 -64.515 -89.125 ;
        RECT -62.060 -89.215 -61.890 -88.615 ;
        RECT -60.230 -88.615 -59.535 -87.985 ;
        RECT -60.230 -89.215 -60.060 -88.615 ;
        RECT -59.890 -89.055 -59.555 -88.805 ;
        RECT -57.195 -88.965 -56.865 -87.985 ;
        RECT -55.335 -88.965 -55.005 -87.985 ;
        RECT -52.665 -88.615 -51.970 -87.985 ;
        RECT -65.190 -90.195 -64.495 -89.565 ;
        RECT -62.155 -90.195 -61.825 -89.215 ;
        RECT -60.295 -90.195 -59.965 -89.215 ;
        RECT -57.605 -89.375 -57.270 -89.125 ;
        RECT -57.100 -89.565 -56.930 -88.965 ;
        RECT -57.625 -90.195 -56.930 -89.565 ;
        RECT -55.270 -89.565 -55.100 -88.965 ;
        RECT -52.645 -89.055 -52.310 -88.805 ;
        RECT -54.930 -89.375 -54.595 -89.125 ;
        RECT -52.140 -89.215 -51.970 -88.615 ;
        RECT -50.310 -88.615 -49.615 -87.985 ;
        RECT -50.310 -89.215 -50.140 -88.615 ;
        RECT -49.970 -89.055 -49.635 -88.805 ;
        RECT -47.275 -88.965 -46.945 -87.985 ;
        RECT -45.415 -88.965 -45.085 -87.985 ;
        RECT -42.745 -88.615 -42.050 -87.985 ;
        RECT -55.270 -90.195 -54.575 -89.565 ;
        RECT -52.235 -90.195 -51.905 -89.215 ;
        RECT -50.375 -90.195 -50.045 -89.215 ;
        RECT -47.685 -89.375 -47.350 -89.125 ;
        RECT -47.180 -89.565 -47.010 -88.965 ;
        RECT -47.705 -90.195 -47.010 -89.565 ;
        RECT -45.350 -89.565 -45.180 -88.965 ;
        RECT -42.725 -89.055 -42.390 -88.805 ;
        RECT -45.010 -89.375 -44.675 -89.125 ;
        RECT -42.220 -89.215 -42.050 -88.615 ;
        RECT -40.390 -88.615 -39.695 -87.985 ;
        RECT -40.390 -89.215 -40.220 -88.615 ;
        RECT -40.050 -89.055 -39.715 -88.805 ;
        RECT -37.355 -88.965 -37.025 -87.985 ;
        RECT -35.495 -88.965 -35.165 -87.985 ;
        RECT -32.825 -88.615 -32.130 -87.985 ;
        RECT -45.350 -90.195 -44.655 -89.565 ;
        RECT -42.315 -90.195 -41.985 -89.215 ;
        RECT -40.455 -90.195 -40.125 -89.215 ;
        RECT -37.765 -89.375 -37.430 -89.125 ;
        RECT -37.260 -89.565 -37.090 -88.965 ;
        RECT -37.785 -90.195 -37.090 -89.565 ;
        RECT -35.430 -89.565 -35.260 -88.965 ;
        RECT -32.805 -89.055 -32.470 -88.805 ;
        RECT -35.090 -89.375 -34.755 -89.125 ;
        RECT -32.300 -89.215 -32.130 -88.615 ;
        RECT -30.470 -88.615 -29.775 -87.985 ;
        RECT -30.470 -89.215 -30.300 -88.615 ;
        RECT -30.130 -89.055 -29.795 -88.805 ;
        RECT -27.435 -88.965 -27.105 -87.985 ;
        RECT -25.575 -88.965 -25.245 -87.985 ;
        RECT -22.905 -88.615 -22.210 -87.985 ;
        RECT -35.430 -90.195 -34.735 -89.565 ;
        RECT -32.395 -90.195 -32.065 -89.215 ;
        RECT -30.535 -90.195 -30.205 -89.215 ;
        RECT -27.845 -89.375 -27.510 -89.125 ;
        RECT -27.340 -89.565 -27.170 -88.965 ;
        RECT -27.865 -90.195 -27.170 -89.565 ;
        RECT -25.510 -89.565 -25.340 -88.965 ;
        RECT -22.885 -89.055 -22.550 -88.805 ;
        RECT -25.170 -89.375 -24.835 -89.125 ;
        RECT -22.380 -89.215 -22.210 -88.615 ;
        RECT -20.550 -88.615 -19.855 -87.985 ;
        RECT -20.550 -89.215 -20.380 -88.615 ;
        RECT -20.210 -89.055 -19.875 -88.805 ;
        RECT -17.515 -88.965 -17.185 -87.985 ;
        RECT -15.655 -88.965 -15.325 -87.985 ;
        RECT -12.985 -88.615 -12.290 -87.985 ;
        RECT -25.510 -90.195 -24.815 -89.565 ;
        RECT -22.475 -90.195 -22.145 -89.215 ;
        RECT -20.615 -90.195 -20.285 -89.215 ;
        RECT -17.925 -89.375 -17.590 -89.125 ;
        RECT -17.420 -89.565 -17.250 -88.965 ;
        RECT -17.945 -90.195 -17.250 -89.565 ;
        RECT -15.590 -89.565 -15.420 -88.965 ;
        RECT -12.965 -89.055 -12.630 -88.805 ;
        RECT -15.250 -89.375 -14.915 -89.125 ;
        RECT -12.460 -89.215 -12.290 -88.615 ;
        RECT -10.630 -88.615 -9.935 -87.985 ;
        RECT -10.630 -89.215 -10.460 -88.615 ;
        RECT -10.290 -89.055 -9.955 -88.805 ;
        RECT -7.595 -88.965 -7.265 -87.985 ;
        RECT -5.735 -88.965 -5.405 -87.985 ;
        RECT -3.065 -88.615 -2.370 -87.985 ;
        RECT -15.590 -90.195 -14.895 -89.565 ;
        RECT -12.555 -90.195 -12.225 -89.215 ;
        RECT -10.695 -90.195 -10.365 -89.215 ;
        RECT -8.005 -89.375 -7.670 -89.125 ;
        RECT -7.500 -89.565 -7.330 -88.965 ;
        RECT -8.025 -90.195 -7.330 -89.565 ;
        RECT -5.670 -89.565 -5.500 -88.965 ;
        RECT -3.045 -89.055 -2.710 -88.805 ;
        RECT -5.330 -89.375 -4.995 -89.125 ;
        RECT -2.540 -89.215 -2.370 -88.615 ;
        RECT -0.710 -88.615 -0.015 -87.985 ;
        RECT -0.710 -89.215 -0.540 -88.615 ;
        RECT -0.370 -89.055 -0.035 -88.805 ;
        RECT 2.325 -88.965 2.655 -87.985 ;
        RECT 4.185 -88.965 4.515 -87.985 ;
        RECT 6.855 -88.615 7.550 -87.985 ;
        RECT -5.670 -90.195 -4.975 -89.565 ;
        RECT -2.635 -90.195 -2.305 -89.215 ;
        RECT -0.775 -90.195 -0.445 -89.215 ;
        RECT 1.915 -89.375 2.250 -89.125 ;
        RECT 2.420 -89.565 2.590 -88.965 ;
        RECT 1.895 -90.195 2.590 -89.565 ;
        RECT 4.250 -89.565 4.420 -88.965 ;
        RECT 6.875 -89.055 7.210 -88.805 ;
        RECT 4.590 -89.375 4.925 -89.125 ;
        RECT 7.380 -89.215 7.550 -88.615 ;
        RECT 9.210 -88.615 9.905 -87.985 ;
        RECT 9.210 -89.215 9.380 -88.615 ;
        RECT 9.550 -89.055 9.885 -88.805 ;
        RECT 12.245 -88.965 12.575 -87.985 ;
        RECT 14.105 -88.965 14.435 -87.985 ;
        RECT 16.775 -88.615 17.470 -87.985 ;
        RECT 4.250 -90.195 4.945 -89.565 ;
        RECT 7.285 -90.195 7.615 -89.215 ;
        RECT 9.145 -90.195 9.475 -89.215 ;
        RECT 11.835 -89.375 12.170 -89.125 ;
        RECT 12.340 -89.565 12.510 -88.965 ;
        RECT 11.815 -90.195 12.510 -89.565 ;
        RECT 14.170 -89.565 14.340 -88.965 ;
        RECT 16.795 -89.055 17.130 -88.805 ;
        RECT 14.510 -89.375 14.845 -89.125 ;
        RECT 17.300 -89.215 17.470 -88.615 ;
        RECT 19.130 -88.615 19.825 -87.985 ;
        RECT 19.130 -89.215 19.300 -88.615 ;
        RECT 19.470 -89.055 19.805 -88.805 ;
        RECT 22.165 -88.965 22.495 -87.985 ;
        RECT 24.025 -88.965 24.355 -87.985 ;
        RECT 26.695 -88.615 27.390 -87.985 ;
        RECT 27.595 -88.615 27.905 -87.815 ;
        RECT 28.075 -88.540 28.365 -87.815 ;
        RECT 14.170 -90.195 14.865 -89.565 ;
        RECT 17.205 -90.195 17.535 -89.215 ;
        RECT 19.065 -90.195 19.395 -89.215 ;
        RECT 21.755 -89.375 22.090 -89.125 ;
        RECT 22.260 -89.565 22.430 -88.965 ;
        RECT 21.735 -90.195 22.430 -89.565 ;
        RECT 24.090 -89.565 24.260 -88.965 ;
        RECT 26.715 -89.055 27.050 -88.805 ;
        RECT 24.430 -89.375 24.765 -89.125 ;
        RECT 27.220 -89.215 27.390 -88.615 ;
        RECT 24.090 -90.195 24.785 -89.565 ;
        RECT 27.125 -90.195 27.455 -89.215 ;
        RECT -289.450 -90.535 -287.610 -90.365 ;
        RECT -288.065 -91.920 -287.775 -91.210 ;
        RECT -287.535 -91.405 -287.365 -90.880 ;
        RECT -287.195 -91.225 -286.645 -91.055 ;
        RECT -287.535 -91.735 -286.985 -91.405 ;
        RECT -286.815 -91.550 -286.645 -91.225 ;
        RECT -286.465 -91.325 -286.095 -90.985 ;
        RECT -285.915 -91.225 -284.985 -91.045 ;
        RECT -283.535 -91.225 -282.605 -91.045 ;
        RECT -285.915 -91.550 -285.745 -91.225 ;
        RECT -286.815 -91.720 -285.745 -91.550 ;
        RECT -282.775 -91.550 -282.605 -91.225 ;
        RECT -282.425 -91.325 -282.055 -90.985 ;
        RECT -281.875 -91.225 -281.325 -91.055 ;
        RECT -277.275 -91.225 -276.725 -91.055 ;
        RECT -281.875 -91.550 -281.705 -91.225 ;
        RECT -282.775 -91.720 -281.705 -91.550 ;
        RECT -276.895 -91.550 -276.725 -91.225 ;
        RECT -276.545 -91.325 -276.175 -90.985 ;
        RECT -275.995 -91.225 -275.065 -91.045 ;
        RECT -273.615 -91.225 -272.685 -91.045 ;
        RECT -275.995 -91.550 -275.825 -91.225 ;
        RECT -276.895 -91.720 -275.825 -91.550 ;
        RECT -272.855 -91.550 -272.685 -91.225 ;
        RECT -272.505 -91.325 -272.135 -90.985 ;
        RECT -271.955 -91.225 -271.405 -91.055 ;
        RECT -267.355 -91.225 -266.805 -91.055 ;
        RECT -271.955 -91.550 -271.785 -91.225 ;
        RECT -272.855 -91.720 -271.785 -91.550 ;
        RECT -266.975 -91.550 -266.805 -91.225 ;
        RECT -266.625 -91.325 -266.255 -90.985 ;
        RECT -266.075 -91.225 -265.145 -91.045 ;
        RECT -263.695 -91.225 -262.765 -91.045 ;
        RECT -266.075 -91.550 -265.905 -91.225 ;
        RECT -266.975 -91.720 -265.905 -91.550 ;
        RECT -262.935 -91.550 -262.765 -91.225 ;
        RECT -262.585 -91.325 -262.215 -90.985 ;
        RECT -262.035 -91.225 -261.485 -91.055 ;
        RECT -257.435 -91.225 -256.885 -91.055 ;
        RECT -262.035 -91.550 -261.865 -91.225 ;
        RECT -262.935 -91.720 -261.865 -91.550 ;
        RECT -257.055 -91.550 -256.885 -91.225 ;
        RECT -256.705 -91.325 -256.335 -90.985 ;
        RECT -256.155 -91.225 -255.225 -91.045 ;
        RECT -253.775 -91.225 -252.845 -91.045 ;
        RECT -256.155 -91.550 -255.985 -91.225 ;
        RECT -257.055 -91.720 -255.985 -91.550 ;
        RECT -253.015 -91.550 -252.845 -91.225 ;
        RECT -252.665 -91.325 -252.295 -90.985 ;
        RECT -252.115 -91.225 -251.565 -91.055 ;
        RECT -247.515 -91.225 -246.965 -91.055 ;
        RECT -252.115 -91.550 -251.945 -91.225 ;
        RECT -253.015 -91.720 -251.945 -91.550 ;
        RECT -247.135 -91.550 -246.965 -91.225 ;
        RECT -246.785 -91.325 -246.415 -90.985 ;
        RECT -246.235 -91.225 -245.305 -91.045 ;
        RECT -243.855 -91.225 -242.925 -91.045 ;
        RECT -246.235 -91.550 -246.065 -91.225 ;
        RECT -247.135 -91.720 -246.065 -91.550 ;
        RECT -243.095 -91.550 -242.925 -91.225 ;
        RECT -242.745 -91.325 -242.375 -90.985 ;
        RECT -242.195 -91.225 -241.645 -91.055 ;
        RECT -237.595 -91.225 -237.045 -91.055 ;
        RECT -242.195 -91.550 -242.025 -91.225 ;
        RECT -243.095 -91.720 -242.025 -91.550 ;
        RECT -237.215 -91.550 -237.045 -91.225 ;
        RECT -236.865 -91.325 -236.495 -90.985 ;
        RECT -236.315 -91.225 -235.385 -91.045 ;
        RECT -233.935 -91.225 -233.005 -91.045 ;
        RECT -236.315 -91.550 -236.145 -91.225 ;
        RECT -237.215 -91.720 -236.145 -91.550 ;
        RECT -233.175 -91.550 -233.005 -91.225 ;
        RECT -232.825 -91.325 -232.455 -90.985 ;
        RECT -232.275 -91.225 -231.725 -91.055 ;
        RECT -227.675 -91.225 -227.125 -91.055 ;
        RECT -232.275 -91.550 -232.105 -91.225 ;
        RECT -233.175 -91.720 -232.105 -91.550 ;
        RECT -227.295 -91.550 -227.125 -91.225 ;
        RECT -226.945 -91.325 -226.575 -90.985 ;
        RECT -226.395 -91.225 -225.465 -91.045 ;
        RECT -224.015 -91.225 -223.085 -91.045 ;
        RECT -226.395 -91.550 -226.225 -91.225 ;
        RECT -227.295 -91.720 -226.225 -91.550 ;
        RECT -223.255 -91.550 -223.085 -91.225 ;
        RECT -222.905 -91.325 -222.535 -90.985 ;
        RECT -222.355 -91.225 -221.805 -91.055 ;
        RECT -217.755 -91.225 -217.205 -91.055 ;
        RECT -222.355 -91.550 -222.185 -91.225 ;
        RECT -223.255 -91.720 -222.185 -91.550 ;
        RECT -217.375 -91.550 -217.205 -91.225 ;
        RECT -217.025 -91.325 -216.655 -90.985 ;
        RECT -216.475 -91.225 -215.545 -91.045 ;
        RECT -214.095 -91.225 -213.165 -91.045 ;
        RECT -216.475 -91.550 -216.305 -91.225 ;
        RECT -217.375 -91.720 -216.305 -91.550 ;
        RECT -213.335 -91.550 -213.165 -91.225 ;
        RECT -212.985 -91.325 -212.615 -90.985 ;
        RECT -212.435 -91.225 -211.885 -91.055 ;
        RECT -207.835 -91.225 -207.285 -91.055 ;
        RECT -212.435 -91.550 -212.265 -91.225 ;
        RECT -213.335 -91.720 -212.265 -91.550 ;
        RECT -207.455 -91.550 -207.285 -91.225 ;
        RECT -207.105 -91.325 -206.735 -90.985 ;
        RECT -206.555 -91.225 -205.625 -91.045 ;
        RECT -204.175 -91.225 -203.245 -91.045 ;
        RECT -206.555 -91.550 -206.385 -91.225 ;
        RECT -207.455 -91.720 -206.385 -91.550 ;
        RECT -203.415 -91.550 -203.245 -91.225 ;
        RECT -203.065 -91.325 -202.695 -90.985 ;
        RECT -202.515 -91.225 -201.965 -91.055 ;
        RECT -197.915 -91.225 -197.365 -91.055 ;
        RECT -202.515 -91.550 -202.345 -91.225 ;
        RECT -203.415 -91.720 -202.345 -91.550 ;
        RECT -197.535 -91.550 -197.365 -91.225 ;
        RECT -197.185 -91.325 -196.815 -90.985 ;
        RECT -196.635 -91.225 -195.705 -91.045 ;
        RECT -194.255 -91.225 -193.325 -91.045 ;
        RECT -196.635 -91.550 -196.465 -91.225 ;
        RECT -197.535 -91.720 -196.465 -91.550 ;
        RECT -193.495 -91.550 -193.325 -91.225 ;
        RECT -193.145 -91.325 -192.775 -90.985 ;
        RECT -192.595 -91.225 -192.045 -91.055 ;
        RECT -187.995 -91.225 -187.445 -91.055 ;
        RECT -192.595 -91.550 -192.425 -91.225 ;
        RECT -193.495 -91.720 -192.425 -91.550 ;
        RECT -187.615 -91.550 -187.445 -91.225 ;
        RECT -187.265 -91.325 -186.895 -90.985 ;
        RECT -186.715 -91.225 -185.785 -91.045 ;
        RECT -184.335 -91.225 -183.405 -91.045 ;
        RECT -186.715 -91.550 -186.545 -91.225 ;
        RECT -187.615 -91.720 -186.545 -91.550 ;
        RECT -183.575 -91.550 -183.405 -91.225 ;
        RECT -183.225 -91.325 -182.855 -90.985 ;
        RECT -182.675 -91.225 -182.125 -91.055 ;
        RECT -178.075 -91.225 -177.525 -91.055 ;
        RECT -182.675 -91.550 -182.505 -91.225 ;
        RECT -183.575 -91.720 -182.505 -91.550 ;
        RECT -177.695 -91.550 -177.525 -91.225 ;
        RECT -177.345 -91.325 -176.975 -90.985 ;
        RECT -176.795 -91.225 -175.865 -91.045 ;
        RECT -174.415 -91.225 -173.485 -91.045 ;
        RECT -176.795 -91.550 -176.625 -91.225 ;
        RECT -177.695 -91.720 -176.625 -91.550 ;
        RECT -173.655 -91.550 -173.485 -91.225 ;
        RECT -173.305 -91.325 -172.935 -90.985 ;
        RECT -172.755 -91.225 -172.205 -91.055 ;
        RECT -168.155 -91.225 -167.605 -91.055 ;
        RECT -172.755 -91.550 -172.585 -91.225 ;
        RECT -173.655 -91.720 -172.585 -91.550 ;
        RECT -167.775 -91.550 -167.605 -91.225 ;
        RECT -167.425 -91.325 -167.055 -90.985 ;
        RECT -166.875 -91.225 -165.945 -91.045 ;
        RECT -164.495 -91.225 -163.565 -91.045 ;
        RECT -166.875 -91.550 -166.705 -91.225 ;
        RECT -167.775 -91.720 -166.705 -91.550 ;
        RECT -163.735 -91.550 -163.565 -91.225 ;
        RECT -163.385 -91.325 -163.015 -90.985 ;
        RECT -162.835 -91.225 -162.285 -91.055 ;
        RECT -158.235 -91.225 -157.685 -91.055 ;
        RECT -162.835 -91.550 -162.665 -91.225 ;
        RECT -163.735 -91.720 -162.665 -91.550 ;
        RECT -157.855 -91.550 -157.685 -91.225 ;
        RECT -157.505 -91.325 -157.135 -90.985 ;
        RECT -156.955 -91.225 -156.025 -91.045 ;
        RECT -154.575 -91.225 -153.645 -91.045 ;
        RECT -156.955 -91.550 -156.785 -91.225 ;
        RECT -157.855 -91.720 -156.785 -91.550 ;
        RECT -153.815 -91.550 -153.645 -91.225 ;
        RECT -153.465 -91.325 -153.095 -90.985 ;
        RECT -152.915 -91.225 -152.365 -91.055 ;
        RECT -148.315 -91.225 -147.765 -91.055 ;
        RECT -152.915 -91.550 -152.745 -91.225 ;
        RECT -153.815 -91.720 -152.745 -91.550 ;
        RECT -147.935 -91.550 -147.765 -91.225 ;
        RECT -147.585 -91.325 -147.215 -90.985 ;
        RECT -147.035 -91.225 -146.105 -91.045 ;
        RECT -144.655 -91.225 -143.725 -91.045 ;
        RECT -147.035 -91.550 -146.865 -91.225 ;
        RECT -147.935 -91.720 -146.865 -91.550 ;
        RECT -143.895 -91.550 -143.725 -91.225 ;
        RECT -143.545 -91.325 -143.175 -90.985 ;
        RECT -142.995 -91.225 -142.445 -91.055 ;
        RECT -138.395 -91.225 -137.845 -91.055 ;
        RECT -142.995 -91.550 -142.825 -91.225 ;
        RECT -143.895 -91.720 -142.825 -91.550 ;
        RECT -138.015 -91.550 -137.845 -91.225 ;
        RECT -137.665 -91.325 -137.295 -90.985 ;
        RECT -137.115 -91.225 -136.185 -91.045 ;
        RECT -134.735 -91.225 -133.805 -91.045 ;
        RECT -137.115 -91.550 -136.945 -91.225 ;
        RECT -138.015 -91.720 -136.945 -91.550 ;
        RECT -133.975 -91.550 -133.805 -91.225 ;
        RECT -133.625 -91.325 -133.255 -90.985 ;
        RECT -133.075 -91.225 -132.525 -91.055 ;
        RECT -128.475 -91.225 -127.925 -91.055 ;
        RECT -133.075 -91.550 -132.905 -91.225 ;
        RECT -133.975 -91.720 -132.905 -91.550 ;
        RECT -128.095 -91.550 -127.925 -91.225 ;
        RECT -127.745 -91.325 -127.375 -90.985 ;
        RECT -127.195 -91.225 -126.265 -91.045 ;
        RECT -124.815 -91.225 -123.885 -91.045 ;
        RECT -127.195 -91.550 -127.025 -91.225 ;
        RECT -128.095 -91.720 -127.025 -91.550 ;
        RECT -124.055 -91.550 -123.885 -91.225 ;
        RECT -123.705 -91.325 -123.335 -90.985 ;
        RECT -123.155 -91.225 -122.605 -91.055 ;
        RECT -118.555 -91.225 -118.005 -91.055 ;
        RECT -123.155 -91.550 -122.985 -91.225 ;
        RECT -124.055 -91.720 -122.985 -91.550 ;
        RECT -118.175 -91.550 -118.005 -91.225 ;
        RECT -117.825 -91.325 -117.455 -90.985 ;
        RECT -117.275 -91.225 -116.345 -91.045 ;
        RECT -114.895 -91.225 -113.965 -91.045 ;
        RECT -117.275 -91.550 -117.105 -91.225 ;
        RECT -118.175 -91.720 -117.105 -91.550 ;
        RECT -114.135 -91.550 -113.965 -91.225 ;
        RECT -113.785 -91.325 -113.415 -90.985 ;
        RECT -113.235 -91.225 -112.685 -91.055 ;
        RECT -108.635 -91.225 -108.085 -91.055 ;
        RECT -113.235 -91.550 -113.065 -91.225 ;
        RECT -114.135 -91.720 -113.065 -91.550 ;
        RECT -108.255 -91.550 -108.085 -91.225 ;
        RECT -107.905 -91.325 -107.535 -90.985 ;
        RECT -107.355 -91.225 -106.425 -91.045 ;
        RECT -104.975 -91.225 -104.045 -91.045 ;
        RECT -107.355 -91.550 -107.185 -91.225 ;
        RECT -108.255 -91.720 -107.185 -91.550 ;
        RECT -104.215 -91.550 -104.045 -91.225 ;
        RECT -103.865 -91.325 -103.495 -90.985 ;
        RECT -103.315 -91.225 -102.765 -91.055 ;
        RECT -98.715 -91.225 -98.165 -91.055 ;
        RECT -103.315 -91.550 -103.145 -91.225 ;
        RECT -104.215 -91.720 -103.145 -91.550 ;
        RECT -98.335 -91.550 -98.165 -91.225 ;
        RECT -97.985 -91.325 -97.615 -90.985 ;
        RECT -97.435 -91.225 -96.505 -91.045 ;
        RECT -95.055 -91.225 -94.125 -91.045 ;
        RECT -97.435 -91.550 -97.265 -91.225 ;
        RECT -98.335 -91.720 -97.265 -91.550 ;
        RECT -94.295 -91.550 -94.125 -91.225 ;
        RECT -93.945 -91.325 -93.575 -90.985 ;
        RECT -93.395 -91.225 -92.845 -91.055 ;
        RECT -88.795 -91.225 -88.245 -91.055 ;
        RECT -93.395 -91.550 -93.225 -91.225 ;
        RECT -94.295 -91.720 -93.225 -91.550 ;
        RECT -88.415 -91.550 -88.245 -91.225 ;
        RECT -88.065 -91.325 -87.695 -90.985 ;
        RECT -87.515 -91.225 -86.585 -91.045 ;
        RECT -85.135 -91.225 -84.205 -91.045 ;
        RECT -87.515 -91.550 -87.345 -91.225 ;
        RECT -88.415 -91.720 -87.345 -91.550 ;
        RECT -84.375 -91.550 -84.205 -91.225 ;
        RECT -84.025 -91.325 -83.655 -90.985 ;
        RECT -83.475 -91.225 -82.925 -91.055 ;
        RECT -78.875 -91.225 -78.325 -91.055 ;
        RECT -83.475 -91.550 -83.305 -91.225 ;
        RECT -84.375 -91.720 -83.305 -91.550 ;
        RECT -78.495 -91.550 -78.325 -91.225 ;
        RECT -78.145 -91.325 -77.775 -90.985 ;
        RECT -77.595 -91.225 -76.665 -91.045 ;
        RECT -75.215 -91.225 -74.285 -91.045 ;
        RECT -77.595 -91.550 -77.425 -91.225 ;
        RECT -78.495 -91.720 -77.425 -91.550 ;
        RECT -74.455 -91.550 -74.285 -91.225 ;
        RECT -74.105 -91.325 -73.735 -90.985 ;
        RECT -73.555 -91.225 -73.005 -91.055 ;
        RECT -68.955 -91.225 -68.405 -91.055 ;
        RECT -73.555 -91.550 -73.385 -91.225 ;
        RECT -74.455 -91.720 -73.385 -91.550 ;
        RECT -68.575 -91.550 -68.405 -91.225 ;
        RECT -68.225 -91.325 -67.855 -90.985 ;
        RECT -67.675 -91.225 -66.745 -91.045 ;
        RECT -65.295 -91.225 -64.365 -91.045 ;
        RECT -67.675 -91.550 -67.505 -91.225 ;
        RECT -68.575 -91.720 -67.505 -91.550 ;
        RECT -64.535 -91.550 -64.365 -91.225 ;
        RECT -64.185 -91.325 -63.815 -90.985 ;
        RECT -63.635 -91.225 -63.085 -91.055 ;
        RECT -59.035 -91.225 -58.485 -91.055 ;
        RECT -63.635 -91.550 -63.465 -91.225 ;
        RECT -64.535 -91.720 -63.465 -91.550 ;
        RECT -58.655 -91.550 -58.485 -91.225 ;
        RECT -58.305 -91.325 -57.935 -90.985 ;
        RECT -57.755 -91.225 -56.825 -91.045 ;
        RECT -55.375 -91.225 -54.445 -91.045 ;
        RECT -57.755 -91.550 -57.585 -91.225 ;
        RECT -58.655 -91.720 -57.585 -91.550 ;
        RECT -54.615 -91.550 -54.445 -91.225 ;
        RECT -54.265 -91.325 -53.895 -90.985 ;
        RECT -53.715 -91.225 -53.165 -91.055 ;
        RECT -49.115 -91.225 -48.565 -91.055 ;
        RECT -53.715 -91.550 -53.545 -91.225 ;
        RECT -54.615 -91.720 -53.545 -91.550 ;
        RECT -48.735 -91.550 -48.565 -91.225 ;
        RECT -48.385 -91.325 -48.015 -90.985 ;
        RECT -47.835 -91.225 -46.905 -91.045 ;
        RECT -45.455 -91.225 -44.525 -91.045 ;
        RECT -47.835 -91.550 -47.665 -91.225 ;
        RECT -48.735 -91.720 -47.665 -91.550 ;
        RECT -44.695 -91.550 -44.525 -91.225 ;
        RECT -44.345 -91.325 -43.975 -90.985 ;
        RECT -43.795 -91.225 -43.245 -91.055 ;
        RECT -39.195 -91.225 -38.645 -91.055 ;
        RECT -43.795 -91.550 -43.625 -91.225 ;
        RECT -44.695 -91.720 -43.625 -91.550 ;
        RECT -38.815 -91.550 -38.645 -91.225 ;
        RECT -38.465 -91.325 -38.095 -90.985 ;
        RECT -37.915 -91.225 -36.985 -91.045 ;
        RECT -35.535 -91.225 -34.605 -91.045 ;
        RECT -37.915 -91.550 -37.745 -91.225 ;
        RECT -38.815 -91.720 -37.745 -91.550 ;
        RECT -34.775 -91.550 -34.605 -91.225 ;
        RECT -34.425 -91.325 -34.055 -90.985 ;
        RECT -33.875 -91.225 -33.325 -91.055 ;
        RECT -29.275 -91.225 -28.725 -91.055 ;
        RECT -33.875 -91.550 -33.705 -91.225 ;
        RECT -34.775 -91.720 -33.705 -91.550 ;
        RECT -28.895 -91.550 -28.725 -91.225 ;
        RECT -28.545 -91.325 -28.175 -90.985 ;
        RECT -27.995 -91.225 -27.065 -91.045 ;
        RECT -25.615 -91.225 -24.685 -91.045 ;
        RECT -27.995 -91.550 -27.825 -91.225 ;
        RECT -28.895 -91.720 -27.825 -91.550 ;
        RECT -24.855 -91.550 -24.685 -91.225 ;
        RECT -24.505 -91.325 -24.135 -90.985 ;
        RECT -23.955 -91.225 -23.405 -91.055 ;
        RECT -19.355 -91.225 -18.805 -91.055 ;
        RECT -23.955 -91.550 -23.785 -91.225 ;
        RECT -24.855 -91.720 -23.785 -91.550 ;
        RECT -18.975 -91.550 -18.805 -91.225 ;
        RECT -18.625 -91.325 -18.255 -90.985 ;
        RECT -18.075 -91.225 -17.145 -91.045 ;
        RECT -15.695 -91.225 -14.765 -91.045 ;
        RECT -18.075 -91.550 -17.905 -91.225 ;
        RECT -18.975 -91.720 -17.905 -91.550 ;
        RECT -14.935 -91.550 -14.765 -91.225 ;
        RECT -14.585 -91.325 -14.215 -90.985 ;
        RECT -14.035 -91.225 -13.485 -91.055 ;
        RECT -9.435 -91.225 -8.885 -91.055 ;
        RECT -14.035 -91.550 -13.865 -91.225 ;
        RECT -14.935 -91.720 -13.865 -91.550 ;
        RECT -9.055 -91.550 -8.885 -91.225 ;
        RECT -8.705 -91.325 -8.335 -90.985 ;
        RECT -8.155 -91.225 -7.225 -91.045 ;
        RECT -5.775 -91.225 -4.845 -91.045 ;
        RECT -8.155 -91.550 -7.985 -91.225 ;
        RECT -9.055 -91.720 -7.985 -91.550 ;
        RECT -5.015 -91.550 -4.845 -91.225 ;
        RECT -4.665 -91.325 -4.295 -90.985 ;
        RECT -4.115 -91.225 -3.565 -91.055 ;
        RECT 0.485 -91.225 1.035 -91.055 ;
        RECT -4.115 -91.550 -3.945 -91.225 ;
        RECT -5.015 -91.720 -3.945 -91.550 ;
        RECT 0.865 -91.550 1.035 -91.225 ;
        RECT 1.215 -91.325 1.585 -90.985 ;
        RECT 1.765 -91.225 2.695 -91.045 ;
        RECT 4.145 -91.225 5.075 -91.045 ;
        RECT 1.765 -91.550 1.935 -91.225 ;
        RECT 0.865 -91.720 1.935 -91.550 ;
        RECT 4.905 -91.550 5.075 -91.225 ;
        RECT 5.255 -91.325 5.625 -90.985 ;
        RECT 5.805 -91.225 6.355 -91.055 ;
        RECT 10.405 -91.225 10.955 -91.055 ;
        RECT 5.805 -91.550 5.975 -91.225 ;
        RECT 4.905 -91.720 5.975 -91.550 ;
        RECT 10.785 -91.550 10.955 -91.225 ;
        RECT 11.135 -91.325 11.505 -90.985 ;
        RECT 11.685 -91.225 12.615 -91.045 ;
        RECT 14.065 -91.225 14.995 -91.045 ;
        RECT 11.685 -91.550 11.855 -91.225 ;
        RECT 10.785 -91.720 11.855 -91.550 ;
        RECT 14.825 -91.550 14.995 -91.225 ;
        RECT 15.175 -91.325 15.545 -90.985 ;
        RECT 15.725 -91.225 16.275 -91.055 ;
        RECT 20.325 -91.225 20.875 -91.055 ;
        RECT 15.725 -91.550 15.895 -91.225 ;
        RECT 14.825 -91.720 15.895 -91.550 ;
        RECT 20.705 -91.550 20.875 -91.225 ;
        RECT 21.055 -91.325 21.425 -90.985 ;
        RECT 21.605 -91.225 22.535 -91.045 ;
        RECT 23.985 -91.225 24.915 -91.045 ;
        RECT 21.605 -91.550 21.775 -91.225 ;
        RECT 20.705 -91.720 21.775 -91.550 ;
        RECT 24.745 -91.550 24.915 -91.225 ;
        RECT 25.095 -91.325 25.465 -90.985 ;
        RECT 25.645 -91.225 26.195 -91.055 ;
        RECT 25.645 -91.550 25.815 -91.225 ;
        RECT 26.365 -91.405 26.535 -90.880 ;
        RECT 24.745 -91.720 25.815 -91.550 ;
        RECT -287.535 -91.920 -287.365 -91.735 ;
        RECT -286.390 -91.825 -286.060 -91.720 ;
        RECT -282.460 -91.825 -282.130 -91.720 ;
        RECT -276.470 -91.825 -276.140 -91.720 ;
        RECT -272.540 -91.825 -272.210 -91.720 ;
        RECT -266.550 -91.825 -266.220 -91.720 ;
        RECT -262.620 -91.825 -262.290 -91.720 ;
        RECT -256.630 -91.825 -256.300 -91.720 ;
        RECT -252.700 -91.825 -252.370 -91.720 ;
        RECT -246.710 -91.825 -246.380 -91.720 ;
        RECT -242.780 -91.825 -242.450 -91.720 ;
        RECT -236.790 -91.825 -236.460 -91.720 ;
        RECT -232.860 -91.825 -232.530 -91.720 ;
        RECT -226.870 -91.825 -226.540 -91.720 ;
        RECT -222.940 -91.825 -222.610 -91.720 ;
        RECT -216.950 -91.825 -216.620 -91.720 ;
        RECT -213.020 -91.825 -212.690 -91.720 ;
        RECT -207.030 -91.825 -206.700 -91.720 ;
        RECT -203.100 -91.825 -202.770 -91.720 ;
        RECT -197.110 -91.825 -196.780 -91.720 ;
        RECT -193.180 -91.825 -192.850 -91.720 ;
        RECT -187.190 -91.825 -186.860 -91.720 ;
        RECT -183.260 -91.825 -182.930 -91.720 ;
        RECT -177.270 -91.825 -176.940 -91.720 ;
        RECT -173.340 -91.825 -173.010 -91.720 ;
        RECT -167.350 -91.825 -167.020 -91.720 ;
        RECT -163.420 -91.825 -163.090 -91.720 ;
        RECT -157.430 -91.825 -157.100 -91.720 ;
        RECT -153.500 -91.825 -153.170 -91.720 ;
        RECT -147.510 -91.825 -147.180 -91.720 ;
        RECT -143.580 -91.825 -143.250 -91.720 ;
        RECT -137.590 -91.825 -137.260 -91.720 ;
        RECT -133.660 -91.825 -133.330 -91.720 ;
        RECT -127.670 -91.825 -127.340 -91.720 ;
        RECT -123.740 -91.825 -123.410 -91.720 ;
        RECT -117.750 -91.825 -117.420 -91.720 ;
        RECT -113.820 -91.825 -113.490 -91.720 ;
        RECT -107.830 -91.825 -107.500 -91.720 ;
        RECT -103.900 -91.825 -103.570 -91.720 ;
        RECT -97.910 -91.825 -97.580 -91.720 ;
        RECT -93.980 -91.825 -93.650 -91.720 ;
        RECT -87.990 -91.825 -87.660 -91.720 ;
        RECT -84.060 -91.825 -83.730 -91.720 ;
        RECT -78.070 -91.825 -77.740 -91.720 ;
        RECT -74.140 -91.825 -73.810 -91.720 ;
        RECT -68.150 -91.825 -67.820 -91.720 ;
        RECT -64.220 -91.825 -63.890 -91.720 ;
        RECT -58.230 -91.825 -57.900 -91.720 ;
        RECT -54.300 -91.825 -53.970 -91.720 ;
        RECT -48.310 -91.825 -47.980 -91.720 ;
        RECT -44.380 -91.825 -44.050 -91.720 ;
        RECT -38.390 -91.825 -38.060 -91.720 ;
        RECT -34.460 -91.825 -34.130 -91.720 ;
        RECT -28.470 -91.825 -28.140 -91.720 ;
        RECT -24.540 -91.825 -24.210 -91.720 ;
        RECT -18.550 -91.825 -18.220 -91.720 ;
        RECT -14.620 -91.825 -14.290 -91.720 ;
        RECT -8.630 -91.825 -8.300 -91.720 ;
        RECT -4.700 -91.825 -4.370 -91.720 ;
        RECT 1.290 -91.825 1.620 -91.720 ;
        RECT 5.220 -91.825 5.550 -91.720 ;
        RECT 11.210 -91.825 11.540 -91.720 ;
        RECT 15.140 -91.825 15.470 -91.720 ;
        RECT 21.130 -91.825 21.460 -91.720 ;
        RECT 25.060 -91.825 25.390 -91.720 ;
        RECT 25.985 -91.735 26.535 -91.405 ;
        RECT -288.065 -91.935 -287.365 -91.920 ;
        RECT -288.150 -92.105 -287.365 -91.935 ;
        RECT -287.830 -92.110 -287.365 -92.105 ;
        RECT -287.535 -92.260 -287.365 -92.110 ;
        RECT -283.535 -91.995 -282.630 -91.905 ;
        RECT -281.830 -91.995 -281.325 -91.915 ;
        RECT -283.535 -92.175 -281.325 -91.995 ;
        RECT -273.615 -91.995 -272.710 -91.905 ;
        RECT -271.910 -91.995 -271.405 -91.915 ;
        RECT -273.615 -92.175 -271.405 -91.995 ;
        RECT -263.695 -91.995 -262.790 -91.905 ;
        RECT -261.990 -91.995 -261.485 -91.915 ;
        RECT -263.695 -92.175 -261.485 -91.995 ;
        RECT -253.775 -91.995 -252.870 -91.905 ;
        RECT -252.070 -91.995 -251.565 -91.915 ;
        RECT -253.775 -92.175 -251.565 -91.995 ;
        RECT -243.855 -91.995 -242.950 -91.905 ;
        RECT -242.150 -91.995 -241.645 -91.915 ;
        RECT -243.855 -92.175 -241.645 -91.995 ;
        RECT -233.935 -91.995 -233.030 -91.905 ;
        RECT -232.230 -91.995 -231.725 -91.915 ;
        RECT -233.935 -92.175 -231.725 -91.995 ;
        RECT -224.015 -91.995 -223.110 -91.905 ;
        RECT -222.310 -91.995 -221.805 -91.915 ;
        RECT -224.015 -92.175 -221.805 -91.995 ;
        RECT -214.095 -91.995 -213.190 -91.905 ;
        RECT -212.390 -91.995 -211.885 -91.915 ;
        RECT -214.095 -92.175 -211.885 -91.995 ;
        RECT -204.175 -91.995 -203.270 -91.905 ;
        RECT -202.470 -91.995 -201.965 -91.915 ;
        RECT -204.175 -92.175 -201.965 -91.995 ;
        RECT -194.255 -91.995 -193.350 -91.905 ;
        RECT -192.550 -91.995 -192.045 -91.915 ;
        RECT -194.255 -92.175 -192.045 -91.995 ;
        RECT -184.335 -91.995 -183.430 -91.905 ;
        RECT -182.630 -91.995 -182.125 -91.915 ;
        RECT -184.335 -92.175 -182.125 -91.995 ;
        RECT -174.415 -91.995 -173.510 -91.905 ;
        RECT -172.710 -91.995 -172.205 -91.915 ;
        RECT -174.415 -92.175 -172.205 -91.995 ;
        RECT -164.495 -91.995 -163.590 -91.905 ;
        RECT -162.790 -91.995 -162.285 -91.915 ;
        RECT -164.495 -92.175 -162.285 -91.995 ;
        RECT -154.575 -91.995 -153.670 -91.905 ;
        RECT -152.870 -91.995 -152.365 -91.915 ;
        RECT -154.575 -92.175 -152.365 -91.995 ;
        RECT -144.655 -91.995 -143.750 -91.905 ;
        RECT -142.950 -91.995 -142.445 -91.915 ;
        RECT -144.655 -92.175 -142.445 -91.995 ;
        RECT -134.735 -91.995 -133.830 -91.905 ;
        RECT -133.030 -91.995 -132.525 -91.915 ;
        RECT -134.735 -92.175 -132.525 -91.995 ;
        RECT -124.815 -91.995 -123.910 -91.905 ;
        RECT -123.110 -91.995 -122.605 -91.915 ;
        RECT -124.815 -92.175 -122.605 -91.995 ;
        RECT -114.895 -91.995 -113.990 -91.905 ;
        RECT -113.190 -91.995 -112.685 -91.915 ;
        RECT -114.895 -92.175 -112.685 -91.995 ;
        RECT -104.975 -91.995 -104.070 -91.905 ;
        RECT -103.270 -91.995 -102.765 -91.915 ;
        RECT -104.975 -92.175 -102.765 -91.995 ;
        RECT -95.055 -91.995 -94.150 -91.905 ;
        RECT -93.350 -91.995 -92.845 -91.915 ;
        RECT -95.055 -92.175 -92.845 -91.995 ;
        RECT -85.135 -91.995 -84.230 -91.905 ;
        RECT -83.430 -91.995 -82.925 -91.915 ;
        RECT -85.135 -92.175 -82.925 -91.995 ;
        RECT -75.215 -91.995 -74.310 -91.905 ;
        RECT -73.510 -91.995 -73.005 -91.915 ;
        RECT -75.215 -92.175 -73.005 -91.995 ;
        RECT -65.295 -91.995 -64.390 -91.905 ;
        RECT -63.590 -91.995 -63.085 -91.915 ;
        RECT -65.295 -92.175 -63.085 -91.995 ;
        RECT -55.375 -91.995 -54.470 -91.905 ;
        RECT -53.670 -91.995 -53.165 -91.915 ;
        RECT -55.375 -92.175 -53.165 -91.995 ;
        RECT -45.455 -91.995 -44.550 -91.905 ;
        RECT -43.750 -91.995 -43.245 -91.915 ;
        RECT -45.455 -92.175 -43.245 -91.995 ;
        RECT -35.535 -91.995 -34.630 -91.905 ;
        RECT -33.830 -91.995 -33.325 -91.915 ;
        RECT -35.535 -92.175 -33.325 -91.995 ;
        RECT -25.615 -91.995 -24.710 -91.905 ;
        RECT -23.910 -91.995 -23.405 -91.915 ;
        RECT -25.615 -92.175 -23.405 -91.995 ;
        RECT -15.695 -91.995 -14.790 -91.905 ;
        RECT -13.990 -91.995 -13.485 -91.915 ;
        RECT -15.695 -92.175 -13.485 -91.995 ;
        RECT -5.775 -91.995 -4.870 -91.905 ;
        RECT -4.070 -91.995 -3.565 -91.915 ;
        RECT -5.775 -92.175 -3.565 -91.995 ;
        RECT 4.145 -91.995 5.050 -91.905 ;
        RECT 5.850 -91.995 6.355 -91.915 ;
        RECT 4.145 -92.175 6.355 -91.995 ;
        RECT 14.065 -91.995 14.970 -91.905 ;
        RECT 15.770 -91.995 16.275 -91.915 ;
        RECT 14.065 -92.175 16.275 -91.995 ;
        RECT 23.985 -91.995 24.890 -91.905 ;
        RECT 25.690 -91.995 26.195 -91.915 ;
        RECT 23.985 -92.175 26.195 -91.995 ;
        RECT 26.365 -91.930 26.535 -91.735 ;
        RECT 26.775 -91.930 27.065 -91.210 ;
        RECT 26.365 -91.935 27.065 -91.930 ;
        RECT 26.365 -92.105 27.150 -91.935 ;
        RECT 26.365 -92.110 26.830 -92.105 ;
        RECT 26.365 -92.260 26.535 -92.110 ;
        RECT -288.585 -173.780 -288.415 -173.630 ;
        RECT -289.200 -173.950 -288.415 -173.780 ;
        RECT -289.115 -175.115 -288.825 -173.950 ;
        RECT -288.585 -174.155 -288.415 -173.950 ;
        RECT -288.245 -173.895 -286.035 -173.715 ;
        RECT -288.245 -173.985 -287.340 -173.895 ;
        RECT -286.540 -173.975 -286.035 -173.895 ;
        RECT -278.325 -173.895 -276.115 -173.715 ;
        RECT -278.325 -173.985 -277.420 -173.895 ;
        RECT -276.620 -173.975 -276.115 -173.895 ;
        RECT -268.405 -173.895 -266.195 -173.715 ;
        RECT -268.405 -173.985 -267.500 -173.895 ;
        RECT -266.700 -173.975 -266.195 -173.895 ;
        RECT -258.485 -173.895 -256.275 -173.715 ;
        RECT -258.485 -173.985 -257.580 -173.895 ;
        RECT -256.780 -173.975 -256.275 -173.895 ;
        RECT -248.565 -173.895 -246.355 -173.715 ;
        RECT -248.565 -173.985 -247.660 -173.895 ;
        RECT -246.860 -173.975 -246.355 -173.895 ;
        RECT -238.645 -173.895 -236.435 -173.715 ;
        RECT -238.645 -173.985 -237.740 -173.895 ;
        RECT -236.940 -173.975 -236.435 -173.895 ;
        RECT -228.725 -173.895 -226.515 -173.715 ;
        RECT -228.725 -173.985 -227.820 -173.895 ;
        RECT -227.020 -173.975 -226.515 -173.895 ;
        RECT -218.805 -173.895 -216.595 -173.715 ;
        RECT -218.805 -173.985 -217.900 -173.895 ;
        RECT -217.100 -173.975 -216.595 -173.895 ;
        RECT -208.885 -173.895 -206.675 -173.715 ;
        RECT -208.885 -173.985 -207.980 -173.895 ;
        RECT -207.180 -173.975 -206.675 -173.895 ;
        RECT -198.965 -173.895 -196.755 -173.715 ;
        RECT -198.965 -173.985 -198.060 -173.895 ;
        RECT -197.260 -173.975 -196.755 -173.895 ;
        RECT -189.045 -173.895 -186.835 -173.715 ;
        RECT -189.045 -173.985 -188.140 -173.895 ;
        RECT -187.340 -173.975 -186.835 -173.895 ;
        RECT -179.125 -173.895 -176.915 -173.715 ;
        RECT -179.125 -173.985 -178.220 -173.895 ;
        RECT -177.420 -173.975 -176.915 -173.895 ;
        RECT -169.205 -173.895 -166.995 -173.715 ;
        RECT -169.205 -173.985 -168.300 -173.895 ;
        RECT -167.500 -173.975 -166.995 -173.895 ;
        RECT -159.285 -173.895 -157.075 -173.715 ;
        RECT -159.285 -173.985 -158.380 -173.895 ;
        RECT -157.580 -173.975 -157.075 -173.895 ;
        RECT -149.365 -173.895 -147.155 -173.715 ;
        RECT -149.365 -173.985 -148.460 -173.895 ;
        RECT -147.660 -173.975 -147.155 -173.895 ;
        RECT -139.445 -173.895 -137.235 -173.715 ;
        RECT -139.445 -173.985 -138.540 -173.895 ;
        RECT -137.740 -173.975 -137.235 -173.895 ;
        RECT -129.525 -173.895 -127.315 -173.715 ;
        RECT -129.525 -173.985 -128.620 -173.895 ;
        RECT -127.820 -173.975 -127.315 -173.895 ;
        RECT -119.605 -173.895 -117.395 -173.715 ;
        RECT -119.605 -173.985 -118.700 -173.895 ;
        RECT -117.900 -173.975 -117.395 -173.895 ;
        RECT -109.685 -173.895 -107.475 -173.715 ;
        RECT -109.685 -173.985 -108.780 -173.895 ;
        RECT -107.980 -173.975 -107.475 -173.895 ;
        RECT -99.765 -173.895 -97.555 -173.715 ;
        RECT -99.765 -173.985 -98.860 -173.895 ;
        RECT -98.060 -173.975 -97.555 -173.895 ;
        RECT -89.845 -173.895 -87.635 -173.715 ;
        RECT -89.845 -173.985 -88.940 -173.895 ;
        RECT -88.140 -173.975 -87.635 -173.895 ;
        RECT -79.925 -173.895 -77.715 -173.715 ;
        RECT -79.925 -173.985 -79.020 -173.895 ;
        RECT -78.220 -173.975 -77.715 -173.895 ;
        RECT -70.005 -173.895 -67.795 -173.715 ;
        RECT -70.005 -173.985 -69.100 -173.895 ;
        RECT -68.300 -173.975 -67.795 -173.895 ;
        RECT -60.085 -173.895 -57.875 -173.715 ;
        RECT -60.085 -173.985 -59.180 -173.895 ;
        RECT -58.380 -173.975 -57.875 -173.895 ;
        RECT -50.165 -173.895 -47.955 -173.715 ;
        RECT -50.165 -173.985 -49.260 -173.895 ;
        RECT -48.460 -173.975 -47.955 -173.895 ;
        RECT -40.245 -173.895 -38.035 -173.715 ;
        RECT -40.245 -173.985 -39.340 -173.895 ;
        RECT -38.540 -173.975 -38.035 -173.895 ;
        RECT -30.325 -173.895 -28.115 -173.715 ;
        RECT -30.325 -173.985 -29.420 -173.895 ;
        RECT -28.620 -173.975 -28.115 -173.895 ;
        RECT -20.405 -173.895 -18.195 -173.715 ;
        RECT -20.405 -173.985 -19.500 -173.895 ;
        RECT -18.700 -173.975 -18.195 -173.895 ;
        RECT -10.485 -173.895 -8.275 -173.715 ;
        RECT -10.485 -173.985 -9.580 -173.895 ;
        RECT -8.780 -173.975 -8.275 -173.895 ;
        RECT -0.565 -173.895 1.645 -173.715 ;
        RECT -0.565 -173.985 0.340 -173.895 ;
        RECT 1.140 -173.975 1.645 -173.895 ;
        RECT 9.355 -173.895 11.565 -173.715 ;
        RECT 9.355 -173.985 10.260 -173.895 ;
        RECT 11.060 -173.975 11.565 -173.895 ;
        RECT 19.275 -173.895 21.485 -173.715 ;
        RECT 19.275 -173.985 20.180 -173.895 ;
        RECT 20.980 -173.975 21.485 -173.895 ;
        RECT -288.585 -174.485 -287.655 -174.155 ;
        RECT -287.170 -174.170 -286.840 -174.065 ;
        RECT -281.180 -174.170 -280.850 -174.065 ;
        RECT -277.250 -174.170 -276.920 -174.065 ;
        RECT -271.260 -174.170 -270.930 -174.065 ;
        RECT -267.330 -174.170 -267.000 -174.065 ;
        RECT -261.340 -174.170 -261.010 -174.065 ;
        RECT -257.410 -174.170 -257.080 -174.065 ;
        RECT -251.420 -174.170 -251.090 -174.065 ;
        RECT -247.490 -174.170 -247.160 -174.065 ;
        RECT -241.500 -174.170 -241.170 -174.065 ;
        RECT -237.570 -174.170 -237.240 -174.065 ;
        RECT -231.580 -174.170 -231.250 -174.065 ;
        RECT -227.650 -174.170 -227.320 -174.065 ;
        RECT -221.660 -174.170 -221.330 -174.065 ;
        RECT -217.730 -174.170 -217.400 -174.065 ;
        RECT -211.740 -174.170 -211.410 -174.065 ;
        RECT -207.810 -174.170 -207.480 -174.065 ;
        RECT -201.820 -174.170 -201.490 -174.065 ;
        RECT -197.890 -174.170 -197.560 -174.065 ;
        RECT -191.900 -174.170 -191.570 -174.065 ;
        RECT -187.970 -174.170 -187.640 -174.065 ;
        RECT -181.980 -174.170 -181.650 -174.065 ;
        RECT -178.050 -174.170 -177.720 -174.065 ;
        RECT -172.060 -174.170 -171.730 -174.065 ;
        RECT -168.130 -174.170 -167.800 -174.065 ;
        RECT -162.140 -174.170 -161.810 -174.065 ;
        RECT -158.210 -174.170 -157.880 -174.065 ;
        RECT -152.220 -174.170 -151.890 -174.065 ;
        RECT -148.290 -174.170 -147.960 -174.065 ;
        RECT -142.300 -174.170 -141.970 -174.065 ;
        RECT -138.370 -174.170 -138.040 -174.065 ;
        RECT -132.380 -174.170 -132.050 -174.065 ;
        RECT -128.450 -174.170 -128.120 -174.065 ;
        RECT -122.460 -174.170 -122.130 -174.065 ;
        RECT -118.530 -174.170 -118.200 -174.065 ;
        RECT -112.540 -174.170 -112.210 -174.065 ;
        RECT -108.610 -174.170 -108.280 -174.065 ;
        RECT -102.620 -174.170 -102.290 -174.065 ;
        RECT -98.690 -174.170 -98.360 -174.065 ;
        RECT -92.700 -174.170 -92.370 -174.065 ;
        RECT -88.770 -174.170 -88.440 -174.065 ;
        RECT -82.780 -174.170 -82.450 -174.065 ;
        RECT -78.850 -174.170 -78.520 -174.065 ;
        RECT -72.860 -174.170 -72.530 -174.065 ;
        RECT -68.930 -174.170 -68.600 -174.065 ;
        RECT -62.940 -174.170 -62.610 -174.065 ;
        RECT -59.010 -174.170 -58.680 -174.065 ;
        RECT -53.020 -174.170 -52.690 -174.065 ;
        RECT -49.090 -174.170 -48.760 -174.065 ;
        RECT -43.100 -174.170 -42.770 -174.065 ;
        RECT -39.170 -174.170 -38.840 -174.065 ;
        RECT -33.180 -174.170 -32.850 -174.065 ;
        RECT -29.250 -174.170 -28.920 -174.065 ;
        RECT -23.260 -174.170 -22.930 -174.065 ;
        RECT -19.330 -174.170 -19.000 -174.065 ;
        RECT -13.340 -174.170 -13.010 -174.065 ;
        RECT -9.410 -174.170 -9.080 -174.065 ;
        RECT -3.420 -174.170 -3.090 -174.065 ;
        RECT 0.510 -174.170 0.840 -174.065 ;
        RECT 6.500 -174.170 6.830 -174.065 ;
        RECT 10.430 -174.170 10.760 -174.065 ;
        RECT 16.420 -174.170 16.750 -174.065 ;
        RECT 20.350 -174.170 20.680 -174.065 ;
        RECT 26.340 -174.170 26.670 -174.065 ;
        RECT -287.485 -174.340 -286.415 -174.170 ;
        RECT -288.585 -175.010 -288.415 -174.485 ;
        RECT -287.485 -174.665 -287.315 -174.340 ;
        RECT -288.245 -174.845 -287.315 -174.665 ;
        RECT -287.135 -174.905 -286.765 -174.565 ;
        RECT -286.585 -174.665 -286.415 -174.340 ;
        RECT -281.605 -174.340 -280.535 -174.170 ;
        RECT -281.605 -174.665 -281.435 -174.340 ;
        RECT -286.585 -174.835 -286.035 -174.665 ;
        RECT -281.985 -174.835 -281.435 -174.665 ;
        RECT -281.255 -174.905 -280.885 -174.565 ;
        RECT -280.705 -174.665 -280.535 -174.340 ;
        RECT -277.565 -174.340 -276.495 -174.170 ;
        RECT -277.565 -174.665 -277.395 -174.340 ;
        RECT -280.705 -174.845 -279.775 -174.665 ;
        RECT -278.325 -174.845 -277.395 -174.665 ;
        RECT -277.215 -174.905 -276.845 -174.565 ;
        RECT -276.665 -174.665 -276.495 -174.340 ;
        RECT -271.685 -174.340 -270.615 -174.170 ;
        RECT -271.685 -174.665 -271.515 -174.340 ;
        RECT -276.665 -174.835 -276.115 -174.665 ;
        RECT -272.065 -174.835 -271.515 -174.665 ;
        RECT -271.335 -174.905 -270.965 -174.565 ;
        RECT -270.785 -174.665 -270.615 -174.340 ;
        RECT -267.645 -174.340 -266.575 -174.170 ;
        RECT -267.645 -174.665 -267.475 -174.340 ;
        RECT -270.785 -174.845 -269.855 -174.665 ;
        RECT -268.405 -174.845 -267.475 -174.665 ;
        RECT -267.295 -174.905 -266.925 -174.565 ;
        RECT -266.745 -174.665 -266.575 -174.340 ;
        RECT -261.765 -174.340 -260.695 -174.170 ;
        RECT -261.765 -174.665 -261.595 -174.340 ;
        RECT -266.745 -174.835 -266.195 -174.665 ;
        RECT -262.145 -174.835 -261.595 -174.665 ;
        RECT -261.415 -174.905 -261.045 -174.565 ;
        RECT -260.865 -174.665 -260.695 -174.340 ;
        RECT -257.725 -174.340 -256.655 -174.170 ;
        RECT -257.725 -174.665 -257.555 -174.340 ;
        RECT -260.865 -174.845 -259.935 -174.665 ;
        RECT -258.485 -174.845 -257.555 -174.665 ;
        RECT -257.375 -174.905 -257.005 -174.565 ;
        RECT -256.825 -174.665 -256.655 -174.340 ;
        RECT -251.845 -174.340 -250.775 -174.170 ;
        RECT -251.845 -174.665 -251.675 -174.340 ;
        RECT -256.825 -174.835 -256.275 -174.665 ;
        RECT -252.225 -174.835 -251.675 -174.665 ;
        RECT -251.495 -174.905 -251.125 -174.565 ;
        RECT -250.945 -174.665 -250.775 -174.340 ;
        RECT -247.805 -174.340 -246.735 -174.170 ;
        RECT -247.805 -174.665 -247.635 -174.340 ;
        RECT -250.945 -174.845 -250.015 -174.665 ;
        RECT -248.565 -174.845 -247.635 -174.665 ;
        RECT -247.455 -174.905 -247.085 -174.565 ;
        RECT -246.905 -174.665 -246.735 -174.340 ;
        RECT -241.925 -174.340 -240.855 -174.170 ;
        RECT -241.925 -174.665 -241.755 -174.340 ;
        RECT -246.905 -174.835 -246.355 -174.665 ;
        RECT -242.305 -174.835 -241.755 -174.665 ;
        RECT -241.575 -174.905 -241.205 -174.565 ;
        RECT -241.025 -174.665 -240.855 -174.340 ;
        RECT -237.885 -174.340 -236.815 -174.170 ;
        RECT -237.885 -174.665 -237.715 -174.340 ;
        RECT -241.025 -174.845 -240.095 -174.665 ;
        RECT -238.645 -174.845 -237.715 -174.665 ;
        RECT -237.535 -174.905 -237.165 -174.565 ;
        RECT -236.985 -174.665 -236.815 -174.340 ;
        RECT -232.005 -174.340 -230.935 -174.170 ;
        RECT -232.005 -174.665 -231.835 -174.340 ;
        RECT -236.985 -174.835 -236.435 -174.665 ;
        RECT -232.385 -174.835 -231.835 -174.665 ;
        RECT -231.655 -174.905 -231.285 -174.565 ;
        RECT -231.105 -174.665 -230.935 -174.340 ;
        RECT -227.965 -174.340 -226.895 -174.170 ;
        RECT -227.965 -174.665 -227.795 -174.340 ;
        RECT -231.105 -174.845 -230.175 -174.665 ;
        RECT -228.725 -174.845 -227.795 -174.665 ;
        RECT -227.615 -174.905 -227.245 -174.565 ;
        RECT -227.065 -174.665 -226.895 -174.340 ;
        RECT -222.085 -174.340 -221.015 -174.170 ;
        RECT -222.085 -174.665 -221.915 -174.340 ;
        RECT -227.065 -174.835 -226.515 -174.665 ;
        RECT -222.465 -174.835 -221.915 -174.665 ;
        RECT -221.735 -174.905 -221.365 -174.565 ;
        RECT -221.185 -174.665 -221.015 -174.340 ;
        RECT -218.045 -174.340 -216.975 -174.170 ;
        RECT -218.045 -174.665 -217.875 -174.340 ;
        RECT -221.185 -174.845 -220.255 -174.665 ;
        RECT -218.805 -174.845 -217.875 -174.665 ;
        RECT -217.695 -174.905 -217.325 -174.565 ;
        RECT -217.145 -174.665 -216.975 -174.340 ;
        RECT -212.165 -174.340 -211.095 -174.170 ;
        RECT -212.165 -174.665 -211.995 -174.340 ;
        RECT -217.145 -174.835 -216.595 -174.665 ;
        RECT -212.545 -174.835 -211.995 -174.665 ;
        RECT -211.815 -174.905 -211.445 -174.565 ;
        RECT -211.265 -174.665 -211.095 -174.340 ;
        RECT -208.125 -174.340 -207.055 -174.170 ;
        RECT -208.125 -174.665 -207.955 -174.340 ;
        RECT -211.265 -174.845 -210.335 -174.665 ;
        RECT -208.885 -174.845 -207.955 -174.665 ;
        RECT -207.775 -174.905 -207.405 -174.565 ;
        RECT -207.225 -174.665 -207.055 -174.340 ;
        RECT -202.245 -174.340 -201.175 -174.170 ;
        RECT -202.245 -174.665 -202.075 -174.340 ;
        RECT -207.225 -174.835 -206.675 -174.665 ;
        RECT -202.625 -174.835 -202.075 -174.665 ;
        RECT -201.895 -174.905 -201.525 -174.565 ;
        RECT -201.345 -174.665 -201.175 -174.340 ;
        RECT -198.205 -174.340 -197.135 -174.170 ;
        RECT -198.205 -174.665 -198.035 -174.340 ;
        RECT -201.345 -174.845 -200.415 -174.665 ;
        RECT -198.965 -174.845 -198.035 -174.665 ;
        RECT -197.855 -174.905 -197.485 -174.565 ;
        RECT -197.305 -174.665 -197.135 -174.340 ;
        RECT -192.325 -174.340 -191.255 -174.170 ;
        RECT -192.325 -174.665 -192.155 -174.340 ;
        RECT -197.305 -174.835 -196.755 -174.665 ;
        RECT -192.705 -174.835 -192.155 -174.665 ;
        RECT -191.975 -174.905 -191.605 -174.565 ;
        RECT -191.425 -174.665 -191.255 -174.340 ;
        RECT -188.285 -174.340 -187.215 -174.170 ;
        RECT -188.285 -174.665 -188.115 -174.340 ;
        RECT -191.425 -174.845 -190.495 -174.665 ;
        RECT -189.045 -174.845 -188.115 -174.665 ;
        RECT -187.935 -174.905 -187.565 -174.565 ;
        RECT -187.385 -174.665 -187.215 -174.340 ;
        RECT -182.405 -174.340 -181.335 -174.170 ;
        RECT -182.405 -174.665 -182.235 -174.340 ;
        RECT -187.385 -174.835 -186.835 -174.665 ;
        RECT -182.785 -174.835 -182.235 -174.665 ;
        RECT -182.055 -174.905 -181.685 -174.565 ;
        RECT -181.505 -174.665 -181.335 -174.340 ;
        RECT -178.365 -174.340 -177.295 -174.170 ;
        RECT -178.365 -174.665 -178.195 -174.340 ;
        RECT -181.505 -174.845 -180.575 -174.665 ;
        RECT -179.125 -174.845 -178.195 -174.665 ;
        RECT -178.015 -174.905 -177.645 -174.565 ;
        RECT -177.465 -174.665 -177.295 -174.340 ;
        RECT -172.485 -174.340 -171.415 -174.170 ;
        RECT -172.485 -174.665 -172.315 -174.340 ;
        RECT -177.465 -174.835 -176.915 -174.665 ;
        RECT -172.865 -174.835 -172.315 -174.665 ;
        RECT -172.135 -174.905 -171.765 -174.565 ;
        RECT -171.585 -174.665 -171.415 -174.340 ;
        RECT -168.445 -174.340 -167.375 -174.170 ;
        RECT -168.445 -174.665 -168.275 -174.340 ;
        RECT -171.585 -174.845 -170.655 -174.665 ;
        RECT -169.205 -174.845 -168.275 -174.665 ;
        RECT -168.095 -174.905 -167.725 -174.565 ;
        RECT -167.545 -174.665 -167.375 -174.340 ;
        RECT -162.565 -174.340 -161.495 -174.170 ;
        RECT -162.565 -174.665 -162.395 -174.340 ;
        RECT -167.545 -174.835 -166.995 -174.665 ;
        RECT -162.945 -174.835 -162.395 -174.665 ;
        RECT -162.215 -174.905 -161.845 -174.565 ;
        RECT -161.665 -174.665 -161.495 -174.340 ;
        RECT -158.525 -174.340 -157.455 -174.170 ;
        RECT -158.525 -174.665 -158.355 -174.340 ;
        RECT -161.665 -174.845 -160.735 -174.665 ;
        RECT -159.285 -174.845 -158.355 -174.665 ;
        RECT -158.175 -174.905 -157.805 -174.565 ;
        RECT -157.625 -174.665 -157.455 -174.340 ;
        RECT -152.645 -174.340 -151.575 -174.170 ;
        RECT -152.645 -174.665 -152.475 -174.340 ;
        RECT -157.625 -174.835 -157.075 -174.665 ;
        RECT -153.025 -174.835 -152.475 -174.665 ;
        RECT -152.295 -174.905 -151.925 -174.565 ;
        RECT -151.745 -174.665 -151.575 -174.340 ;
        RECT -148.605 -174.340 -147.535 -174.170 ;
        RECT -148.605 -174.665 -148.435 -174.340 ;
        RECT -151.745 -174.845 -150.815 -174.665 ;
        RECT -149.365 -174.845 -148.435 -174.665 ;
        RECT -148.255 -174.905 -147.885 -174.565 ;
        RECT -147.705 -174.665 -147.535 -174.340 ;
        RECT -142.725 -174.340 -141.655 -174.170 ;
        RECT -142.725 -174.665 -142.555 -174.340 ;
        RECT -147.705 -174.835 -147.155 -174.665 ;
        RECT -143.105 -174.835 -142.555 -174.665 ;
        RECT -142.375 -174.905 -142.005 -174.565 ;
        RECT -141.825 -174.665 -141.655 -174.340 ;
        RECT -138.685 -174.340 -137.615 -174.170 ;
        RECT -138.685 -174.665 -138.515 -174.340 ;
        RECT -141.825 -174.845 -140.895 -174.665 ;
        RECT -139.445 -174.845 -138.515 -174.665 ;
        RECT -138.335 -174.905 -137.965 -174.565 ;
        RECT -137.785 -174.665 -137.615 -174.340 ;
        RECT -132.805 -174.340 -131.735 -174.170 ;
        RECT -132.805 -174.665 -132.635 -174.340 ;
        RECT -137.785 -174.835 -137.235 -174.665 ;
        RECT -133.185 -174.835 -132.635 -174.665 ;
        RECT -132.455 -174.905 -132.085 -174.565 ;
        RECT -131.905 -174.665 -131.735 -174.340 ;
        RECT -128.765 -174.340 -127.695 -174.170 ;
        RECT -128.765 -174.665 -128.595 -174.340 ;
        RECT -131.905 -174.845 -130.975 -174.665 ;
        RECT -129.525 -174.845 -128.595 -174.665 ;
        RECT -128.415 -174.905 -128.045 -174.565 ;
        RECT -127.865 -174.665 -127.695 -174.340 ;
        RECT -122.885 -174.340 -121.815 -174.170 ;
        RECT -122.885 -174.665 -122.715 -174.340 ;
        RECT -127.865 -174.835 -127.315 -174.665 ;
        RECT -123.265 -174.835 -122.715 -174.665 ;
        RECT -122.535 -174.905 -122.165 -174.565 ;
        RECT -121.985 -174.665 -121.815 -174.340 ;
        RECT -118.845 -174.340 -117.775 -174.170 ;
        RECT -118.845 -174.665 -118.675 -174.340 ;
        RECT -121.985 -174.845 -121.055 -174.665 ;
        RECT -119.605 -174.845 -118.675 -174.665 ;
        RECT -118.495 -174.905 -118.125 -174.565 ;
        RECT -117.945 -174.665 -117.775 -174.340 ;
        RECT -112.965 -174.340 -111.895 -174.170 ;
        RECT -112.965 -174.665 -112.795 -174.340 ;
        RECT -117.945 -174.835 -117.395 -174.665 ;
        RECT -113.345 -174.835 -112.795 -174.665 ;
        RECT -112.615 -174.905 -112.245 -174.565 ;
        RECT -112.065 -174.665 -111.895 -174.340 ;
        RECT -108.925 -174.340 -107.855 -174.170 ;
        RECT -108.925 -174.665 -108.755 -174.340 ;
        RECT -112.065 -174.845 -111.135 -174.665 ;
        RECT -109.685 -174.845 -108.755 -174.665 ;
        RECT -108.575 -174.905 -108.205 -174.565 ;
        RECT -108.025 -174.665 -107.855 -174.340 ;
        RECT -103.045 -174.340 -101.975 -174.170 ;
        RECT -103.045 -174.665 -102.875 -174.340 ;
        RECT -108.025 -174.835 -107.475 -174.665 ;
        RECT -103.425 -174.835 -102.875 -174.665 ;
        RECT -102.695 -174.905 -102.325 -174.565 ;
        RECT -102.145 -174.665 -101.975 -174.340 ;
        RECT -99.005 -174.340 -97.935 -174.170 ;
        RECT -99.005 -174.665 -98.835 -174.340 ;
        RECT -102.145 -174.845 -101.215 -174.665 ;
        RECT -99.765 -174.845 -98.835 -174.665 ;
        RECT -98.655 -174.905 -98.285 -174.565 ;
        RECT -98.105 -174.665 -97.935 -174.340 ;
        RECT -93.125 -174.340 -92.055 -174.170 ;
        RECT -93.125 -174.665 -92.955 -174.340 ;
        RECT -98.105 -174.835 -97.555 -174.665 ;
        RECT -93.505 -174.835 -92.955 -174.665 ;
        RECT -92.775 -174.905 -92.405 -174.565 ;
        RECT -92.225 -174.665 -92.055 -174.340 ;
        RECT -89.085 -174.340 -88.015 -174.170 ;
        RECT -89.085 -174.665 -88.915 -174.340 ;
        RECT -92.225 -174.845 -91.295 -174.665 ;
        RECT -89.845 -174.845 -88.915 -174.665 ;
        RECT -88.735 -174.905 -88.365 -174.565 ;
        RECT -88.185 -174.665 -88.015 -174.340 ;
        RECT -83.205 -174.340 -82.135 -174.170 ;
        RECT -83.205 -174.665 -83.035 -174.340 ;
        RECT -88.185 -174.835 -87.635 -174.665 ;
        RECT -83.585 -174.835 -83.035 -174.665 ;
        RECT -82.855 -174.905 -82.485 -174.565 ;
        RECT -82.305 -174.665 -82.135 -174.340 ;
        RECT -79.165 -174.340 -78.095 -174.170 ;
        RECT -79.165 -174.665 -78.995 -174.340 ;
        RECT -82.305 -174.845 -81.375 -174.665 ;
        RECT -79.925 -174.845 -78.995 -174.665 ;
        RECT -78.815 -174.905 -78.445 -174.565 ;
        RECT -78.265 -174.665 -78.095 -174.340 ;
        RECT -73.285 -174.340 -72.215 -174.170 ;
        RECT -73.285 -174.665 -73.115 -174.340 ;
        RECT -78.265 -174.835 -77.715 -174.665 ;
        RECT -73.665 -174.835 -73.115 -174.665 ;
        RECT -72.935 -174.905 -72.565 -174.565 ;
        RECT -72.385 -174.665 -72.215 -174.340 ;
        RECT -69.245 -174.340 -68.175 -174.170 ;
        RECT -69.245 -174.665 -69.075 -174.340 ;
        RECT -72.385 -174.845 -71.455 -174.665 ;
        RECT -70.005 -174.845 -69.075 -174.665 ;
        RECT -68.895 -174.905 -68.525 -174.565 ;
        RECT -68.345 -174.665 -68.175 -174.340 ;
        RECT -63.365 -174.340 -62.295 -174.170 ;
        RECT -63.365 -174.665 -63.195 -174.340 ;
        RECT -68.345 -174.835 -67.795 -174.665 ;
        RECT -63.745 -174.835 -63.195 -174.665 ;
        RECT -63.015 -174.905 -62.645 -174.565 ;
        RECT -62.465 -174.665 -62.295 -174.340 ;
        RECT -59.325 -174.340 -58.255 -174.170 ;
        RECT -59.325 -174.665 -59.155 -174.340 ;
        RECT -62.465 -174.845 -61.535 -174.665 ;
        RECT -60.085 -174.845 -59.155 -174.665 ;
        RECT -58.975 -174.905 -58.605 -174.565 ;
        RECT -58.425 -174.665 -58.255 -174.340 ;
        RECT -53.445 -174.340 -52.375 -174.170 ;
        RECT -53.445 -174.665 -53.275 -174.340 ;
        RECT -58.425 -174.835 -57.875 -174.665 ;
        RECT -53.825 -174.835 -53.275 -174.665 ;
        RECT -53.095 -174.905 -52.725 -174.565 ;
        RECT -52.545 -174.665 -52.375 -174.340 ;
        RECT -49.405 -174.340 -48.335 -174.170 ;
        RECT -49.405 -174.665 -49.235 -174.340 ;
        RECT -52.545 -174.845 -51.615 -174.665 ;
        RECT -50.165 -174.845 -49.235 -174.665 ;
        RECT -49.055 -174.905 -48.685 -174.565 ;
        RECT -48.505 -174.665 -48.335 -174.340 ;
        RECT -43.525 -174.340 -42.455 -174.170 ;
        RECT -43.525 -174.665 -43.355 -174.340 ;
        RECT -48.505 -174.835 -47.955 -174.665 ;
        RECT -43.905 -174.835 -43.355 -174.665 ;
        RECT -43.175 -174.905 -42.805 -174.565 ;
        RECT -42.625 -174.665 -42.455 -174.340 ;
        RECT -39.485 -174.340 -38.415 -174.170 ;
        RECT -39.485 -174.665 -39.315 -174.340 ;
        RECT -42.625 -174.845 -41.695 -174.665 ;
        RECT -40.245 -174.845 -39.315 -174.665 ;
        RECT -39.135 -174.905 -38.765 -174.565 ;
        RECT -38.585 -174.665 -38.415 -174.340 ;
        RECT -33.605 -174.340 -32.535 -174.170 ;
        RECT -33.605 -174.665 -33.435 -174.340 ;
        RECT -38.585 -174.835 -38.035 -174.665 ;
        RECT -33.985 -174.835 -33.435 -174.665 ;
        RECT -33.255 -174.905 -32.885 -174.565 ;
        RECT -32.705 -174.665 -32.535 -174.340 ;
        RECT -29.565 -174.340 -28.495 -174.170 ;
        RECT -29.565 -174.665 -29.395 -174.340 ;
        RECT -32.705 -174.845 -31.775 -174.665 ;
        RECT -30.325 -174.845 -29.395 -174.665 ;
        RECT -29.215 -174.905 -28.845 -174.565 ;
        RECT -28.665 -174.665 -28.495 -174.340 ;
        RECT -23.685 -174.340 -22.615 -174.170 ;
        RECT -23.685 -174.665 -23.515 -174.340 ;
        RECT -28.665 -174.835 -28.115 -174.665 ;
        RECT -24.065 -174.835 -23.515 -174.665 ;
        RECT -23.335 -174.905 -22.965 -174.565 ;
        RECT -22.785 -174.665 -22.615 -174.340 ;
        RECT -19.645 -174.340 -18.575 -174.170 ;
        RECT -19.645 -174.665 -19.475 -174.340 ;
        RECT -22.785 -174.845 -21.855 -174.665 ;
        RECT -20.405 -174.845 -19.475 -174.665 ;
        RECT -19.295 -174.905 -18.925 -174.565 ;
        RECT -18.745 -174.665 -18.575 -174.340 ;
        RECT -13.765 -174.340 -12.695 -174.170 ;
        RECT -13.765 -174.665 -13.595 -174.340 ;
        RECT -18.745 -174.835 -18.195 -174.665 ;
        RECT -14.145 -174.835 -13.595 -174.665 ;
        RECT -13.415 -174.905 -13.045 -174.565 ;
        RECT -12.865 -174.665 -12.695 -174.340 ;
        RECT -9.725 -174.340 -8.655 -174.170 ;
        RECT -9.725 -174.665 -9.555 -174.340 ;
        RECT -12.865 -174.845 -11.935 -174.665 ;
        RECT -10.485 -174.845 -9.555 -174.665 ;
        RECT -9.375 -174.905 -9.005 -174.565 ;
        RECT -8.825 -174.665 -8.655 -174.340 ;
        RECT -3.845 -174.340 -2.775 -174.170 ;
        RECT -3.845 -174.665 -3.675 -174.340 ;
        RECT -8.825 -174.835 -8.275 -174.665 ;
        RECT -4.225 -174.835 -3.675 -174.665 ;
        RECT -3.495 -174.905 -3.125 -174.565 ;
        RECT -2.945 -174.665 -2.775 -174.340 ;
        RECT 0.195 -174.340 1.265 -174.170 ;
        RECT 0.195 -174.665 0.365 -174.340 ;
        RECT -2.945 -174.845 -2.015 -174.665 ;
        RECT -0.565 -174.845 0.365 -174.665 ;
        RECT 0.545 -174.905 0.915 -174.565 ;
        RECT 1.095 -174.665 1.265 -174.340 ;
        RECT 6.075 -174.340 7.145 -174.170 ;
        RECT 6.075 -174.665 6.245 -174.340 ;
        RECT 1.095 -174.835 1.645 -174.665 ;
        RECT 5.695 -174.835 6.245 -174.665 ;
        RECT 6.425 -174.905 6.795 -174.565 ;
        RECT 6.975 -174.665 7.145 -174.340 ;
        RECT 10.115 -174.340 11.185 -174.170 ;
        RECT 10.115 -174.665 10.285 -174.340 ;
        RECT 6.975 -174.845 7.905 -174.665 ;
        RECT 9.355 -174.845 10.285 -174.665 ;
        RECT 10.465 -174.905 10.835 -174.565 ;
        RECT 11.015 -174.665 11.185 -174.340 ;
        RECT 15.995 -174.340 17.065 -174.170 ;
        RECT 15.995 -174.665 16.165 -174.340 ;
        RECT 11.015 -174.835 11.565 -174.665 ;
        RECT 15.615 -174.835 16.165 -174.665 ;
        RECT 16.345 -174.905 16.715 -174.565 ;
        RECT 16.895 -174.665 17.065 -174.340 ;
        RECT 20.035 -174.340 21.105 -174.170 ;
        RECT 20.035 -174.665 20.205 -174.340 ;
        RECT 16.895 -174.845 17.825 -174.665 ;
        RECT 19.275 -174.845 20.205 -174.665 ;
        RECT 20.385 -174.905 20.755 -174.565 ;
        RECT 20.935 -174.665 21.105 -174.340 ;
        RECT 25.915 -174.340 26.985 -174.170 ;
        RECT 25.915 -174.665 26.085 -174.340 ;
        RECT 20.935 -174.835 21.485 -174.665 ;
        RECT 25.535 -174.835 26.085 -174.665 ;
        RECT 26.265 -174.905 26.635 -174.565 ;
        RECT 26.815 -174.665 26.985 -174.340 ;
        RECT 26.815 -174.845 27.745 -174.665 ;
        RECT -289.200 -175.525 -287.360 -175.355 ;
        RECT 26.860 -175.525 28.700 -175.355 ;
        RECT -289.115 -176.250 -288.825 -175.525 ;
        RECT -288.655 -176.325 -288.345 -175.525 ;
        RECT -288.140 -176.325 -287.445 -175.695 ;
        RECT -289.115 -178.075 -288.825 -176.910 ;
        RECT -288.140 -176.925 -287.970 -176.325 ;
        RECT -287.800 -176.765 -287.465 -176.515 ;
        RECT -285.105 -176.675 -284.775 -175.695 ;
        RECT -283.245 -176.675 -282.915 -175.695 ;
        RECT -280.575 -176.325 -279.880 -175.695 ;
        RECT -288.655 -178.075 -288.375 -176.935 ;
        RECT -288.205 -177.905 -287.875 -176.925 ;
        RECT -287.705 -178.075 -287.445 -176.935 ;
        RECT -285.515 -177.085 -285.180 -176.835 ;
        RECT -285.010 -177.275 -284.840 -176.675 ;
        RECT -285.535 -177.905 -284.840 -177.275 ;
        RECT -283.180 -177.275 -283.010 -176.675 ;
        RECT -280.555 -176.765 -280.220 -176.515 ;
        RECT -282.840 -177.085 -282.505 -176.835 ;
        RECT -280.050 -176.925 -279.880 -176.325 ;
        RECT -278.220 -176.325 -277.525 -175.695 ;
        RECT -278.220 -176.925 -278.050 -176.325 ;
        RECT -277.880 -176.765 -277.545 -176.515 ;
        RECT -275.185 -176.675 -274.855 -175.695 ;
        RECT -273.325 -176.675 -272.995 -175.695 ;
        RECT -270.655 -176.325 -269.960 -175.695 ;
        RECT -283.180 -177.905 -282.485 -177.275 ;
        RECT -280.145 -177.905 -279.815 -176.925 ;
        RECT -278.285 -177.905 -277.955 -176.925 ;
        RECT -275.595 -177.085 -275.260 -176.835 ;
        RECT -275.090 -177.275 -274.920 -176.675 ;
        RECT -275.615 -177.905 -274.920 -177.275 ;
        RECT -273.260 -177.275 -273.090 -176.675 ;
        RECT -270.635 -176.765 -270.300 -176.515 ;
        RECT -272.920 -177.085 -272.585 -176.835 ;
        RECT -270.130 -176.925 -269.960 -176.325 ;
        RECT -268.300 -176.325 -267.605 -175.695 ;
        RECT -268.300 -176.925 -268.130 -176.325 ;
        RECT -267.960 -176.765 -267.625 -176.515 ;
        RECT -265.265 -176.675 -264.935 -175.695 ;
        RECT -263.405 -176.675 -263.075 -175.695 ;
        RECT -260.735 -176.325 -260.040 -175.695 ;
        RECT -273.260 -177.905 -272.565 -177.275 ;
        RECT -270.225 -177.905 -269.895 -176.925 ;
        RECT -268.365 -177.905 -268.035 -176.925 ;
        RECT -265.675 -177.085 -265.340 -176.835 ;
        RECT -265.170 -177.275 -265.000 -176.675 ;
        RECT -265.695 -177.905 -265.000 -177.275 ;
        RECT -263.340 -177.275 -263.170 -176.675 ;
        RECT -260.715 -176.765 -260.380 -176.515 ;
        RECT -263.000 -177.085 -262.665 -176.835 ;
        RECT -260.210 -176.925 -260.040 -176.325 ;
        RECT -258.380 -176.325 -257.685 -175.695 ;
        RECT -258.380 -176.925 -258.210 -176.325 ;
        RECT -258.040 -176.765 -257.705 -176.515 ;
        RECT -255.345 -176.675 -255.015 -175.695 ;
        RECT -253.485 -176.675 -253.155 -175.695 ;
        RECT -250.815 -176.325 -250.120 -175.695 ;
        RECT -263.340 -177.905 -262.645 -177.275 ;
        RECT -260.305 -177.905 -259.975 -176.925 ;
        RECT -258.445 -177.905 -258.115 -176.925 ;
        RECT -255.755 -177.085 -255.420 -176.835 ;
        RECT -255.250 -177.275 -255.080 -176.675 ;
        RECT -255.775 -177.905 -255.080 -177.275 ;
        RECT -253.420 -177.275 -253.250 -176.675 ;
        RECT -250.795 -176.765 -250.460 -176.515 ;
        RECT -253.080 -177.085 -252.745 -176.835 ;
        RECT -250.290 -176.925 -250.120 -176.325 ;
        RECT -248.460 -176.325 -247.765 -175.695 ;
        RECT -248.460 -176.925 -248.290 -176.325 ;
        RECT -248.120 -176.765 -247.785 -176.515 ;
        RECT -245.425 -176.675 -245.095 -175.695 ;
        RECT -243.565 -176.675 -243.235 -175.695 ;
        RECT -240.895 -176.325 -240.200 -175.695 ;
        RECT -253.420 -177.905 -252.725 -177.275 ;
        RECT -250.385 -177.905 -250.055 -176.925 ;
        RECT -248.525 -177.905 -248.195 -176.925 ;
        RECT -245.835 -177.085 -245.500 -176.835 ;
        RECT -245.330 -177.275 -245.160 -176.675 ;
        RECT -245.855 -177.905 -245.160 -177.275 ;
        RECT -243.500 -177.275 -243.330 -176.675 ;
        RECT -240.875 -176.765 -240.540 -176.515 ;
        RECT -243.160 -177.085 -242.825 -176.835 ;
        RECT -240.370 -176.925 -240.200 -176.325 ;
        RECT -238.540 -176.325 -237.845 -175.695 ;
        RECT -238.540 -176.925 -238.370 -176.325 ;
        RECT -238.200 -176.765 -237.865 -176.515 ;
        RECT -235.505 -176.675 -235.175 -175.695 ;
        RECT -233.645 -176.675 -233.315 -175.695 ;
        RECT -230.975 -176.325 -230.280 -175.695 ;
        RECT -243.500 -177.905 -242.805 -177.275 ;
        RECT -240.465 -177.905 -240.135 -176.925 ;
        RECT -238.605 -177.905 -238.275 -176.925 ;
        RECT -235.915 -177.085 -235.580 -176.835 ;
        RECT -235.410 -177.275 -235.240 -176.675 ;
        RECT -235.935 -177.905 -235.240 -177.275 ;
        RECT -233.580 -177.275 -233.410 -176.675 ;
        RECT -230.955 -176.765 -230.620 -176.515 ;
        RECT -233.240 -177.085 -232.905 -176.835 ;
        RECT -230.450 -176.925 -230.280 -176.325 ;
        RECT -228.620 -176.325 -227.925 -175.695 ;
        RECT -228.620 -176.925 -228.450 -176.325 ;
        RECT -228.280 -176.765 -227.945 -176.515 ;
        RECT -225.585 -176.675 -225.255 -175.695 ;
        RECT -223.725 -176.675 -223.395 -175.695 ;
        RECT -221.055 -176.325 -220.360 -175.695 ;
        RECT -233.580 -177.905 -232.885 -177.275 ;
        RECT -230.545 -177.905 -230.215 -176.925 ;
        RECT -228.685 -177.905 -228.355 -176.925 ;
        RECT -225.995 -177.085 -225.660 -176.835 ;
        RECT -225.490 -177.275 -225.320 -176.675 ;
        RECT -226.015 -177.905 -225.320 -177.275 ;
        RECT -223.660 -177.275 -223.490 -176.675 ;
        RECT -221.035 -176.765 -220.700 -176.515 ;
        RECT -223.320 -177.085 -222.985 -176.835 ;
        RECT -220.530 -176.925 -220.360 -176.325 ;
        RECT -218.700 -176.325 -218.005 -175.695 ;
        RECT -218.700 -176.925 -218.530 -176.325 ;
        RECT -218.360 -176.765 -218.025 -176.515 ;
        RECT -215.665 -176.675 -215.335 -175.695 ;
        RECT -213.805 -176.675 -213.475 -175.695 ;
        RECT -211.135 -176.325 -210.440 -175.695 ;
        RECT -223.660 -177.905 -222.965 -177.275 ;
        RECT -220.625 -177.905 -220.295 -176.925 ;
        RECT -218.765 -177.905 -218.435 -176.925 ;
        RECT -216.075 -177.085 -215.740 -176.835 ;
        RECT -215.570 -177.275 -215.400 -176.675 ;
        RECT -216.095 -177.905 -215.400 -177.275 ;
        RECT -213.740 -177.275 -213.570 -176.675 ;
        RECT -211.115 -176.765 -210.780 -176.515 ;
        RECT -213.400 -177.085 -213.065 -176.835 ;
        RECT -210.610 -176.925 -210.440 -176.325 ;
        RECT -208.780 -176.325 -208.085 -175.695 ;
        RECT -208.780 -176.925 -208.610 -176.325 ;
        RECT -208.440 -176.765 -208.105 -176.515 ;
        RECT -205.745 -176.675 -205.415 -175.695 ;
        RECT -203.885 -176.675 -203.555 -175.695 ;
        RECT -201.215 -176.325 -200.520 -175.695 ;
        RECT -213.740 -177.905 -213.045 -177.275 ;
        RECT -210.705 -177.905 -210.375 -176.925 ;
        RECT -208.845 -177.905 -208.515 -176.925 ;
        RECT -206.155 -177.085 -205.820 -176.835 ;
        RECT -205.650 -177.275 -205.480 -176.675 ;
        RECT -206.175 -177.905 -205.480 -177.275 ;
        RECT -203.820 -177.275 -203.650 -176.675 ;
        RECT -201.195 -176.765 -200.860 -176.515 ;
        RECT -203.480 -177.085 -203.145 -176.835 ;
        RECT -200.690 -176.925 -200.520 -176.325 ;
        RECT -198.860 -176.325 -198.165 -175.695 ;
        RECT -198.860 -176.925 -198.690 -176.325 ;
        RECT -198.520 -176.765 -198.185 -176.515 ;
        RECT -195.825 -176.675 -195.495 -175.695 ;
        RECT -193.965 -176.675 -193.635 -175.695 ;
        RECT -191.295 -176.325 -190.600 -175.695 ;
        RECT -203.820 -177.905 -203.125 -177.275 ;
        RECT -200.785 -177.905 -200.455 -176.925 ;
        RECT -198.925 -177.905 -198.595 -176.925 ;
        RECT -196.235 -177.085 -195.900 -176.835 ;
        RECT -195.730 -177.275 -195.560 -176.675 ;
        RECT -196.255 -177.905 -195.560 -177.275 ;
        RECT -193.900 -177.275 -193.730 -176.675 ;
        RECT -191.275 -176.765 -190.940 -176.515 ;
        RECT -193.560 -177.085 -193.225 -176.835 ;
        RECT -190.770 -176.925 -190.600 -176.325 ;
        RECT -188.940 -176.325 -188.245 -175.695 ;
        RECT -188.940 -176.925 -188.770 -176.325 ;
        RECT -188.600 -176.765 -188.265 -176.515 ;
        RECT -185.905 -176.675 -185.575 -175.695 ;
        RECT -184.045 -176.675 -183.715 -175.695 ;
        RECT -181.375 -176.325 -180.680 -175.695 ;
        RECT -193.900 -177.905 -193.205 -177.275 ;
        RECT -190.865 -177.905 -190.535 -176.925 ;
        RECT -189.005 -177.905 -188.675 -176.925 ;
        RECT -186.315 -177.085 -185.980 -176.835 ;
        RECT -185.810 -177.275 -185.640 -176.675 ;
        RECT -186.335 -177.905 -185.640 -177.275 ;
        RECT -183.980 -177.275 -183.810 -176.675 ;
        RECT -181.355 -176.765 -181.020 -176.515 ;
        RECT -183.640 -177.085 -183.305 -176.835 ;
        RECT -180.850 -176.925 -180.680 -176.325 ;
        RECT -179.020 -176.325 -178.325 -175.695 ;
        RECT -179.020 -176.925 -178.850 -176.325 ;
        RECT -178.680 -176.765 -178.345 -176.515 ;
        RECT -175.985 -176.675 -175.655 -175.695 ;
        RECT -174.125 -176.675 -173.795 -175.695 ;
        RECT -171.455 -176.325 -170.760 -175.695 ;
        RECT -183.980 -177.905 -183.285 -177.275 ;
        RECT -180.945 -177.905 -180.615 -176.925 ;
        RECT -179.085 -177.905 -178.755 -176.925 ;
        RECT -176.395 -177.085 -176.060 -176.835 ;
        RECT -175.890 -177.275 -175.720 -176.675 ;
        RECT -176.415 -177.905 -175.720 -177.275 ;
        RECT -174.060 -177.275 -173.890 -176.675 ;
        RECT -171.435 -176.765 -171.100 -176.515 ;
        RECT -173.720 -177.085 -173.385 -176.835 ;
        RECT -170.930 -176.925 -170.760 -176.325 ;
        RECT -169.100 -176.325 -168.405 -175.695 ;
        RECT -169.100 -176.925 -168.930 -176.325 ;
        RECT -168.760 -176.765 -168.425 -176.515 ;
        RECT -166.065 -176.675 -165.735 -175.695 ;
        RECT -164.205 -176.675 -163.875 -175.695 ;
        RECT -161.535 -176.325 -160.840 -175.695 ;
        RECT -174.060 -177.905 -173.365 -177.275 ;
        RECT -171.025 -177.905 -170.695 -176.925 ;
        RECT -169.165 -177.905 -168.835 -176.925 ;
        RECT -166.475 -177.085 -166.140 -176.835 ;
        RECT -165.970 -177.275 -165.800 -176.675 ;
        RECT -166.495 -177.905 -165.800 -177.275 ;
        RECT -164.140 -177.275 -163.970 -176.675 ;
        RECT -161.515 -176.765 -161.180 -176.515 ;
        RECT -163.800 -177.085 -163.465 -176.835 ;
        RECT -161.010 -176.925 -160.840 -176.325 ;
        RECT -159.180 -176.325 -158.485 -175.695 ;
        RECT -159.180 -176.925 -159.010 -176.325 ;
        RECT -158.840 -176.765 -158.505 -176.515 ;
        RECT -156.145 -176.675 -155.815 -175.695 ;
        RECT -154.285 -176.675 -153.955 -175.695 ;
        RECT -151.615 -176.325 -150.920 -175.695 ;
        RECT -164.140 -177.905 -163.445 -177.275 ;
        RECT -161.105 -177.905 -160.775 -176.925 ;
        RECT -159.245 -177.905 -158.915 -176.925 ;
        RECT -156.555 -177.085 -156.220 -176.835 ;
        RECT -156.050 -177.275 -155.880 -176.675 ;
        RECT -156.575 -177.905 -155.880 -177.275 ;
        RECT -154.220 -177.275 -154.050 -176.675 ;
        RECT -151.595 -176.765 -151.260 -176.515 ;
        RECT -153.880 -177.085 -153.545 -176.835 ;
        RECT -151.090 -176.925 -150.920 -176.325 ;
        RECT -149.260 -176.325 -148.565 -175.695 ;
        RECT -149.260 -176.925 -149.090 -176.325 ;
        RECT -148.920 -176.765 -148.585 -176.515 ;
        RECT -146.225 -176.675 -145.895 -175.695 ;
        RECT -144.365 -176.675 -144.035 -175.695 ;
        RECT -141.695 -176.325 -141.000 -175.695 ;
        RECT -154.220 -177.905 -153.525 -177.275 ;
        RECT -151.185 -177.905 -150.855 -176.925 ;
        RECT -149.325 -177.905 -148.995 -176.925 ;
        RECT -146.635 -177.085 -146.300 -176.835 ;
        RECT -146.130 -177.275 -145.960 -176.675 ;
        RECT -146.655 -177.905 -145.960 -177.275 ;
        RECT -144.300 -177.275 -144.130 -176.675 ;
        RECT -141.675 -176.765 -141.340 -176.515 ;
        RECT -143.960 -177.085 -143.625 -176.835 ;
        RECT -141.170 -176.925 -141.000 -176.325 ;
        RECT -139.340 -176.325 -138.645 -175.695 ;
        RECT -139.340 -176.925 -139.170 -176.325 ;
        RECT -139.000 -176.765 -138.665 -176.515 ;
        RECT -136.305 -176.675 -135.975 -175.695 ;
        RECT -134.445 -176.675 -134.115 -175.695 ;
        RECT -131.775 -176.325 -131.080 -175.695 ;
        RECT -144.300 -177.905 -143.605 -177.275 ;
        RECT -141.265 -177.905 -140.935 -176.925 ;
        RECT -139.405 -177.905 -139.075 -176.925 ;
        RECT -136.715 -177.085 -136.380 -176.835 ;
        RECT -136.210 -177.275 -136.040 -176.675 ;
        RECT -136.735 -177.905 -136.040 -177.275 ;
        RECT -134.380 -177.275 -134.210 -176.675 ;
        RECT -131.755 -176.765 -131.420 -176.515 ;
        RECT -134.040 -177.085 -133.705 -176.835 ;
        RECT -131.250 -176.925 -131.080 -176.325 ;
        RECT -129.420 -176.325 -128.725 -175.695 ;
        RECT -129.420 -176.925 -129.250 -176.325 ;
        RECT -129.080 -176.765 -128.745 -176.515 ;
        RECT -126.385 -176.675 -126.055 -175.695 ;
        RECT -124.525 -176.675 -124.195 -175.695 ;
        RECT -121.855 -176.325 -121.160 -175.695 ;
        RECT -134.380 -177.905 -133.685 -177.275 ;
        RECT -131.345 -177.905 -131.015 -176.925 ;
        RECT -129.485 -177.905 -129.155 -176.925 ;
        RECT -126.795 -177.085 -126.460 -176.835 ;
        RECT -126.290 -177.275 -126.120 -176.675 ;
        RECT -126.815 -177.905 -126.120 -177.275 ;
        RECT -124.460 -177.275 -124.290 -176.675 ;
        RECT -121.835 -176.765 -121.500 -176.515 ;
        RECT -124.120 -177.085 -123.785 -176.835 ;
        RECT -121.330 -176.925 -121.160 -176.325 ;
        RECT -119.500 -176.325 -118.805 -175.695 ;
        RECT -119.500 -176.925 -119.330 -176.325 ;
        RECT -119.160 -176.765 -118.825 -176.515 ;
        RECT -116.465 -176.675 -116.135 -175.695 ;
        RECT -114.605 -176.675 -114.275 -175.695 ;
        RECT -111.935 -176.325 -111.240 -175.695 ;
        RECT -124.460 -177.905 -123.765 -177.275 ;
        RECT -121.425 -177.905 -121.095 -176.925 ;
        RECT -119.565 -177.905 -119.235 -176.925 ;
        RECT -116.875 -177.085 -116.540 -176.835 ;
        RECT -116.370 -177.275 -116.200 -176.675 ;
        RECT -116.895 -177.905 -116.200 -177.275 ;
        RECT -114.540 -177.275 -114.370 -176.675 ;
        RECT -111.915 -176.765 -111.580 -176.515 ;
        RECT -114.200 -177.085 -113.865 -176.835 ;
        RECT -111.410 -176.925 -111.240 -176.325 ;
        RECT -109.580 -176.325 -108.885 -175.695 ;
        RECT -109.580 -176.925 -109.410 -176.325 ;
        RECT -109.240 -176.765 -108.905 -176.515 ;
        RECT -106.545 -176.675 -106.215 -175.695 ;
        RECT -104.685 -176.675 -104.355 -175.695 ;
        RECT -102.015 -176.325 -101.320 -175.695 ;
        RECT -114.540 -177.905 -113.845 -177.275 ;
        RECT -111.505 -177.905 -111.175 -176.925 ;
        RECT -109.645 -177.905 -109.315 -176.925 ;
        RECT -106.955 -177.085 -106.620 -176.835 ;
        RECT -106.450 -177.275 -106.280 -176.675 ;
        RECT -106.975 -177.905 -106.280 -177.275 ;
        RECT -104.620 -177.275 -104.450 -176.675 ;
        RECT -101.995 -176.765 -101.660 -176.515 ;
        RECT -104.280 -177.085 -103.945 -176.835 ;
        RECT -101.490 -176.925 -101.320 -176.325 ;
        RECT -99.660 -176.325 -98.965 -175.695 ;
        RECT -99.660 -176.925 -99.490 -176.325 ;
        RECT -99.320 -176.765 -98.985 -176.515 ;
        RECT -96.625 -176.675 -96.295 -175.695 ;
        RECT -94.765 -176.675 -94.435 -175.695 ;
        RECT -92.095 -176.325 -91.400 -175.695 ;
        RECT -104.620 -177.905 -103.925 -177.275 ;
        RECT -101.585 -177.905 -101.255 -176.925 ;
        RECT -99.725 -177.905 -99.395 -176.925 ;
        RECT -97.035 -177.085 -96.700 -176.835 ;
        RECT -96.530 -177.275 -96.360 -176.675 ;
        RECT -97.055 -177.905 -96.360 -177.275 ;
        RECT -94.700 -177.275 -94.530 -176.675 ;
        RECT -92.075 -176.765 -91.740 -176.515 ;
        RECT -94.360 -177.085 -94.025 -176.835 ;
        RECT -91.570 -176.925 -91.400 -176.325 ;
        RECT -89.740 -176.325 -89.045 -175.695 ;
        RECT -89.740 -176.925 -89.570 -176.325 ;
        RECT -89.400 -176.765 -89.065 -176.515 ;
        RECT -86.705 -176.675 -86.375 -175.695 ;
        RECT -84.845 -176.675 -84.515 -175.695 ;
        RECT -82.175 -176.325 -81.480 -175.695 ;
        RECT -94.700 -177.905 -94.005 -177.275 ;
        RECT -91.665 -177.905 -91.335 -176.925 ;
        RECT -89.805 -177.905 -89.475 -176.925 ;
        RECT -87.115 -177.085 -86.780 -176.835 ;
        RECT -86.610 -177.275 -86.440 -176.675 ;
        RECT -87.135 -177.905 -86.440 -177.275 ;
        RECT -84.780 -177.275 -84.610 -176.675 ;
        RECT -82.155 -176.765 -81.820 -176.515 ;
        RECT -84.440 -177.085 -84.105 -176.835 ;
        RECT -81.650 -176.925 -81.480 -176.325 ;
        RECT -79.820 -176.325 -79.125 -175.695 ;
        RECT -79.820 -176.925 -79.650 -176.325 ;
        RECT -79.480 -176.765 -79.145 -176.515 ;
        RECT -76.785 -176.675 -76.455 -175.695 ;
        RECT -74.925 -176.675 -74.595 -175.695 ;
        RECT -72.255 -176.325 -71.560 -175.695 ;
        RECT -84.780 -177.905 -84.085 -177.275 ;
        RECT -81.745 -177.905 -81.415 -176.925 ;
        RECT -79.885 -177.905 -79.555 -176.925 ;
        RECT -77.195 -177.085 -76.860 -176.835 ;
        RECT -76.690 -177.275 -76.520 -176.675 ;
        RECT -77.215 -177.905 -76.520 -177.275 ;
        RECT -74.860 -177.275 -74.690 -176.675 ;
        RECT -72.235 -176.765 -71.900 -176.515 ;
        RECT -74.520 -177.085 -74.185 -176.835 ;
        RECT -71.730 -176.925 -71.560 -176.325 ;
        RECT -69.900 -176.325 -69.205 -175.695 ;
        RECT -69.900 -176.925 -69.730 -176.325 ;
        RECT -69.560 -176.765 -69.225 -176.515 ;
        RECT -66.865 -176.675 -66.535 -175.695 ;
        RECT -65.005 -176.675 -64.675 -175.695 ;
        RECT -62.335 -176.325 -61.640 -175.695 ;
        RECT -74.860 -177.905 -74.165 -177.275 ;
        RECT -71.825 -177.905 -71.495 -176.925 ;
        RECT -69.965 -177.905 -69.635 -176.925 ;
        RECT -67.275 -177.085 -66.940 -176.835 ;
        RECT -66.770 -177.275 -66.600 -176.675 ;
        RECT -67.295 -177.905 -66.600 -177.275 ;
        RECT -64.940 -177.275 -64.770 -176.675 ;
        RECT -62.315 -176.765 -61.980 -176.515 ;
        RECT -64.600 -177.085 -64.265 -176.835 ;
        RECT -61.810 -176.925 -61.640 -176.325 ;
        RECT -59.980 -176.325 -59.285 -175.695 ;
        RECT -59.980 -176.925 -59.810 -176.325 ;
        RECT -59.640 -176.765 -59.305 -176.515 ;
        RECT -56.945 -176.675 -56.615 -175.695 ;
        RECT -55.085 -176.675 -54.755 -175.695 ;
        RECT -52.415 -176.325 -51.720 -175.695 ;
        RECT -64.940 -177.905 -64.245 -177.275 ;
        RECT -61.905 -177.905 -61.575 -176.925 ;
        RECT -60.045 -177.905 -59.715 -176.925 ;
        RECT -57.355 -177.085 -57.020 -176.835 ;
        RECT -56.850 -177.275 -56.680 -176.675 ;
        RECT -57.375 -177.905 -56.680 -177.275 ;
        RECT -55.020 -177.275 -54.850 -176.675 ;
        RECT -52.395 -176.765 -52.060 -176.515 ;
        RECT -54.680 -177.085 -54.345 -176.835 ;
        RECT -51.890 -176.925 -51.720 -176.325 ;
        RECT -50.060 -176.325 -49.365 -175.695 ;
        RECT -50.060 -176.925 -49.890 -176.325 ;
        RECT -49.720 -176.765 -49.385 -176.515 ;
        RECT -47.025 -176.675 -46.695 -175.695 ;
        RECT -45.165 -176.675 -44.835 -175.695 ;
        RECT -42.495 -176.325 -41.800 -175.695 ;
        RECT -55.020 -177.905 -54.325 -177.275 ;
        RECT -51.985 -177.905 -51.655 -176.925 ;
        RECT -50.125 -177.905 -49.795 -176.925 ;
        RECT -47.435 -177.085 -47.100 -176.835 ;
        RECT -46.930 -177.275 -46.760 -176.675 ;
        RECT -47.455 -177.905 -46.760 -177.275 ;
        RECT -45.100 -177.275 -44.930 -176.675 ;
        RECT -42.475 -176.765 -42.140 -176.515 ;
        RECT -44.760 -177.085 -44.425 -176.835 ;
        RECT -41.970 -176.925 -41.800 -176.325 ;
        RECT -40.140 -176.325 -39.445 -175.695 ;
        RECT -40.140 -176.925 -39.970 -176.325 ;
        RECT -39.800 -176.765 -39.465 -176.515 ;
        RECT -37.105 -176.675 -36.775 -175.695 ;
        RECT -35.245 -176.675 -34.915 -175.695 ;
        RECT -32.575 -176.325 -31.880 -175.695 ;
        RECT -45.100 -177.905 -44.405 -177.275 ;
        RECT -42.065 -177.905 -41.735 -176.925 ;
        RECT -40.205 -177.905 -39.875 -176.925 ;
        RECT -37.515 -177.085 -37.180 -176.835 ;
        RECT -37.010 -177.275 -36.840 -176.675 ;
        RECT -37.535 -177.905 -36.840 -177.275 ;
        RECT -35.180 -177.275 -35.010 -176.675 ;
        RECT -32.555 -176.765 -32.220 -176.515 ;
        RECT -34.840 -177.085 -34.505 -176.835 ;
        RECT -32.050 -176.925 -31.880 -176.325 ;
        RECT -30.220 -176.325 -29.525 -175.695 ;
        RECT -30.220 -176.925 -30.050 -176.325 ;
        RECT -29.880 -176.765 -29.545 -176.515 ;
        RECT -27.185 -176.675 -26.855 -175.695 ;
        RECT -25.325 -176.675 -24.995 -175.695 ;
        RECT -22.655 -176.325 -21.960 -175.695 ;
        RECT -35.180 -177.905 -34.485 -177.275 ;
        RECT -32.145 -177.905 -31.815 -176.925 ;
        RECT -30.285 -177.905 -29.955 -176.925 ;
        RECT -27.595 -177.085 -27.260 -176.835 ;
        RECT -27.090 -177.275 -26.920 -176.675 ;
        RECT -27.615 -177.905 -26.920 -177.275 ;
        RECT -25.260 -177.275 -25.090 -176.675 ;
        RECT -22.635 -176.765 -22.300 -176.515 ;
        RECT -24.920 -177.085 -24.585 -176.835 ;
        RECT -22.130 -176.925 -21.960 -176.325 ;
        RECT -20.300 -176.325 -19.605 -175.695 ;
        RECT -20.300 -176.925 -20.130 -176.325 ;
        RECT -19.960 -176.765 -19.625 -176.515 ;
        RECT -17.265 -176.675 -16.935 -175.695 ;
        RECT -15.405 -176.675 -15.075 -175.695 ;
        RECT -12.735 -176.325 -12.040 -175.695 ;
        RECT -25.260 -177.905 -24.565 -177.275 ;
        RECT -22.225 -177.905 -21.895 -176.925 ;
        RECT -20.365 -177.905 -20.035 -176.925 ;
        RECT -17.675 -177.085 -17.340 -176.835 ;
        RECT -17.170 -177.275 -17.000 -176.675 ;
        RECT -17.695 -177.905 -17.000 -177.275 ;
        RECT -15.340 -177.275 -15.170 -176.675 ;
        RECT -12.715 -176.765 -12.380 -176.515 ;
        RECT -15.000 -177.085 -14.665 -176.835 ;
        RECT -12.210 -176.925 -12.040 -176.325 ;
        RECT -10.380 -176.325 -9.685 -175.695 ;
        RECT -10.380 -176.925 -10.210 -176.325 ;
        RECT -10.040 -176.765 -9.705 -176.515 ;
        RECT -7.345 -176.675 -7.015 -175.695 ;
        RECT -5.485 -176.675 -5.155 -175.695 ;
        RECT -2.815 -176.325 -2.120 -175.695 ;
        RECT -15.340 -177.905 -14.645 -177.275 ;
        RECT -12.305 -177.905 -11.975 -176.925 ;
        RECT -10.445 -177.905 -10.115 -176.925 ;
        RECT -7.755 -177.085 -7.420 -176.835 ;
        RECT -7.250 -177.275 -7.080 -176.675 ;
        RECT -7.775 -177.905 -7.080 -177.275 ;
        RECT -5.420 -177.275 -5.250 -176.675 ;
        RECT -2.795 -176.765 -2.460 -176.515 ;
        RECT -5.080 -177.085 -4.745 -176.835 ;
        RECT -2.290 -176.925 -2.120 -176.325 ;
        RECT -0.460 -176.325 0.235 -175.695 ;
        RECT -0.460 -176.925 -0.290 -176.325 ;
        RECT -0.120 -176.765 0.215 -176.515 ;
        RECT 2.575 -176.675 2.905 -175.695 ;
        RECT 4.435 -176.675 4.765 -175.695 ;
        RECT 7.105 -176.325 7.800 -175.695 ;
        RECT -5.420 -177.905 -4.725 -177.275 ;
        RECT -2.385 -177.905 -2.055 -176.925 ;
        RECT -0.525 -177.905 -0.195 -176.925 ;
        RECT 2.165 -177.085 2.500 -176.835 ;
        RECT 2.670 -177.275 2.840 -176.675 ;
        RECT 2.145 -177.905 2.840 -177.275 ;
        RECT 4.500 -177.275 4.670 -176.675 ;
        RECT 7.125 -176.765 7.460 -176.515 ;
        RECT 4.840 -177.085 5.175 -176.835 ;
        RECT 7.630 -176.925 7.800 -176.325 ;
        RECT 9.460 -176.325 10.155 -175.695 ;
        RECT 9.460 -176.925 9.630 -176.325 ;
        RECT 9.800 -176.765 10.135 -176.515 ;
        RECT 12.495 -176.675 12.825 -175.695 ;
        RECT 14.355 -176.675 14.685 -175.695 ;
        RECT 17.025 -176.325 17.720 -175.695 ;
        RECT 4.500 -177.905 5.195 -177.275 ;
        RECT 7.535 -177.905 7.865 -176.925 ;
        RECT 9.395 -177.905 9.725 -176.925 ;
        RECT 12.085 -177.085 12.420 -176.835 ;
        RECT 12.590 -177.275 12.760 -176.675 ;
        RECT 12.065 -177.905 12.760 -177.275 ;
        RECT 14.420 -177.275 14.590 -176.675 ;
        RECT 17.045 -176.765 17.380 -176.515 ;
        RECT 14.760 -177.085 15.095 -176.835 ;
        RECT 17.550 -176.925 17.720 -176.325 ;
        RECT 19.380 -176.325 20.075 -175.695 ;
        RECT 19.380 -176.925 19.550 -176.325 ;
        RECT 19.720 -176.765 20.055 -176.515 ;
        RECT 22.415 -176.675 22.745 -175.695 ;
        RECT 24.275 -176.675 24.605 -175.695 ;
        RECT 26.945 -176.325 27.640 -175.695 ;
        RECT 27.845 -176.325 28.155 -175.525 ;
        RECT 28.325 -176.250 28.615 -175.525 ;
        RECT 14.420 -177.905 15.115 -177.275 ;
        RECT 17.455 -177.905 17.785 -176.925 ;
        RECT 19.315 -177.905 19.645 -176.925 ;
        RECT 22.005 -177.085 22.340 -176.835 ;
        RECT 22.510 -177.275 22.680 -176.675 ;
        RECT 21.985 -177.905 22.680 -177.275 ;
        RECT 24.340 -177.275 24.510 -176.675 ;
        RECT 26.965 -176.765 27.300 -176.515 ;
        RECT 24.680 -177.085 25.015 -176.835 ;
        RECT 27.470 -176.925 27.640 -176.325 ;
        RECT 24.340 -177.905 25.035 -177.275 ;
        RECT 27.375 -177.905 27.705 -176.925 ;
        RECT -289.200 -178.245 -287.360 -178.075 ;
        RECT -287.815 -179.630 -287.525 -178.920 ;
        RECT -287.285 -179.115 -287.115 -178.590 ;
        RECT -286.945 -178.935 -286.395 -178.765 ;
        RECT -287.285 -179.445 -286.735 -179.115 ;
        RECT -286.565 -179.260 -286.395 -178.935 ;
        RECT -286.215 -179.035 -285.845 -178.695 ;
        RECT -285.665 -178.935 -284.735 -178.755 ;
        RECT -283.285 -178.935 -282.355 -178.755 ;
        RECT -285.665 -179.260 -285.495 -178.935 ;
        RECT -286.565 -179.430 -285.495 -179.260 ;
        RECT -282.525 -179.260 -282.355 -178.935 ;
        RECT -282.175 -179.035 -281.805 -178.695 ;
        RECT -281.625 -178.935 -281.075 -178.765 ;
        RECT -277.025 -178.935 -276.475 -178.765 ;
        RECT -281.625 -179.260 -281.455 -178.935 ;
        RECT -282.525 -179.430 -281.455 -179.260 ;
        RECT -276.645 -179.260 -276.475 -178.935 ;
        RECT -276.295 -179.035 -275.925 -178.695 ;
        RECT -275.745 -178.935 -274.815 -178.755 ;
        RECT -273.365 -178.935 -272.435 -178.755 ;
        RECT -275.745 -179.260 -275.575 -178.935 ;
        RECT -276.645 -179.430 -275.575 -179.260 ;
        RECT -272.605 -179.260 -272.435 -178.935 ;
        RECT -272.255 -179.035 -271.885 -178.695 ;
        RECT -271.705 -178.935 -271.155 -178.765 ;
        RECT -267.105 -178.935 -266.555 -178.765 ;
        RECT -271.705 -179.260 -271.535 -178.935 ;
        RECT -272.605 -179.430 -271.535 -179.260 ;
        RECT -266.725 -179.260 -266.555 -178.935 ;
        RECT -266.375 -179.035 -266.005 -178.695 ;
        RECT -265.825 -178.935 -264.895 -178.755 ;
        RECT -263.445 -178.935 -262.515 -178.755 ;
        RECT -265.825 -179.260 -265.655 -178.935 ;
        RECT -266.725 -179.430 -265.655 -179.260 ;
        RECT -262.685 -179.260 -262.515 -178.935 ;
        RECT -262.335 -179.035 -261.965 -178.695 ;
        RECT -261.785 -178.935 -261.235 -178.765 ;
        RECT -257.185 -178.935 -256.635 -178.765 ;
        RECT -261.785 -179.260 -261.615 -178.935 ;
        RECT -262.685 -179.430 -261.615 -179.260 ;
        RECT -256.805 -179.260 -256.635 -178.935 ;
        RECT -256.455 -179.035 -256.085 -178.695 ;
        RECT -255.905 -178.935 -254.975 -178.755 ;
        RECT -253.525 -178.935 -252.595 -178.755 ;
        RECT -255.905 -179.260 -255.735 -178.935 ;
        RECT -256.805 -179.430 -255.735 -179.260 ;
        RECT -252.765 -179.260 -252.595 -178.935 ;
        RECT -252.415 -179.035 -252.045 -178.695 ;
        RECT -251.865 -178.935 -251.315 -178.765 ;
        RECT -247.265 -178.935 -246.715 -178.765 ;
        RECT -251.865 -179.260 -251.695 -178.935 ;
        RECT -252.765 -179.430 -251.695 -179.260 ;
        RECT -246.885 -179.260 -246.715 -178.935 ;
        RECT -246.535 -179.035 -246.165 -178.695 ;
        RECT -245.985 -178.935 -245.055 -178.755 ;
        RECT -243.605 -178.935 -242.675 -178.755 ;
        RECT -245.985 -179.260 -245.815 -178.935 ;
        RECT -246.885 -179.430 -245.815 -179.260 ;
        RECT -242.845 -179.260 -242.675 -178.935 ;
        RECT -242.495 -179.035 -242.125 -178.695 ;
        RECT -241.945 -178.935 -241.395 -178.765 ;
        RECT -237.345 -178.935 -236.795 -178.765 ;
        RECT -241.945 -179.260 -241.775 -178.935 ;
        RECT -242.845 -179.430 -241.775 -179.260 ;
        RECT -236.965 -179.260 -236.795 -178.935 ;
        RECT -236.615 -179.035 -236.245 -178.695 ;
        RECT -236.065 -178.935 -235.135 -178.755 ;
        RECT -233.685 -178.935 -232.755 -178.755 ;
        RECT -236.065 -179.260 -235.895 -178.935 ;
        RECT -236.965 -179.430 -235.895 -179.260 ;
        RECT -232.925 -179.260 -232.755 -178.935 ;
        RECT -232.575 -179.035 -232.205 -178.695 ;
        RECT -232.025 -178.935 -231.475 -178.765 ;
        RECT -227.425 -178.935 -226.875 -178.765 ;
        RECT -232.025 -179.260 -231.855 -178.935 ;
        RECT -232.925 -179.430 -231.855 -179.260 ;
        RECT -227.045 -179.260 -226.875 -178.935 ;
        RECT -226.695 -179.035 -226.325 -178.695 ;
        RECT -226.145 -178.935 -225.215 -178.755 ;
        RECT -223.765 -178.935 -222.835 -178.755 ;
        RECT -226.145 -179.260 -225.975 -178.935 ;
        RECT -227.045 -179.430 -225.975 -179.260 ;
        RECT -223.005 -179.260 -222.835 -178.935 ;
        RECT -222.655 -179.035 -222.285 -178.695 ;
        RECT -222.105 -178.935 -221.555 -178.765 ;
        RECT -217.505 -178.935 -216.955 -178.765 ;
        RECT -222.105 -179.260 -221.935 -178.935 ;
        RECT -223.005 -179.430 -221.935 -179.260 ;
        RECT -217.125 -179.260 -216.955 -178.935 ;
        RECT -216.775 -179.035 -216.405 -178.695 ;
        RECT -216.225 -178.935 -215.295 -178.755 ;
        RECT -213.845 -178.935 -212.915 -178.755 ;
        RECT -216.225 -179.260 -216.055 -178.935 ;
        RECT -217.125 -179.430 -216.055 -179.260 ;
        RECT -213.085 -179.260 -212.915 -178.935 ;
        RECT -212.735 -179.035 -212.365 -178.695 ;
        RECT -212.185 -178.935 -211.635 -178.765 ;
        RECT -207.585 -178.935 -207.035 -178.765 ;
        RECT -212.185 -179.260 -212.015 -178.935 ;
        RECT -213.085 -179.430 -212.015 -179.260 ;
        RECT -207.205 -179.260 -207.035 -178.935 ;
        RECT -206.855 -179.035 -206.485 -178.695 ;
        RECT -206.305 -178.935 -205.375 -178.755 ;
        RECT -203.925 -178.935 -202.995 -178.755 ;
        RECT -206.305 -179.260 -206.135 -178.935 ;
        RECT -207.205 -179.430 -206.135 -179.260 ;
        RECT -203.165 -179.260 -202.995 -178.935 ;
        RECT -202.815 -179.035 -202.445 -178.695 ;
        RECT -202.265 -178.935 -201.715 -178.765 ;
        RECT -197.665 -178.935 -197.115 -178.765 ;
        RECT -202.265 -179.260 -202.095 -178.935 ;
        RECT -203.165 -179.430 -202.095 -179.260 ;
        RECT -197.285 -179.260 -197.115 -178.935 ;
        RECT -196.935 -179.035 -196.565 -178.695 ;
        RECT -196.385 -178.935 -195.455 -178.755 ;
        RECT -194.005 -178.935 -193.075 -178.755 ;
        RECT -196.385 -179.260 -196.215 -178.935 ;
        RECT -197.285 -179.430 -196.215 -179.260 ;
        RECT -193.245 -179.260 -193.075 -178.935 ;
        RECT -192.895 -179.035 -192.525 -178.695 ;
        RECT -192.345 -178.935 -191.795 -178.765 ;
        RECT -187.745 -178.935 -187.195 -178.765 ;
        RECT -192.345 -179.260 -192.175 -178.935 ;
        RECT -193.245 -179.430 -192.175 -179.260 ;
        RECT -187.365 -179.260 -187.195 -178.935 ;
        RECT -187.015 -179.035 -186.645 -178.695 ;
        RECT -186.465 -178.935 -185.535 -178.755 ;
        RECT -184.085 -178.935 -183.155 -178.755 ;
        RECT -186.465 -179.260 -186.295 -178.935 ;
        RECT -187.365 -179.430 -186.295 -179.260 ;
        RECT -183.325 -179.260 -183.155 -178.935 ;
        RECT -182.975 -179.035 -182.605 -178.695 ;
        RECT -182.425 -178.935 -181.875 -178.765 ;
        RECT -177.825 -178.935 -177.275 -178.765 ;
        RECT -182.425 -179.260 -182.255 -178.935 ;
        RECT -183.325 -179.430 -182.255 -179.260 ;
        RECT -177.445 -179.260 -177.275 -178.935 ;
        RECT -177.095 -179.035 -176.725 -178.695 ;
        RECT -176.545 -178.935 -175.615 -178.755 ;
        RECT -174.165 -178.935 -173.235 -178.755 ;
        RECT -176.545 -179.260 -176.375 -178.935 ;
        RECT -177.445 -179.430 -176.375 -179.260 ;
        RECT -173.405 -179.260 -173.235 -178.935 ;
        RECT -173.055 -179.035 -172.685 -178.695 ;
        RECT -172.505 -178.935 -171.955 -178.765 ;
        RECT -167.905 -178.935 -167.355 -178.765 ;
        RECT -172.505 -179.260 -172.335 -178.935 ;
        RECT -173.405 -179.430 -172.335 -179.260 ;
        RECT -167.525 -179.260 -167.355 -178.935 ;
        RECT -167.175 -179.035 -166.805 -178.695 ;
        RECT -166.625 -178.935 -165.695 -178.755 ;
        RECT -164.245 -178.935 -163.315 -178.755 ;
        RECT -166.625 -179.260 -166.455 -178.935 ;
        RECT -167.525 -179.430 -166.455 -179.260 ;
        RECT -163.485 -179.260 -163.315 -178.935 ;
        RECT -163.135 -179.035 -162.765 -178.695 ;
        RECT -162.585 -178.935 -162.035 -178.765 ;
        RECT -157.985 -178.935 -157.435 -178.765 ;
        RECT -162.585 -179.260 -162.415 -178.935 ;
        RECT -163.485 -179.430 -162.415 -179.260 ;
        RECT -157.605 -179.260 -157.435 -178.935 ;
        RECT -157.255 -179.035 -156.885 -178.695 ;
        RECT -156.705 -178.935 -155.775 -178.755 ;
        RECT -154.325 -178.935 -153.395 -178.755 ;
        RECT -156.705 -179.260 -156.535 -178.935 ;
        RECT -157.605 -179.430 -156.535 -179.260 ;
        RECT -153.565 -179.260 -153.395 -178.935 ;
        RECT -153.215 -179.035 -152.845 -178.695 ;
        RECT -152.665 -178.935 -152.115 -178.765 ;
        RECT -148.065 -178.935 -147.515 -178.765 ;
        RECT -152.665 -179.260 -152.495 -178.935 ;
        RECT -153.565 -179.430 -152.495 -179.260 ;
        RECT -147.685 -179.260 -147.515 -178.935 ;
        RECT -147.335 -179.035 -146.965 -178.695 ;
        RECT -146.785 -178.935 -145.855 -178.755 ;
        RECT -144.405 -178.935 -143.475 -178.755 ;
        RECT -146.785 -179.260 -146.615 -178.935 ;
        RECT -147.685 -179.430 -146.615 -179.260 ;
        RECT -143.645 -179.260 -143.475 -178.935 ;
        RECT -143.295 -179.035 -142.925 -178.695 ;
        RECT -142.745 -178.935 -142.195 -178.765 ;
        RECT -138.145 -178.935 -137.595 -178.765 ;
        RECT -142.745 -179.260 -142.575 -178.935 ;
        RECT -143.645 -179.430 -142.575 -179.260 ;
        RECT -137.765 -179.260 -137.595 -178.935 ;
        RECT -137.415 -179.035 -137.045 -178.695 ;
        RECT -136.865 -178.935 -135.935 -178.755 ;
        RECT -134.485 -178.935 -133.555 -178.755 ;
        RECT -136.865 -179.260 -136.695 -178.935 ;
        RECT -137.765 -179.430 -136.695 -179.260 ;
        RECT -133.725 -179.260 -133.555 -178.935 ;
        RECT -133.375 -179.035 -133.005 -178.695 ;
        RECT -132.825 -178.935 -132.275 -178.765 ;
        RECT -128.225 -178.935 -127.675 -178.765 ;
        RECT -132.825 -179.260 -132.655 -178.935 ;
        RECT -133.725 -179.430 -132.655 -179.260 ;
        RECT -127.845 -179.260 -127.675 -178.935 ;
        RECT -127.495 -179.035 -127.125 -178.695 ;
        RECT -126.945 -178.935 -126.015 -178.755 ;
        RECT -124.565 -178.935 -123.635 -178.755 ;
        RECT -126.945 -179.260 -126.775 -178.935 ;
        RECT -127.845 -179.430 -126.775 -179.260 ;
        RECT -123.805 -179.260 -123.635 -178.935 ;
        RECT -123.455 -179.035 -123.085 -178.695 ;
        RECT -122.905 -178.935 -122.355 -178.765 ;
        RECT -118.305 -178.935 -117.755 -178.765 ;
        RECT -122.905 -179.260 -122.735 -178.935 ;
        RECT -123.805 -179.430 -122.735 -179.260 ;
        RECT -117.925 -179.260 -117.755 -178.935 ;
        RECT -117.575 -179.035 -117.205 -178.695 ;
        RECT -117.025 -178.935 -116.095 -178.755 ;
        RECT -114.645 -178.935 -113.715 -178.755 ;
        RECT -117.025 -179.260 -116.855 -178.935 ;
        RECT -117.925 -179.430 -116.855 -179.260 ;
        RECT -113.885 -179.260 -113.715 -178.935 ;
        RECT -113.535 -179.035 -113.165 -178.695 ;
        RECT -112.985 -178.935 -112.435 -178.765 ;
        RECT -108.385 -178.935 -107.835 -178.765 ;
        RECT -112.985 -179.260 -112.815 -178.935 ;
        RECT -113.885 -179.430 -112.815 -179.260 ;
        RECT -108.005 -179.260 -107.835 -178.935 ;
        RECT -107.655 -179.035 -107.285 -178.695 ;
        RECT -107.105 -178.935 -106.175 -178.755 ;
        RECT -104.725 -178.935 -103.795 -178.755 ;
        RECT -107.105 -179.260 -106.935 -178.935 ;
        RECT -108.005 -179.430 -106.935 -179.260 ;
        RECT -103.965 -179.260 -103.795 -178.935 ;
        RECT -103.615 -179.035 -103.245 -178.695 ;
        RECT -103.065 -178.935 -102.515 -178.765 ;
        RECT -98.465 -178.935 -97.915 -178.765 ;
        RECT -103.065 -179.260 -102.895 -178.935 ;
        RECT -103.965 -179.430 -102.895 -179.260 ;
        RECT -98.085 -179.260 -97.915 -178.935 ;
        RECT -97.735 -179.035 -97.365 -178.695 ;
        RECT -97.185 -178.935 -96.255 -178.755 ;
        RECT -94.805 -178.935 -93.875 -178.755 ;
        RECT -97.185 -179.260 -97.015 -178.935 ;
        RECT -98.085 -179.430 -97.015 -179.260 ;
        RECT -94.045 -179.260 -93.875 -178.935 ;
        RECT -93.695 -179.035 -93.325 -178.695 ;
        RECT -93.145 -178.935 -92.595 -178.765 ;
        RECT -88.545 -178.935 -87.995 -178.765 ;
        RECT -93.145 -179.260 -92.975 -178.935 ;
        RECT -94.045 -179.430 -92.975 -179.260 ;
        RECT -88.165 -179.260 -87.995 -178.935 ;
        RECT -87.815 -179.035 -87.445 -178.695 ;
        RECT -87.265 -178.935 -86.335 -178.755 ;
        RECT -84.885 -178.935 -83.955 -178.755 ;
        RECT -87.265 -179.260 -87.095 -178.935 ;
        RECT -88.165 -179.430 -87.095 -179.260 ;
        RECT -84.125 -179.260 -83.955 -178.935 ;
        RECT -83.775 -179.035 -83.405 -178.695 ;
        RECT -83.225 -178.935 -82.675 -178.765 ;
        RECT -78.625 -178.935 -78.075 -178.765 ;
        RECT -83.225 -179.260 -83.055 -178.935 ;
        RECT -84.125 -179.430 -83.055 -179.260 ;
        RECT -78.245 -179.260 -78.075 -178.935 ;
        RECT -77.895 -179.035 -77.525 -178.695 ;
        RECT -77.345 -178.935 -76.415 -178.755 ;
        RECT -74.965 -178.935 -74.035 -178.755 ;
        RECT -77.345 -179.260 -77.175 -178.935 ;
        RECT -78.245 -179.430 -77.175 -179.260 ;
        RECT -74.205 -179.260 -74.035 -178.935 ;
        RECT -73.855 -179.035 -73.485 -178.695 ;
        RECT -73.305 -178.935 -72.755 -178.765 ;
        RECT -68.705 -178.935 -68.155 -178.765 ;
        RECT -73.305 -179.260 -73.135 -178.935 ;
        RECT -74.205 -179.430 -73.135 -179.260 ;
        RECT -68.325 -179.260 -68.155 -178.935 ;
        RECT -67.975 -179.035 -67.605 -178.695 ;
        RECT -67.425 -178.935 -66.495 -178.755 ;
        RECT -65.045 -178.935 -64.115 -178.755 ;
        RECT -67.425 -179.260 -67.255 -178.935 ;
        RECT -68.325 -179.430 -67.255 -179.260 ;
        RECT -64.285 -179.260 -64.115 -178.935 ;
        RECT -63.935 -179.035 -63.565 -178.695 ;
        RECT -63.385 -178.935 -62.835 -178.765 ;
        RECT -58.785 -178.935 -58.235 -178.765 ;
        RECT -63.385 -179.260 -63.215 -178.935 ;
        RECT -64.285 -179.430 -63.215 -179.260 ;
        RECT -58.405 -179.260 -58.235 -178.935 ;
        RECT -58.055 -179.035 -57.685 -178.695 ;
        RECT -57.505 -178.935 -56.575 -178.755 ;
        RECT -55.125 -178.935 -54.195 -178.755 ;
        RECT -57.505 -179.260 -57.335 -178.935 ;
        RECT -58.405 -179.430 -57.335 -179.260 ;
        RECT -54.365 -179.260 -54.195 -178.935 ;
        RECT -54.015 -179.035 -53.645 -178.695 ;
        RECT -53.465 -178.935 -52.915 -178.765 ;
        RECT -48.865 -178.935 -48.315 -178.765 ;
        RECT -53.465 -179.260 -53.295 -178.935 ;
        RECT -54.365 -179.430 -53.295 -179.260 ;
        RECT -48.485 -179.260 -48.315 -178.935 ;
        RECT -48.135 -179.035 -47.765 -178.695 ;
        RECT -47.585 -178.935 -46.655 -178.755 ;
        RECT -45.205 -178.935 -44.275 -178.755 ;
        RECT -47.585 -179.260 -47.415 -178.935 ;
        RECT -48.485 -179.430 -47.415 -179.260 ;
        RECT -44.445 -179.260 -44.275 -178.935 ;
        RECT -44.095 -179.035 -43.725 -178.695 ;
        RECT -43.545 -178.935 -42.995 -178.765 ;
        RECT -38.945 -178.935 -38.395 -178.765 ;
        RECT -43.545 -179.260 -43.375 -178.935 ;
        RECT -44.445 -179.430 -43.375 -179.260 ;
        RECT -38.565 -179.260 -38.395 -178.935 ;
        RECT -38.215 -179.035 -37.845 -178.695 ;
        RECT -37.665 -178.935 -36.735 -178.755 ;
        RECT -35.285 -178.935 -34.355 -178.755 ;
        RECT -37.665 -179.260 -37.495 -178.935 ;
        RECT -38.565 -179.430 -37.495 -179.260 ;
        RECT -34.525 -179.260 -34.355 -178.935 ;
        RECT -34.175 -179.035 -33.805 -178.695 ;
        RECT -33.625 -178.935 -33.075 -178.765 ;
        RECT -29.025 -178.935 -28.475 -178.765 ;
        RECT -33.625 -179.260 -33.455 -178.935 ;
        RECT -34.525 -179.430 -33.455 -179.260 ;
        RECT -28.645 -179.260 -28.475 -178.935 ;
        RECT -28.295 -179.035 -27.925 -178.695 ;
        RECT -27.745 -178.935 -26.815 -178.755 ;
        RECT -25.365 -178.935 -24.435 -178.755 ;
        RECT -27.745 -179.260 -27.575 -178.935 ;
        RECT -28.645 -179.430 -27.575 -179.260 ;
        RECT -24.605 -179.260 -24.435 -178.935 ;
        RECT -24.255 -179.035 -23.885 -178.695 ;
        RECT -23.705 -178.935 -23.155 -178.765 ;
        RECT -19.105 -178.935 -18.555 -178.765 ;
        RECT -23.705 -179.260 -23.535 -178.935 ;
        RECT -24.605 -179.430 -23.535 -179.260 ;
        RECT -18.725 -179.260 -18.555 -178.935 ;
        RECT -18.375 -179.035 -18.005 -178.695 ;
        RECT -17.825 -178.935 -16.895 -178.755 ;
        RECT -15.445 -178.935 -14.515 -178.755 ;
        RECT -17.825 -179.260 -17.655 -178.935 ;
        RECT -18.725 -179.430 -17.655 -179.260 ;
        RECT -14.685 -179.260 -14.515 -178.935 ;
        RECT -14.335 -179.035 -13.965 -178.695 ;
        RECT -13.785 -178.935 -13.235 -178.765 ;
        RECT -9.185 -178.935 -8.635 -178.765 ;
        RECT -13.785 -179.260 -13.615 -178.935 ;
        RECT -14.685 -179.430 -13.615 -179.260 ;
        RECT -8.805 -179.260 -8.635 -178.935 ;
        RECT -8.455 -179.035 -8.085 -178.695 ;
        RECT -7.905 -178.935 -6.975 -178.755 ;
        RECT -5.525 -178.935 -4.595 -178.755 ;
        RECT -7.905 -179.260 -7.735 -178.935 ;
        RECT -8.805 -179.430 -7.735 -179.260 ;
        RECT -4.765 -179.260 -4.595 -178.935 ;
        RECT -4.415 -179.035 -4.045 -178.695 ;
        RECT -3.865 -178.935 -3.315 -178.765 ;
        RECT 0.735 -178.935 1.285 -178.765 ;
        RECT -3.865 -179.260 -3.695 -178.935 ;
        RECT -4.765 -179.430 -3.695 -179.260 ;
        RECT 1.115 -179.260 1.285 -178.935 ;
        RECT 1.465 -179.035 1.835 -178.695 ;
        RECT 2.015 -178.935 2.945 -178.755 ;
        RECT 4.395 -178.935 5.325 -178.755 ;
        RECT 2.015 -179.260 2.185 -178.935 ;
        RECT 1.115 -179.430 2.185 -179.260 ;
        RECT 5.155 -179.260 5.325 -178.935 ;
        RECT 5.505 -179.035 5.875 -178.695 ;
        RECT 6.055 -178.935 6.605 -178.765 ;
        RECT 10.655 -178.935 11.205 -178.765 ;
        RECT 6.055 -179.260 6.225 -178.935 ;
        RECT 5.155 -179.430 6.225 -179.260 ;
        RECT 11.035 -179.260 11.205 -178.935 ;
        RECT 11.385 -179.035 11.755 -178.695 ;
        RECT 11.935 -178.935 12.865 -178.755 ;
        RECT 14.315 -178.935 15.245 -178.755 ;
        RECT 11.935 -179.260 12.105 -178.935 ;
        RECT 11.035 -179.430 12.105 -179.260 ;
        RECT 15.075 -179.260 15.245 -178.935 ;
        RECT 15.425 -179.035 15.795 -178.695 ;
        RECT 15.975 -178.935 16.525 -178.765 ;
        RECT 20.575 -178.935 21.125 -178.765 ;
        RECT 15.975 -179.260 16.145 -178.935 ;
        RECT 15.075 -179.430 16.145 -179.260 ;
        RECT 20.955 -179.260 21.125 -178.935 ;
        RECT 21.305 -179.035 21.675 -178.695 ;
        RECT 21.855 -178.935 22.785 -178.755 ;
        RECT 24.235 -178.935 25.165 -178.755 ;
        RECT 21.855 -179.260 22.025 -178.935 ;
        RECT 20.955 -179.430 22.025 -179.260 ;
        RECT 24.995 -179.260 25.165 -178.935 ;
        RECT 25.345 -179.035 25.715 -178.695 ;
        RECT 25.895 -178.935 26.445 -178.765 ;
        RECT 25.895 -179.260 26.065 -178.935 ;
        RECT 26.615 -179.115 26.785 -178.590 ;
        RECT 24.995 -179.430 26.065 -179.260 ;
        RECT -287.285 -179.630 -287.115 -179.445 ;
        RECT -286.140 -179.535 -285.810 -179.430 ;
        RECT -282.210 -179.535 -281.880 -179.430 ;
        RECT -276.220 -179.535 -275.890 -179.430 ;
        RECT -272.290 -179.535 -271.960 -179.430 ;
        RECT -266.300 -179.535 -265.970 -179.430 ;
        RECT -262.370 -179.535 -262.040 -179.430 ;
        RECT -256.380 -179.535 -256.050 -179.430 ;
        RECT -252.450 -179.535 -252.120 -179.430 ;
        RECT -246.460 -179.535 -246.130 -179.430 ;
        RECT -242.530 -179.535 -242.200 -179.430 ;
        RECT -236.540 -179.535 -236.210 -179.430 ;
        RECT -232.610 -179.535 -232.280 -179.430 ;
        RECT -226.620 -179.535 -226.290 -179.430 ;
        RECT -222.690 -179.535 -222.360 -179.430 ;
        RECT -216.700 -179.535 -216.370 -179.430 ;
        RECT -212.770 -179.535 -212.440 -179.430 ;
        RECT -206.780 -179.535 -206.450 -179.430 ;
        RECT -202.850 -179.535 -202.520 -179.430 ;
        RECT -196.860 -179.535 -196.530 -179.430 ;
        RECT -192.930 -179.535 -192.600 -179.430 ;
        RECT -186.940 -179.535 -186.610 -179.430 ;
        RECT -183.010 -179.535 -182.680 -179.430 ;
        RECT -177.020 -179.535 -176.690 -179.430 ;
        RECT -173.090 -179.535 -172.760 -179.430 ;
        RECT -167.100 -179.535 -166.770 -179.430 ;
        RECT -163.170 -179.535 -162.840 -179.430 ;
        RECT -157.180 -179.535 -156.850 -179.430 ;
        RECT -153.250 -179.535 -152.920 -179.430 ;
        RECT -147.260 -179.535 -146.930 -179.430 ;
        RECT -143.330 -179.535 -143.000 -179.430 ;
        RECT -137.340 -179.535 -137.010 -179.430 ;
        RECT -133.410 -179.535 -133.080 -179.430 ;
        RECT -127.420 -179.535 -127.090 -179.430 ;
        RECT -123.490 -179.535 -123.160 -179.430 ;
        RECT -117.500 -179.535 -117.170 -179.430 ;
        RECT -113.570 -179.535 -113.240 -179.430 ;
        RECT -107.580 -179.535 -107.250 -179.430 ;
        RECT -103.650 -179.535 -103.320 -179.430 ;
        RECT -97.660 -179.535 -97.330 -179.430 ;
        RECT -93.730 -179.535 -93.400 -179.430 ;
        RECT -87.740 -179.535 -87.410 -179.430 ;
        RECT -83.810 -179.535 -83.480 -179.430 ;
        RECT -77.820 -179.535 -77.490 -179.430 ;
        RECT -73.890 -179.535 -73.560 -179.430 ;
        RECT -67.900 -179.535 -67.570 -179.430 ;
        RECT -63.970 -179.535 -63.640 -179.430 ;
        RECT -57.980 -179.535 -57.650 -179.430 ;
        RECT -54.050 -179.535 -53.720 -179.430 ;
        RECT -48.060 -179.535 -47.730 -179.430 ;
        RECT -44.130 -179.535 -43.800 -179.430 ;
        RECT -38.140 -179.535 -37.810 -179.430 ;
        RECT -34.210 -179.535 -33.880 -179.430 ;
        RECT -28.220 -179.535 -27.890 -179.430 ;
        RECT -24.290 -179.535 -23.960 -179.430 ;
        RECT -18.300 -179.535 -17.970 -179.430 ;
        RECT -14.370 -179.535 -14.040 -179.430 ;
        RECT -8.380 -179.535 -8.050 -179.430 ;
        RECT -4.450 -179.535 -4.120 -179.430 ;
        RECT 1.540 -179.535 1.870 -179.430 ;
        RECT 5.470 -179.535 5.800 -179.430 ;
        RECT 11.460 -179.535 11.790 -179.430 ;
        RECT 15.390 -179.535 15.720 -179.430 ;
        RECT 21.380 -179.535 21.710 -179.430 ;
        RECT 25.310 -179.535 25.640 -179.430 ;
        RECT 26.235 -179.445 26.785 -179.115 ;
        RECT -287.815 -179.645 -287.115 -179.630 ;
        RECT -287.900 -179.815 -287.115 -179.645 ;
        RECT -287.580 -179.820 -287.115 -179.815 ;
        RECT -287.285 -179.970 -287.115 -179.820 ;
        RECT -283.285 -179.705 -282.380 -179.615 ;
        RECT -281.580 -179.705 -281.075 -179.625 ;
        RECT -283.285 -179.885 -281.075 -179.705 ;
        RECT -273.365 -179.705 -272.460 -179.615 ;
        RECT -271.660 -179.705 -271.155 -179.625 ;
        RECT -273.365 -179.885 -271.155 -179.705 ;
        RECT -263.445 -179.705 -262.540 -179.615 ;
        RECT -261.740 -179.705 -261.235 -179.625 ;
        RECT -263.445 -179.885 -261.235 -179.705 ;
        RECT -253.525 -179.705 -252.620 -179.615 ;
        RECT -251.820 -179.705 -251.315 -179.625 ;
        RECT -253.525 -179.885 -251.315 -179.705 ;
        RECT -243.605 -179.705 -242.700 -179.615 ;
        RECT -241.900 -179.705 -241.395 -179.625 ;
        RECT -243.605 -179.885 -241.395 -179.705 ;
        RECT -233.685 -179.705 -232.780 -179.615 ;
        RECT -231.980 -179.705 -231.475 -179.625 ;
        RECT -233.685 -179.885 -231.475 -179.705 ;
        RECT -223.765 -179.705 -222.860 -179.615 ;
        RECT -222.060 -179.705 -221.555 -179.625 ;
        RECT -223.765 -179.885 -221.555 -179.705 ;
        RECT -213.845 -179.705 -212.940 -179.615 ;
        RECT -212.140 -179.705 -211.635 -179.625 ;
        RECT -213.845 -179.885 -211.635 -179.705 ;
        RECT -203.925 -179.705 -203.020 -179.615 ;
        RECT -202.220 -179.705 -201.715 -179.625 ;
        RECT -203.925 -179.885 -201.715 -179.705 ;
        RECT -194.005 -179.705 -193.100 -179.615 ;
        RECT -192.300 -179.705 -191.795 -179.625 ;
        RECT -194.005 -179.885 -191.795 -179.705 ;
        RECT -184.085 -179.705 -183.180 -179.615 ;
        RECT -182.380 -179.705 -181.875 -179.625 ;
        RECT -184.085 -179.885 -181.875 -179.705 ;
        RECT -174.165 -179.705 -173.260 -179.615 ;
        RECT -172.460 -179.705 -171.955 -179.625 ;
        RECT -174.165 -179.885 -171.955 -179.705 ;
        RECT -164.245 -179.705 -163.340 -179.615 ;
        RECT -162.540 -179.705 -162.035 -179.625 ;
        RECT -164.245 -179.885 -162.035 -179.705 ;
        RECT -154.325 -179.705 -153.420 -179.615 ;
        RECT -152.620 -179.705 -152.115 -179.625 ;
        RECT -154.325 -179.885 -152.115 -179.705 ;
        RECT -144.405 -179.705 -143.500 -179.615 ;
        RECT -142.700 -179.705 -142.195 -179.625 ;
        RECT -144.405 -179.885 -142.195 -179.705 ;
        RECT -134.485 -179.705 -133.580 -179.615 ;
        RECT -132.780 -179.705 -132.275 -179.625 ;
        RECT -134.485 -179.885 -132.275 -179.705 ;
        RECT -124.565 -179.705 -123.660 -179.615 ;
        RECT -122.860 -179.705 -122.355 -179.625 ;
        RECT -124.565 -179.885 -122.355 -179.705 ;
        RECT -114.645 -179.705 -113.740 -179.615 ;
        RECT -112.940 -179.705 -112.435 -179.625 ;
        RECT -114.645 -179.885 -112.435 -179.705 ;
        RECT -104.725 -179.705 -103.820 -179.615 ;
        RECT -103.020 -179.705 -102.515 -179.625 ;
        RECT -104.725 -179.885 -102.515 -179.705 ;
        RECT -94.805 -179.705 -93.900 -179.615 ;
        RECT -93.100 -179.705 -92.595 -179.625 ;
        RECT -94.805 -179.885 -92.595 -179.705 ;
        RECT -84.885 -179.705 -83.980 -179.615 ;
        RECT -83.180 -179.705 -82.675 -179.625 ;
        RECT -84.885 -179.885 -82.675 -179.705 ;
        RECT -74.965 -179.705 -74.060 -179.615 ;
        RECT -73.260 -179.705 -72.755 -179.625 ;
        RECT -74.965 -179.885 -72.755 -179.705 ;
        RECT -65.045 -179.705 -64.140 -179.615 ;
        RECT -63.340 -179.705 -62.835 -179.625 ;
        RECT -65.045 -179.885 -62.835 -179.705 ;
        RECT -55.125 -179.705 -54.220 -179.615 ;
        RECT -53.420 -179.705 -52.915 -179.625 ;
        RECT -55.125 -179.885 -52.915 -179.705 ;
        RECT -45.205 -179.705 -44.300 -179.615 ;
        RECT -43.500 -179.705 -42.995 -179.625 ;
        RECT -45.205 -179.885 -42.995 -179.705 ;
        RECT -35.285 -179.705 -34.380 -179.615 ;
        RECT -33.580 -179.705 -33.075 -179.625 ;
        RECT -35.285 -179.885 -33.075 -179.705 ;
        RECT -25.365 -179.705 -24.460 -179.615 ;
        RECT -23.660 -179.705 -23.155 -179.625 ;
        RECT -25.365 -179.885 -23.155 -179.705 ;
        RECT -15.445 -179.705 -14.540 -179.615 ;
        RECT -13.740 -179.705 -13.235 -179.625 ;
        RECT -15.445 -179.885 -13.235 -179.705 ;
        RECT -5.525 -179.705 -4.620 -179.615 ;
        RECT -3.820 -179.705 -3.315 -179.625 ;
        RECT -5.525 -179.885 -3.315 -179.705 ;
        RECT 4.395 -179.705 5.300 -179.615 ;
        RECT 6.100 -179.705 6.605 -179.625 ;
        RECT 4.395 -179.885 6.605 -179.705 ;
        RECT 14.315 -179.705 15.220 -179.615 ;
        RECT 16.020 -179.705 16.525 -179.625 ;
        RECT 14.315 -179.885 16.525 -179.705 ;
        RECT 24.235 -179.705 25.140 -179.615 ;
        RECT 25.940 -179.705 26.445 -179.625 ;
        RECT 24.235 -179.885 26.445 -179.705 ;
        RECT 26.615 -179.640 26.785 -179.445 ;
        RECT 27.025 -179.640 27.315 -178.920 ;
        RECT 26.615 -179.645 27.315 -179.640 ;
        RECT 26.615 -179.815 27.400 -179.645 ;
        RECT 26.615 -179.820 27.080 -179.815 ;
        RECT 26.615 -179.970 26.785 -179.820 ;
      LAYER mcon ;
        RECT -291.315 94.820 -291.145 94.990 ;
        RECT -290.845 94.825 -290.675 94.995 ;
        RECT -290.020 94.795 -289.850 94.965 ;
        RECT -288.655 94.795 -288.485 94.965 ;
        RECT -280.100 94.795 -279.930 94.965 ;
        RECT -278.735 94.795 -278.565 94.965 ;
        RECT -270.180 94.795 -270.010 94.965 ;
        RECT -268.815 94.795 -268.645 94.965 ;
        RECT -260.260 94.795 -260.090 94.965 ;
        RECT -258.895 94.795 -258.725 94.965 ;
        RECT -250.340 94.795 -250.170 94.965 ;
        RECT -248.975 94.795 -248.805 94.965 ;
        RECT -240.420 94.795 -240.250 94.965 ;
        RECT -239.055 94.795 -238.885 94.965 ;
        RECT -230.500 94.795 -230.330 94.965 ;
        RECT -229.135 94.795 -228.965 94.965 ;
        RECT -220.580 94.795 -220.410 94.965 ;
        RECT -219.215 94.795 -219.045 94.965 ;
        RECT -210.660 94.795 -210.490 94.965 ;
        RECT -209.295 94.795 -209.125 94.965 ;
        RECT -200.740 94.795 -200.570 94.965 ;
        RECT -199.375 94.795 -199.205 94.965 ;
        RECT -190.820 94.795 -190.650 94.965 ;
        RECT -189.455 94.795 -189.285 94.965 ;
        RECT -180.900 94.795 -180.730 94.965 ;
        RECT -179.535 94.795 -179.365 94.965 ;
        RECT -170.980 94.795 -170.810 94.965 ;
        RECT -169.615 94.795 -169.445 94.965 ;
        RECT -161.060 94.795 -160.890 94.965 ;
        RECT -159.695 94.795 -159.525 94.965 ;
        RECT -151.140 94.795 -150.970 94.965 ;
        RECT -149.775 94.795 -149.605 94.965 ;
        RECT -141.220 94.795 -141.050 94.965 ;
        RECT -139.855 94.795 -139.685 94.965 ;
        RECT -131.300 94.795 -131.130 94.965 ;
        RECT -129.935 94.795 -129.765 94.965 ;
        RECT -121.380 94.795 -121.210 94.965 ;
        RECT -120.015 94.795 -119.845 94.965 ;
        RECT -111.460 94.795 -111.290 94.965 ;
        RECT -110.095 94.795 -109.925 94.965 ;
        RECT -101.540 94.795 -101.370 94.965 ;
        RECT -100.175 94.795 -100.005 94.965 ;
        RECT -91.620 94.795 -91.450 94.965 ;
        RECT -90.255 94.795 -90.085 94.965 ;
        RECT -81.700 94.795 -81.530 94.965 ;
        RECT -80.335 94.795 -80.165 94.965 ;
        RECT -71.780 94.795 -71.610 94.965 ;
        RECT -70.415 94.795 -70.245 94.965 ;
        RECT -61.860 94.795 -61.690 94.965 ;
        RECT -60.495 94.795 -60.325 94.965 ;
        RECT -51.940 94.795 -51.770 94.965 ;
        RECT -50.575 94.795 -50.405 94.965 ;
        RECT -42.020 94.795 -41.850 94.965 ;
        RECT -40.655 94.795 -40.485 94.965 ;
        RECT -32.100 94.795 -31.930 94.965 ;
        RECT -30.735 94.795 -30.565 94.965 ;
        RECT -22.180 94.795 -22.010 94.965 ;
        RECT -20.815 94.795 -20.645 94.965 ;
        RECT -12.260 94.795 -12.090 94.965 ;
        RECT -10.895 94.795 -10.725 94.965 ;
        RECT -2.340 94.795 -2.170 94.965 ;
        RECT -0.975 94.795 -0.805 94.965 ;
        RECT 7.580 94.795 7.750 94.965 ;
        RECT 8.945 94.795 9.115 94.965 ;
        RECT 17.500 94.795 17.670 94.965 ;
        RECT 18.865 94.795 19.035 94.965 ;
        RECT -290.845 94.365 -290.675 94.535 ;
        RECT -290.845 93.905 -290.675 94.075 ;
        RECT -289.285 93.945 -289.115 94.115 ;
        RECT -283.425 93.945 -283.255 94.115 ;
        RECT -279.365 93.945 -279.195 94.115 ;
        RECT -273.505 93.945 -273.335 94.115 ;
        RECT -269.445 93.945 -269.275 94.115 ;
        RECT -263.585 93.945 -263.415 94.115 ;
        RECT -259.525 93.945 -259.355 94.115 ;
        RECT -253.665 93.945 -253.495 94.115 ;
        RECT -249.605 93.945 -249.435 94.115 ;
        RECT -243.745 93.945 -243.575 94.115 ;
        RECT -239.685 93.945 -239.515 94.115 ;
        RECT -233.825 93.945 -233.655 94.115 ;
        RECT -229.765 93.945 -229.595 94.115 ;
        RECT -223.905 93.945 -223.735 94.115 ;
        RECT -219.845 93.945 -219.675 94.115 ;
        RECT -213.985 93.945 -213.815 94.115 ;
        RECT -209.925 93.945 -209.755 94.115 ;
        RECT -204.065 93.945 -203.895 94.115 ;
        RECT -200.005 93.945 -199.835 94.115 ;
        RECT -194.145 93.945 -193.975 94.115 ;
        RECT -190.085 93.945 -189.915 94.115 ;
        RECT -184.225 93.945 -184.055 94.115 ;
        RECT -180.165 93.945 -179.995 94.115 ;
        RECT -174.305 93.945 -174.135 94.115 ;
        RECT -170.245 93.945 -170.075 94.115 ;
        RECT -164.385 93.945 -164.215 94.115 ;
        RECT -160.325 93.945 -160.155 94.115 ;
        RECT -154.465 93.945 -154.295 94.115 ;
        RECT -150.405 93.945 -150.235 94.115 ;
        RECT -144.545 93.945 -144.375 94.115 ;
        RECT -140.485 93.945 -140.315 94.115 ;
        RECT -134.625 93.945 -134.455 94.115 ;
        RECT -130.565 93.945 -130.395 94.115 ;
        RECT -124.705 93.945 -124.535 94.115 ;
        RECT -120.645 93.945 -120.475 94.115 ;
        RECT -114.785 93.945 -114.615 94.115 ;
        RECT -110.725 93.945 -110.555 94.115 ;
        RECT -104.865 93.945 -104.695 94.115 ;
        RECT -100.805 93.945 -100.635 94.115 ;
        RECT -94.945 93.945 -94.775 94.115 ;
        RECT -90.885 93.945 -90.715 94.115 ;
        RECT -85.025 93.945 -84.855 94.115 ;
        RECT -80.965 93.945 -80.795 94.115 ;
        RECT -75.105 93.945 -74.935 94.115 ;
        RECT -71.045 93.945 -70.875 94.115 ;
        RECT -65.185 93.945 -65.015 94.115 ;
        RECT -61.125 93.945 -60.955 94.115 ;
        RECT -55.265 93.945 -55.095 94.115 ;
        RECT -51.205 93.945 -51.035 94.115 ;
        RECT -45.345 93.945 -45.175 94.115 ;
        RECT -41.285 93.945 -41.115 94.115 ;
        RECT -35.425 93.945 -35.255 94.115 ;
        RECT -31.365 93.945 -31.195 94.115 ;
        RECT -25.505 93.945 -25.335 94.115 ;
        RECT -21.445 93.945 -21.275 94.115 ;
        RECT -15.585 93.945 -15.415 94.115 ;
        RECT -11.525 93.945 -11.355 94.115 ;
        RECT -5.665 93.945 -5.495 94.115 ;
        RECT -1.605 93.945 -1.435 94.115 ;
        RECT 4.255 93.945 4.425 94.115 ;
        RECT 8.315 93.945 8.485 94.115 ;
        RECT 14.175 93.945 14.345 94.115 ;
        RECT 18.235 93.945 18.405 94.115 ;
        RECT 24.095 93.945 24.265 94.115 ;
        RECT -291.315 93.245 -291.145 93.415 ;
        RECT -290.855 93.245 -290.685 93.415 ;
        RECT -290.395 93.245 -290.225 93.415 ;
        RECT -289.935 93.245 -289.765 93.415 ;
        RECT 24.745 93.245 24.915 93.415 ;
        RECT 25.205 93.245 25.375 93.415 ;
        RECT 25.665 93.245 25.835 93.415 ;
        RECT 26.125 93.245 26.295 93.415 ;
        RECT -289.965 92.525 -289.795 92.695 ;
        RECT -289.980 92.085 -289.810 92.255 ;
        RECT -282.745 92.525 -282.575 92.695 ;
        RECT -287.690 91.685 -287.520 91.855 ;
        RECT -287.705 91.245 -287.535 91.415 ;
        RECT -282.730 92.085 -282.560 92.255 ;
        RECT -285.020 91.685 -284.850 91.855 ;
        RECT -280.045 92.525 -279.875 92.695 ;
        RECT -280.060 92.085 -279.890 92.255 ;
        RECT -272.825 92.525 -272.655 92.695 ;
        RECT -285.005 91.245 -284.835 91.415 ;
        RECT -277.770 91.685 -277.600 91.855 ;
        RECT -277.785 91.245 -277.615 91.415 ;
        RECT -272.810 92.085 -272.640 92.255 ;
        RECT -275.100 91.685 -274.930 91.855 ;
        RECT -270.125 92.525 -269.955 92.695 ;
        RECT -270.140 92.085 -269.970 92.255 ;
        RECT -262.905 92.525 -262.735 92.695 ;
        RECT -275.085 91.245 -274.915 91.415 ;
        RECT -267.850 91.685 -267.680 91.855 ;
        RECT -267.865 91.245 -267.695 91.415 ;
        RECT -262.890 92.085 -262.720 92.255 ;
        RECT -265.180 91.685 -265.010 91.855 ;
        RECT -260.205 92.525 -260.035 92.695 ;
        RECT -260.220 92.085 -260.050 92.255 ;
        RECT -252.985 92.525 -252.815 92.695 ;
        RECT -265.165 91.245 -264.995 91.415 ;
        RECT -257.930 91.685 -257.760 91.855 ;
        RECT -257.945 91.245 -257.775 91.415 ;
        RECT -252.970 92.085 -252.800 92.255 ;
        RECT -255.260 91.685 -255.090 91.855 ;
        RECT -250.285 92.525 -250.115 92.695 ;
        RECT -250.300 92.085 -250.130 92.255 ;
        RECT -243.065 92.525 -242.895 92.695 ;
        RECT -255.245 91.245 -255.075 91.415 ;
        RECT -248.010 91.685 -247.840 91.855 ;
        RECT -248.025 91.245 -247.855 91.415 ;
        RECT -243.050 92.085 -242.880 92.255 ;
        RECT -245.340 91.685 -245.170 91.855 ;
        RECT -240.365 92.525 -240.195 92.695 ;
        RECT -240.380 92.085 -240.210 92.255 ;
        RECT -233.145 92.525 -232.975 92.695 ;
        RECT -245.325 91.245 -245.155 91.415 ;
        RECT -238.090 91.685 -237.920 91.855 ;
        RECT -238.105 91.245 -237.935 91.415 ;
        RECT -233.130 92.085 -232.960 92.255 ;
        RECT -235.420 91.685 -235.250 91.855 ;
        RECT -230.445 92.525 -230.275 92.695 ;
        RECT -230.460 92.085 -230.290 92.255 ;
        RECT -223.225 92.525 -223.055 92.695 ;
        RECT -235.405 91.245 -235.235 91.415 ;
        RECT -228.170 91.685 -228.000 91.855 ;
        RECT -228.185 91.245 -228.015 91.415 ;
        RECT -223.210 92.085 -223.040 92.255 ;
        RECT -225.500 91.685 -225.330 91.855 ;
        RECT -220.525 92.525 -220.355 92.695 ;
        RECT -220.540 92.085 -220.370 92.255 ;
        RECT -213.305 92.525 -213.135 92.695 ;
        RECT -225.485 91.245 -225.315 91.415 ;
        RECT -218.250 91.685 -218.080 91.855 ;
        RECT -218.265 91.245 -218.095 91.415 ;
        RECT -213.290 92.085 -213.120 92.255 ;
        RECT -215.580 91.685 -215.410 91.855 ;
        RECT -210.605 92.525 -210.435 92.695 ;
        RECT -210.620 92.085 -210.450 92.255 ;
        RECT -203.385 92.525 -203.215 92.695 ;
        RECT -215.565 91.245 -215.395 91.415 ;
        RECT -208.330 91.685 -208.160 91.855 ;
        RECT -208.345 91.245 -208.175 91.415 ;
        RECT -203.370 92.085 -203.200 92.255 ;
        RECT -205.660 91.685 -205.490 91.855 ;
        RECT -200.685 92.525 -200.515 92.695 ;
        RECT -200.700 92.085 -200.530 92.255 ;
        RECT -193.465 92.525 -193.295 92.695 ;
        RECT -205.645 91.245 -205.475 91.415 ;
        RECT -198.410 91.685 -198.240 91.855 ;
        RECT -198.425 91.245 -198.255 91.415 ;
        RECT -193.450 92.085 -193.280 92.255 ;
        RECT -195.740 91.685 -195.570 91.855 ;
        RECT -190.765 92.525 -190.595 92.695 ;
        RECT -190.780 92.085 -190.610 92.255 ;
        RECT -183.545 92.525 -183.375 92.695 ;
        RECT -195.725 91.245 -195.555 91.415 ;
        RECT -188.490 91.685 -188.320 91.855 ;
        RECT -188.505 91.245 -188.335 91.415 ;
        RECT -183.530 92.085 -183.360 92.255 ;
        RECT -185.820 91.685 -185.650 91.855 ;
        RECT -180.845 92.525 -180.675 92.695 ;
        RECT -180.860 92.085 -180.690 92.255 ;
        RECT -173.625 92.525 -173.455 92.695 ;
        RECT -185.805 91.245 -185.635 91.415 ;
        RECT -178.570 91.685 -178.400 91.855 ;
        RECT -178.585 91.245 -178.415 91.415 ;
        RECT -173.610 92.085 -173.440 92.255 ;
        RECT -175.900 91.685 -175.730 91.855 ;
        RECT -170.925 92.525 -170.755 92.695 ;
        RECT -170.940 92.085 -170.770 92.255 ;
        RECT -163.705 92.525 -163.535 92.695 ;
        RECT -175.885 91.245 -175.715 91.415 ;
        RECT -168.650 91.685 -168.480 91.855 ;
        RECT -168.665 91.245 -168.495 91.415 ;
        RECT -163.690 92.085 -163.520 92.255 ;
        RECT -165.980 91.685 -165.810 91.855 ;
        RECT -161.005 92.525 -160.835 92.695 ;
        RECT -161.020 92.085 -160.850 92.255 ;
        RECT -153.785 92.525 -153.615 92.695 ;
        RECT -165.965 91.245 -165.795 91.415 ;
        RECT -158.730 91.685 -158.560 91.855 ;
        RECT -158.745 91.245 -158.575 91.415 ;
        RECT -153.770 92.085 -153.600 92.255 ;
        RECT -156.060 91.685 -155.890 91.855 ;
        RECT -151.085 92.525 -150.915 92.695 ;
        RECT -151.100 92.085 -150.930 92.255 ;
        RECT -143.865 92.525 -143.695 92.695 ;
        RECT -156.045 91.245 -155.875 91.415 ;
        RECT -148.810 91.685 -148.640 91.855 ;
        RECT -148.825 91.245 -148.655 91.415 ;
        RECT -143.850 92.085 -143.680 92.255 ;
        RECT -146.140 91.685 -145.970 91.855 ;
        RECT -141.165 92.525 -140.995 92.695 ;
        RECT -141.180 92.085 -141.010 92.255 ;
        RECT -133.945 92.525 -133.775 92.695 ;
        RECT -146.125 91.245 -145.955 91.415 ;
        RECT -138.890 91.685 -138.720 91.855 ;
        RECT -138.905 91.245 -138.735 91.415 ;
        RECT -133.930 92.085 -133.760 92.255 ;
        RECT -136.220 91.685 -136.050 91.855 ;
        RECT -131.245 92.525 -131.075 92.695 ;
        RECT -131.260 92.085 -131.090 92.255 ;
        RECT -124.025 92.525 -123.855 92.695 ;
        RECT -136.205 91.245 -136.035 91.415 ;
        RECT -128.970 91.685 -128.800 91.855 ;
        RECT -128.985 91.245 -128.815 91.415 ;
        RECT -124.010 92.085 -123.840 92.255 ;
        RECT -126.300 91.685 -126.130 91.855 ;
        RECT -121.325 92.525 -121.155 92.695 ;
        RECT -121.340 92.085 -121.170 92.255 ;
        RECT -114.105 92.525 -113.935 92.695 ;
        RECT -126.285 91.245 -126.115 91.415 ;
        RECT -119.050 91.685 -118.880 91.855 ;
        RECT -119.065 91.245 -118.895 91.415 ;
        RECT -114.090 92.085 -113.920 92.255 ;
        RECT -116.380 91.685 -116.210 91.855 ;
        RECT -111.405 92.525 -111.235 92.695 ;
        RECT -111.420 92.085 -111.250 92.255 ;
        RECT -104.185 92.525 -104.015 92.695 ;
        RECT -116.365 91.245 -116.195 91.415 ;
        RECT -109.130 91.685 -108.960 91.855 ;
        RECT -109.145 91.245 -108.975 91.415 ;
        RECT -104.170 92.085 -104.000 92.255 ;
        RECT -106.460 91.685 -106.290 91.855 ;
        RECT -101.485 92.525 -101.315 92.695 ;
        RECT -101.500 92.085 -101.330 92.255 ;
        RECT -94.265 92.525 -94.095 92.695 ;
        RECT -106.445 91.245 -106.275 91.415 ;
        RECT -99.210 91.685 -99.040 91.855 ;
        RECT -99.225 91.245 -99.055 91.415 ;
        RECT -94.250 92.085 -94.080 92.255 ;
        RECT -96.540 91.685 -96.370 91.855 ;
        RECT -91.565 92.525 -91.395 92.695 ;
        RECT -91.580 92.085 -91.410 92.255 ;
        RECT -84.345 92.525 -84.175 92.695 ;
        RECT -96.525 91.245 -96.355 91.415 ;
        RECT -89.290 91.685 -89.120 91.855 ;
        RECT -89.305 91.245 -89.135 91.415 ;
        RECT -84.330 92.085 -84.160 92.255 ;
        RECT -86.620 91.685 -86.450 91.855 ;
        RECT -81.645 92.525 -81.475 92.695 ;
        RECT -81.660 92.085 -81.490 92.255 ;
        RECT -74.425 92.525 -74.255 92.695 ;
        RECT -86.605 91.245 -86.435 91.415 ;
        RECT -79.370 91.685 -79.200 91.855 ;
        RECT -79.385 91.245 -79.215 91.415 ;
        RECT -74.410 92.085 -74.240 92.255 ;
        RECT -76.700 91.685 -76.530 91.855 ;
        RECT -71.725 92.525 -71.555 92.695 ;
        RECT -71.740 92.085 -71.570 92.255 ;
        RECT -64.505 92.525 -64.335 92.695 ;
        RECT -76.685 91.245 -76.515 91.415 ;
        RECT -69.450 91.685 -69.280 91.855 ;
        RECT -69.465 91.245 -69.295 91.415 ;
        RECT -64.490 92.085 -64.320 92.255 ;
        RECT -66.780 91.685 -66.610 91.855 ;
        RECT -61.805 92.525 -61.635 92.695 ;
        RECT -61.820 92.085 -61.650 92.255 ;
        RECT -54.585 92.525 -54.415 92.695 ;
        RECT -66.765 91.245 -66.595 91.415 ;
        RECT -59.530 91.685 -59.360 91.855 ;
        RECT -59.545 91.245 -59.375 91.415 ;
        RECT -54.570 92.085 -54.400 92.255 ;
        RECT -56.860 91.685 -56.690 91.855 ;
        RECT -51.885 92.525 -51.715 92.695 ;
        RECT -51.900 92.085 -51.730 92.255 ;
        RECT -44.665 92.525 -44.495 92.695 ;
        RECT -56.845 91.245 -56.675 91.415 ;
        RECT -49.610 91.685 -49.440 91.855 ;
        RECT -49.625 91.245 -49.455 91.415 ;
        RECT -44.650 92.085 -44.480 92.255 ;
        RECT -46.940 91.685 -46.770 91.855 ;
        RECT -41.965 92.525 -41.795 92.695 ;
        RECT -41.980 92.085 -41.810 92.255 ;
        RECT -34.745 92.525 -34.575 92.695 ;
        RECT -46.925 91.245 -46.755 91.415 ;
        RECT -39.690 91.685 -39.520 91.855 ;
        RECT -39.705 91.245 -39.535 91.415 ;
        RECT -34.730 92.085 -34.560 92.255 ;
        RECT -37.020 91.685 -36.850 91.855 ;
        RECT -32.045 92.525 -31.875 92.695 ;
        RECT -32.060 92.085 -31.890 92.255 ;
        RECT -24.825 92.525 -24.655 92.695 ;
        RECT -37.005 91.245 -36.835 91.415 ;
        RECT -29.770 91.685 -29.600 91.855 ;
        RECT -29.785 91.245 -29.615 91.415 ;
        RECT -24.810 92.085 -24.640 92.255 ;
        RECT -27.100 91.685 -26.930 91.855 ;
        RECT -22.125 92.525 -21.955 92.695 ;
        RECT -22.140 92.085 -21.970 92.255 ;
        RECT -14.905 92.525 -14.735 92.695 ;
        RECT -27.085 91.245 -26.915 91.415 ;
        RECT -19.850 91.685 -19.680 91.855 ;
        RECT -19.865 91.245 -19.695 91.415 ;
        RECT -14.890 92.085 -14.720 92.255 ;
        RECT -17.180 91.685 -17.010 91.855 ;
        RECT -12.205 92.525 -12.035 92.695 ;
        RECT -12.220 92.085 -12.050 92.255 ;
        RECT -4.985 92.525 -4.815 92.695 ;
        RECT -17.165 91.245 -16.995 91.415 ;
        RECT -9.930 91.685 -9.760 91.855 ;
        RECT -9.945 91.245 -9.775 91.415 ;
        RECT -4.970 92.085 -4.800 92.255 ;
        RECT -7.260 91.685 -7.090 91.855 ;
        RECT -2.285 92.525 -2.115 92.695 ;
        RECT -2.300 92.085 -2.130 92.255 ;
        RECT 4.935 92.525 5.105 92.695 ;
        RECT -7.245 91.245 -7.075 91.415 ;
        RECT -0.010 91.685 0.160 91.855 ;
        RECT -0.025 91.245 0.145 91.415 ;
        RECT 4.950 92.085 5.120 92.255 ;
        RECT 2.660 91.685 2.830 91.855 ;
        RECT 7.635 92.525 7.805 92.695 ;
        RECT 7.620 92.085 7.790 92.255 ;
        RECT 14.855 92.525 15.025 92.695 ;
        RECT 2.675 91.245 2.845 91.415 ;
        RECT 9.910 91.685 10.080 91.855 ;
        RECT 9.895 91.245 10.065 91.415 ;
        RECT 14.870 92.085 15.040 92.255 ;
        RECT 12.580 91.685 12.750 91.855 ;
        RECT 17.555 92.525 17.725 92.695 ;
        RECT 17.540 92.085 17.710 92.255 ;
        RECT 24.775 92.525 24.945 92.695 ;
        RECT 12.595 91.245 12.765 91.415 ;
        RECT 19.830 91.685 20.000 91.855 ;
        RECT 19.815 91.245 19.985 91.415 ;
        RECT 24.790 92.085 24.960 92.255 ;
        RECT 22.500 91.685 22.670 91.855 ;
        RECT 22.515 91.245 22.685 91.415 ;
        RECT -291.315 90.525 -291.145 90.695 ;
        RECT -290.855 90.525 -290.685 90.695 ;
        RECT -290.395 90.525 -290.225 90.695 ;
        RECT -289.935 90.525 -289.765 90.695 ;
        RECT -289.545 89.865 -289.375 90.035 ;
        RECT -289.545 89.405 -289.375 89.575 ;
        RECT -288.385 89.825 -288.215 89.995 ;
        RECT -284.325 89.825 -284.155 89.995 ;
        RECT -278.465 89.825 -278.295 89.995 ;
        RECT -274.405 89.825 -274.235 89.995 ;
        RECT -268.545 89.825 -268.375 89.995 ;
        RECT -264.485 89.825 -264.315 89.995 ;
        RECT -258.625 89.825 -258.455 89.995 ;
        RECT -254.565 89.825 -254.395 89.995 ;
        RECT -248.705 89.825 -248.535 89.995 ;
        RECT -244.645 89.825 -244.475 89.995 ;
        RECT -238.785 89.825 -238.615 89.995 ;
        RECT -234.725 89.825 -234.555 89.995 ;
        RECT -228.865 89.825 -228.695 89.995 ;
        RECT -224.805 89.825 -224.635 89.995 ;
        RECT -218.945 89.825 -218.775 89.995 ;
        RECT -214.885 89.825 -214.715 89.995 ;
        RECT -209.025 89.825 -208.855 89.995 ;
        RECT -204.965 89.825 -204.795 89.995 ;
        RECT -199.105 89.825 -198.935 89.995 ;
        RECT -195.045 89.825 -194.875 89.995 ;
        RECT -189.185 89.825 -189.015 89.995 ;
        RECT -185.125 89.825 -184.955 89.995 ;
        RECT -179.265 89.825 -179.095 89.995 ;
        RECT -175.205 89.825 -175.035 89.995 ;
        RECT -169.345 89.825 -169.175 89.995 ;
        RECT -165.285 89.825 -165.115 89.995 ;
        RECT -159.425 89.825 -159.255 89.995 ;
        RECT -155.365 89.825 -155.195 89.995 ;
        RECT -149.505 89.825 -149.335 89.995 ;
        RECT -145.445 89.825 -145.275 89.995 ;
        RECT -139.585 89.825 -139.415 89.995 ;
        RECT -135.525 89.825 -135.355 89.995 ;
        RECT -129.665 89.825 -129.495 89.995 ;
        RECT -125.605 89.825 -125.435 89.995 ;
        RECT -119.745 89.825 -119.575 89.995 ;
        RECT -115.685 89.825 -115.515 89.995 ;
        RECT -109.825 89.825 -109.655 89.995 ;
        RECT -105.765 89.825 -105.595 89.995 ;
        RECT -99.905 89.825 -99.735 89.995 ;
        RECT -95.845 89.825 -95.675 89.995 ;
        RECT -89.985 89.825 -89.815 89.995 ;
        RECT -85.925 89.825 -85.755 89.995 ;
        RECT -80.065 89.825 -79.895 89.995 ;
        RECT -76.005 89.825 -75.835 89.995 ;
        RECT -70.145 89.825 -69.975 89.995 ;
        RECT -66.085 89.825 -65.915 89.995 ;
        RECT -60.225 89.825 -60.055 89.995 ;
        RECT -56.165 89.825 -55.995 89.995 ;
        RECT -50.305 89.825 -50.135 89.995 ;
        RECT -46.245 89.825 -46.075 89.995 ;
        RECT -40.385 89.825 -40.215 89.995 ;
        RECT -36.325 89.825 -36.155 89.995 ;
        RECT -30.465 89.825 -30.295 89.995 ;
        RECT -26.405 89.825 -26.235 89.995 ;
        RECT -20.545 89.825 -20.375 89.995 ;
        RECT -16.485 89.825 -16.315 89.995 ;
        RECT -10.625 89.825 -10.455 89.995 ;
        RECT -6.565 89.825 -6.395 89.995 ;
        RECT -0.705 89.825 -0.535 89.995 ;
        RECT 3.355 89.825 3.525 89.995 ;
        RECT 9.215 89.825 9.385 89.995 ;
        RECT 13.275 89.825 13.445 89.995 ;
        RECT 19.135 89.825 19.305 89.995 ;
        RECT 23.195 89.825 23.365 89.995 ;
        RECT 24.355 89.865 24.525 90.035 ;
        RECT 24.355 89.405 24.525 89.575 ;
        RECT -290.015 88.955 -289.845 89.125 ;
        RECT -289.545 88.945 -289.375 89.115 ;
        RECT -285.060 88.975 -284.890 89.145 ;
        RECT -283.695 88.975 -283.525 89.145 ;
        RECT -275.140 88.975 -274.970 89.145 ;
        RECT -273.775 88.975 -273.605 89.145 ;
        RECT -265.220 88.975 -265.050 89.145 ;
        RECT -263.855 88.975 -263.685 89.145 ;
        RECT -255.300 88.975 -255.130 89.145 ;
        RECT -253.935 88.975 -253.765 89.145 ;
        RECT -245.380 88.975 -245.210 89.145 ;
        RECT -244.015 88.975 -243.845 89.145 ;
        RECT -235.460 88.975 -235.290 89.145 ;
        RECT -234.095 88.975 -233.925 89.145 ;
        RECT -225.540 88.975 -225.370 89.145 ;
        RECT -224.175 88.975 -224.005 89.145 ;
        RECT -215.620 88.975 -215.450 89.145 ;
        RECT -214.255 88.975 -214.085 89.145 ;
        RECT -205.700 88.975 -205.530 89.145 ;
        RECT -204.335 88.975 -204.165 89.145 ;
        RECT -195.780 88.975 -195.610 89.145 ;
        RECT -194.415 88.975 -194.245 89.145 ;
        RECT -185.860 88.975 -185.690 89.145 ;
        RECT -184.495 88.975 -184.325 89.145 ;
        RECT -175.940 88.975 -175.770 89.145 ;
        RECT -174.575 88.975 -174.405 89.145 ;
        RECT -166.020 88.975 -165.850 89.145 ;
        RECT -164.655 88.975 -164.485 89.145 ;
        RECT -156.100 88.975 -155.930 89.145 ;
        RECT -154.735 88.975 -154.565 89.145 ;
        RECT -146.180 88.975 -146.010 89.145 ;
        RECT -144.815 88.975 -144.645 89.145 ;
        RECT -136.260 88.975 -136.090 89.145 ;
        RECT -134.895 88.975 -134.725 89.145 ;
        RECT -126.340 88.975 -126.170 89.145 ;
        RECT -124.975 88.975 -124.805 89.145 ;
        RECT -116.420 88.975 -116.250 89.145 ;
        RECT -115.055 88.975 -114.885 89.145 ;
        RECT -106.500 88.975 -106.330 89.145 ;
        RECT -105.135 88.975 -104.965 89.145 ;
        RECT -96.580 88.975 -96.410 89.145 ;
        RECT -95.215 88.975 -95.045 89.145 ;
        RECT -86.660 88.975 -86.490 89.145 ;
        RECT -85.295 88.975 -85.125 89.145 ;
        RECT -76.740 88.975 -76.570 89.145 ;
        RECT -75.375 88.975 -75.205 89.145 ;
        RECT -66.820 88.975 -66.650 89.145 ;
        RECT -65.455 88.975 -65.285 89.145 ;
        RECT -56.900 88.975 -56.730 89.145 ;
        RECT -55.535 88.975 -55.365 89.145 ;
        RECT -46.980 88.975 -46.810 89.145 ;
        RECT -45.615 88.975 -45.445 89.145 ;
        RECT -37.060 88.975 -36.890 89.145 ;
        RECT -35.695 88.975 -35.525 89.145 ;
        RECT -27.140 88.975 -26.970 89.145 ;
        RECT -25.775 88.975 -25.605 89.145 ;
        RECT -17.220 88.975 -17.050 89.145 ;
        RECT -15.855 88.975 -15.685 89.145 ;
        RECT -7.300 88.975 -7.130 89.145 ;
        RECT -5.935 88.975 -5.765 89.145 ;
        RECT 2.620 88.975 2.790 89.145 ;
        RECT 3.985 88.975 4.155 89.145 ;
        RECT 12.540 88.975 12.710 89.145 ;
        RECT 13.905 88.975 14.075 89.145 ;
        RECT 22.460 88.975 22.630 89.145 ;
        RECT 23.825 88.975 23.995 89.145 ;
        RECT 24.355 88.945 24.525 89.115 ;
        RECT 24.825 88.955 24.995 89.125 ;
        RECT -291.065 7.110 -290.895 7.280 ;
        RECT -290.595 7.115 -290.425 7.285 ;
        RECT -289.770 7.085 -289.600 7.255 ;
        RECT -288.405 7.085 -288.235 7.255 ;
        RECT -279.850 7.085 -279.680 7.255 ;
        RECT -278.485 7.085 -278.315 7.255 ;
        RECT -269.930 7.085 -269.760 7.255 ;
        RECT -268.565 7.085 -268.395 7.255 ;
        RECT -260.010 7.085 -259.840 7.255 ;
        RECT -258.645 7.085 -258.475 7.255 ;
        RECT -250.090 7.085 -249.920 7.255 ;
        RECT -248.725 7.085 -248.555 7.255 ;
        RECT -240.170 7.085 -240.000 7.255 ;
        RECT -238.805 7.085 -238.635 7.255 ;
        RECT -230.250 7.085 -230.080 7.255 ;
        RECT -228.885 7.085 -228.715 7.255 ;
        RECT -220.330 7.085 -220.160 7.255 ;
        RECT -218.965 7.085 -218.795 7.255 ;
        RECT -210.410 7.085 -210.240 7.255 ;
        RECT -209.045 7.085 -208.875 7.255 ;
        RECT -200.490 7.085 -200.320 7.255 ;
        RECT -199.125 7.085 -198.955 7.255 ;
        RECT -190.570 7.085 -190.400 7.255 ;
        RECT -189.205 7.085 -189.035 7.255 ;
        RECT -180.650 7.085 -180.480 7.255 ;
        RECT -179.285 7.085 -179.115 7.255 ;
        RECT -170.730 7.085 -170.560 7.255 ;
        RECT -169.365 7.085 -169.195 7.255 ;
        RECT -160.810 7.085 -160.640 7.255 ;
        RECT -159.445 7.085 -159.275 7.255 ;
        RECT -150.890 7.085 -150.720 7.255 ;
        RECT -149.525 7.085 -149.355 7.255 ;
        RECT -140.970 7.085 -140.800 7.255 ;
        RECT -139.605 7.085 -139.435 7.255 ;
        RECT -131.050 7.085 -130.880 7.255 ;
        RECT -129.685 7.085 -129.515 7.255 ;
        RECT -121.130 7.085 -120.960 7.255 ;
        RECT -119.765 7.085 -119.595 7.255 ;
        RECT -111.210 7.085 -111.040 7.255 ;
        RECT -109.845 7.085 -109.675 7.255 ;
        RECT -101.290 7.085 -101.120 7.255 ;
        RECT -99.925 7.085 -99.755 7.255 ;
        RECT -91.370 7.085 -91.200 7.255 ;
        RECT -90.005 7.085 -89.835 7.255 ;
        RECT -81.450 7.085 -81.280 7.255 ;
        RECT -80.085 7.085 -79.915 7.255 ;
        RECT -71.530 7.085 -71.360 7.255 ;
        RECT -70.165 7.085 -69.995 7.255 ;
        RECT -61.610 7.085 -61.440 7.255 ;
        RECT -60.245 7.085 -60.075 7.255 ;
        RECT -51.690 7.085 -51.520 7.255 ;
        RECT -50.325 7.085 -50.155 7.255 ;
        RECT -41.770 7.085 -41.600 7.255 ;
        RECT -40.405 7.085 -40.235 7.255 ;
        RECT -31.850 7.085 -31.680 7.255 ;
        RECT -30.485 7.085 -30.315 7.255 ;
        RECT -21.930 7.085 -21.760 7.255 ;
        RECT -20.565 7.085 -20.395 7.255 ;
        RECT -12.010 7.085 -11.840 7.255 ;
        RECT -10.645 7.085 -10.475 7.255 ;
        RECT -2.090 7.085 -1.920 7.255 ;
        RECT -0.725 7.085 -0.555 7.255 ;
        RECT 7.830 7.085 8.000 7.255 ;
        RECT 9.195 7.085 9.365 7.255 ;
        RECT 17.750 7.085 17.920 7.255 ;
        RECT 19.115 7.085 19.285 7.255 ;
        RECT -290.595 6.655 -290.425 6.825 ;
        RECT -290.595 6.195 -290.425 6.365 ;
        RECT -289.035 6.235 -288.865 6.405 ;
        RECT -283.175 6.235 -283.005 6.405 ;
        RECT -279.115 6.235 -278.945 6.405 ;
        RECT -273.255 6.235 -273.085 6.405 ;
        RECT -269.195 6.235 -269.025 6.405 ;
        RECT -263.335 6.235 -263.165 6.405 ;
        RECT -259.275 6.235 -259.105 6.405 ;
        RECT -253.415 6.235 -253.245 6.405 ;
        RECT -249.355 6.235 -249.185 6.405 ;
        RECT -243.495 6.235 -243.325 6.405 ;
        RECT -239.435 6.235 -239.265 6.405 ;
        RECT -233.575 6.235 -233.405 6.405 ;
        RECT -229.515 6.235 -229.345 6.405 ;
        RECT -223.655 6.235 -223.485 6.405 ;
        RECT -219.595 6.235 -219.425 6.405 ;
        RECT -213.735 6.235 -213.565 6.405 ;
        RECT -209.675 6.235 -209.505 6.405 ;
        RECT -203.815 6.235 -203.645 6.405 ;
        RECT -199.755 6.235 -199.585 6.405 ;
        RECT -193.895 6.235 -193.725 6.405 ;
        RECT -189.835 6.235 -189.665 6.405 ;
        RECT -183.975 6.235 -183.805 6.405 ;
        RECT -179.915 6.235 -179.745 6.405 ;
        RECT -174.055 6.235 -173.885 6.405 ;
        RECT -169.995 6.235 -169.825 6.405 ;
        RECT -164.135 6.235 -163.965 6.405 ;
        RECT -160.075 6.235 -159.905 6.405 ;
        RECT -154.215 6.235 -154.045 6.405 ;
        RECT -150.155 6.235 -149.985 6.405 ;
        RECT -144.295 6.235 -144.125 6.405 ;
        RECT -140.235 6.235 -140.065 6.405 ;
        RECT -134.375 6.235 -134.205 6.405 ;
        RECT -130.315 6.235 -130.145 6.405 ;
        RECT -124.455 6.235 -124.285 6.405 ;
        RECT -120.395 6.235 -120.225 6.405 ;
        RECT -114.535 6.235 -114.365 6.405 ;
        RECT -110.475 6.235 -110.305 6.405 ;
        RECT -104.615 6.235 -104.445 6.405 ;
        RECT -100.555 6.235 -100.385 6.405 ;
        RECT -94.695 6.235 -94.525 6.405 ;
        RECT -90.635 6.235 -90.465 6.405 ;
        RECT -84.775 6.235 -84.605 6.405 ;
        RECT -80.715 6.235 -80.545 6.405 ;
        RECT -74.855 6.235 -74.685 6.405 ;
        RECT -70.795 6.235 -70.625 6.405 ;
        RECT -64.935 6.235 -64.765 6.405 ;
        RECT -60.875 6.235 -60.705 6.405 ;
        RECT -55.015 6.235 -54.845 6.405 ;
        RECT -50.955 6.235 -50.785 6.405 ;
        RECT -45.095 6.235 -44.925 6.405 ;
        RECT -41.035 6.235 -40.865 6.405 ;
        RECT -35.175 6.235 -35.005 6.405 ;
        RECT -31.115 6.235 -30.945 6.405 ;
        RECT -25.255 6.235 -25.085 6.405 ;
        RECT -21.195 6.235 -21.025 6.405 ;
        RECT -15.335 6.235 -15.165 6.405 ;
        RECT -11.275 6.235 -11.105 6.405 ;
        RECT -5.415 6.235 -5.245 6.405 ;
        RECT -1.355 6.235 -1.185 6.405 ;
        RECT 4.505 6.235 4.675 6.405 ;
        RECT 8.565 6.235 8.735 6.405 ;
        RECT 14.425 6.235 14.595 6.405 ;
        RECT 18.485 6.235 18.655 6.405 ;
        RECT 24.345 6.235 24.515 6.405 ;
        RECT -291.065 5.535 -290.895 5.705 ;
        RECT -290.605 5.535 -290.435 5.705 ;
        RECT -290.145 5.535 -289.975 5.705 ;
        RECT -289.685 5.535 -289.515 5.705 ;
        RECT 24.995 5.535 25.165 5.705 ;
        RECT 25.455 5.535 25.625 5.705 ;
        RECT 25.915 5.535 26.085 5.705 ;
        RECT 26.375 5.535 26.545 5.705 ;
        RECT -289.715 4.815 -289.545 4.985 ;
        RECT -289.730 4.375 -289.560 4.545 ;
        RECT -282.495 4.815 -282.325 4.985 ;
        RECT -287.440 3.975 -287.270 4.145 ;
        RECT -287.455 3.535 -287.285 3.705 ;
        RECT -282.480 4.375 -282.310 4.545 ;
        RECT -284.770 3.975 -284.600 4.145 ;
        RECT -279.795 4.815 -279.625 4.985 ;
        RECT -279.810 4.375 -279.640 4.545 ;
        RECT -272.575 4.815 -272.405 4.985 ;
        RECT -284.755 3.535 -284.585 3.705 ;
        RECT -277.520 3.975 -277.350 4.145 ;
        RECT -277.535 3.535 -277.365 3.705 ;
        RECT -272.560 4.375 -272.390 4.545 ;
        RECT -274.850 3.975 -274.680 4.145 ;
        RECT -269.875 4.815 -269.705 4.985 ;
        RECT -269.890 4.375 -269.720 4.545 ;
        RECT -262.655 4.815 -262.485 4.985 ;
        RECT -274.835 3.535 -274.665 3.705 ;
        RECT -267.600 3.975 -267.430 4.145 ;
        RECT -267.615 3.535 -267.445 3.705 ;
        RECT -262.640 4.375 -262.470 4.545 ;
        RECT -264.930 3.975 -264.760 4.145 ;
        RECT -259.955 4.815 -259.785 4.985 ;
        RECT -259.970 4.375 -259.800 4.545 ;
        RECT -252.735 4.815 -252.565 4.985 ;
        RECT -264.915 3.535 -264.745 3.705 ;
        RECT -257.680 3.975 -257.510 4.145 ;
        RECT -257.695 3.535 -257.525 3.705 ;
        RECT -252.720 4.375 -252.550 4.545 ;
        RECT -255.010 3.975 -254.840 4.145 ;
        RECT -250.035 4.815 -249.865 4.985 ;
        RECT -250.050 4.375 -249.880 4.545 ;
        RECT -242.815 4.815 -242.645 4.985 ;
        RECT -254.995 3.535 -254.825 3.705 ;
        RECT -247.760 3.975 -247.590 4.145 ;
        RECT -247.775 3.535 -247.605 3.705 ;
        RECT -242.800 4.375 -242.630 4.545 ;
        RECT -245.090 3.975 -244.920 4.145 ;
        RECT -240.115 4.815 -239.945 4.985 ;
        RECT -240.130 4.375 -239.960 4.545 ;
        RECT -232.895 4.815 -232.725 4.985 ;
        RECT -245.075 3.535 -244.905 3.705 ;
        RECT -237.840 3.975 -237.670 4.145 ;
        RECT -237.855 3.535 -237.685 3.705 ;
        RECT -232.880 4.375 -232.710 4.545 ;
        RECT -235.170 3.975 -235.000 4.145 ;
        RECT -230.195 4.815 -230.025 4.985 ;
        RECT -230.210 4.375 -230.040 4.545 ;
        RECT -222.975 4.815 -222.805 4.985 ;
        RECT -235.155 3.535 -234.985 3.705 ;
        RECT -227.920 3.975 -227.750 4.145 ;
        RECT -227.935 3.535 -227.765 3.705 ;
        RECT -222.960 4.375 -222.790 4.545 ;
        RECT -225.250 3.975 -225.080 4.145 ;
        RECT -220.275 4.815 -220.105 4.985 ;
        RECT -220.290 4.375 -220.120 4.545 ;
        RECT -213.055 4.815 -212.885 4.985 ;
        RECT -225.235 3.535 -225.065 3.705 ;
        RECT -218.000 3.975 -217.830 4.145 ;
        RECT -218.015 3.535 -217.845 3.705 ;
        RECT -213.040 4.375 -212.870 4.545 ;
        RECT -215.330 3.975 -215.160 4.145 ;
        RECT -210.355 4.815 -210.185 4.985 ;
        RECT -210.370 4.375 -210.200 4.545 ;
        RECT -203.135 4.815 -202.965 4.985 ;
        RECT -215.315 3.535 -215.145 3.705 ;
        RECT -208.080 3.975 -207.910 4.145 ;
        RECT -208.095 3.535 -207.925 3.705 ;
        RECT -203.120 4.375 -202.950 4.545 ;
        RECT -205.410 3.975 -205.240 4.145 ;
        RECT -200.435 4.815 -200.265 4.985 ;
        RECT -200.450 4.375 -200.280 4.545 ;
        RECT -193.215 4.815 -193.045 4.985 ;
        RECT -205.395 3.535 -205.225 3.705 ;
        RECT -198.160 3.975 -197.990 4.145 ;
        RECT -198.175 3.535 -198.005 3.705 ;
        RECT -193.200 4.375 -193.030 4.545 ;
        RECT -195.490 3.975 -195.320 4.145 ;
        RECT -190.515 4.815 -190.345 4.985 ;
        RECT -190.530 4.375 -190.360 4.545 ;
        RECT -183.295 4.815 -183.125 4.985 ;
        RECT -195.475 3.535 -195.305 3.705 ;
        RECT -188.240 3.975 -188.070 4.145 ;
        RECT -188.255 3.535 -188.085 3.705 ;
        RECT -183.280 4.375 -183.110 4.545 ;
        RECT -185.570 3.975 -185.400 4.145 ;
        RECT -180.595 4.815 -180.425 4.985 ;
        RECT -180.610 4.375 -180.440 4.545 ;
        RECT -173.375 4.815 -173.205 4.985 ;
        RECT -185.555 3.535 -185.385 3.705 ;
        RECT -178.320 3.975 -178.150 4.145 ;
        RECT -178.335 3.535 -178.165 3.705 ;
        RECT -173.360 4.375 -173.190 4.545 ;
        RECT -175.650 3.975 -175.480 4.145 ;
        RECT -170.675 4.815 -170.505 4.985 ;
        RECT -170.690 4.375 -170.520 4.545 ;
        RECT -163.455 4.815 -163.285 4.985 ;
        RECT -175.635 3.535 -175.465 3.705 ;
        RECT -168.400 3.975 -168.230 4.145 ;
        RECT -168.415 3.535 -168.245 3.705 ;
        RECT -163.440 4.375 -163.270 4.545 ;
        RECT -165.730 3.975 -165.560 4.145 ;
        RECT -160.755 4.815 -160.585 4.985 ;
        RECT -160.770 4.375 -160.600 4.545 ;
        RECT -153.535 4.815 -153.365 4.985 ;
        RECT -165.715 3.535 -165.545 3.705 ;
        RECT -158.480 3.975 -158.310 4.145 ;
        RECT -158.495 3.535 -158.325 3.705 ;
        RECT -153.520 4.375 -153.350 4.545 ;
        RECT -155.810 3.975 -155.640 4.145 ;
        RECT -150.835 4.815 -150.665 4.985 ;
        RECT -150.850 4.375 -150.680 4.545 ;
        RECT -143.615 4.815 -143.445 4.985 ;
        RECT -155.795 3.535 -155.625 3.705 ;
        RECT -148.560 3.975 -148.390 4.145 ;
        RECT -148.575 3.535 -148.405 3.705 ;
        RECT -143.600 4.375 -143.430 4.545 ;
        RECT -145.890 3.975 -145.720 4.145 ;
        RECT -140.915 4.815 -140.745 4.985 ;
        RECT -140.930 4.375 -140.760 4.545 ;
        RECT -133.695 4.815 -133.525 4.985 ;
        RECT -145.875 3.535 -145.705 3.705 ;
        RECT -138.640 3.975 -138.470 4.145 ;
        RECT -138.655 3.535 -138.485 3.705 ;
        RECT -133.680 4.375 -133.510 4.545 ;
        RECT -135.970 3.975 -135.800 4.145 ;
        RECT -130.995 4.815 -130.825 4.985 ;
        RECT -131.010 4.375 -130.840 4.545 ;
        RECT -123.775 4.815 -123.605 4.985 ;
        RECT -135.955 3.535 -135.785 3.705 ;
        RECT -128.720 3.975 -128.550 4.145 ;
        RECT -128.735 3.535 -128.565 3.705 ;
        RECT -123.760 4.375 -123.590 4.545 ;
        RECT -126.050 3.975 -125.880 4.145 ;
        RECT -121.075 4.815 -120.905 4.985 ;
        RECT -121.090 4.375 -120.920 4.545 ;
        RECT -113.855 4.815 -113.685 4.985 ;
        RECT -126.035 3.535 -125.865 3.705 ;
        RECT -118.800 3.975 -118.630 4.145 ;
        RECT -118.815 3.535 -118.645 3.705 ;
        RECT -113.840 4.375 -113.670 4.545 ;
        RECT -116.130 3.975 -115.960 4.145 ;
        RECT -111.155 4.815 -110.985 4.985 ;
        RECT -111.170 4.375 -111.000 4.545 ;
        RECT -103.935 4.815 -103.765 4.985 ;
        RECT -116.115 3.535 -115.945 3.705 ;
        RECT -108.880 3.975 -108.710 4.145 ;
        RECT -108.895 3.535 -108.725 3.705 ;
        RECT -103.920 4.375 -103.750 4.545 ;
        RECT -106.210 3.975 -106.040 4.145 ;
        RECT -101.235 4.815 -101.065 4.985 ;
        RECT -101.250 4.375 -101.080 4.545 ;
        RECT -94.015 4.815 -93.845 4.985 ;
        RECT -106.195 3.535 -106.025 3.705 ;
        RECT -98.960 3.975 -98.790 4.145 ;
        RECT -98.975 3.535 -98.805 3.705 ;
        RECT -94.000 4.375 -93.830 4.545 ;
        RECT -96.290 3.975 -96.120 4.145 ;
        RECT -91.315 4.815 -91.145 4.985 ;
        RECT -91.330 4.375 -91.160 4.545 ;
        RECT -84.095 4.815 -83.925 4.985 ;
        RECT -96.275 3.535 -96.105 3.705 ;
        RECT -89.040 3.975 -88.870 4.145 ;
        RECT -89.055 3.535 -88.885 3.705 ;
        RECT -84.080 4.375 -83.910 4.545 ;
        RECT -86.370 3.975 -86.200 4.145 ;
        RECT -81.395 4.815 -81.225 4.985 ;
        RECT -81.410 4.375 -81.240 4.545 ;
        RECT -74.175 4.815 -74.005 4.985 ;
        RECT -86.355 3.535 -86.185 3.705 ;
        RECT -79.120 3.975 -78.950 4.145 ;
        RECT -79.135 3.535 -78.965 3.705 ;
        RECT -74.160 4.375 -73.990 4.545 ;
        RECT -76.450 3.975 -76.280 4.145 ;
        RECT -71.475 4.815 -71.305 4.985 ;
        RECT -71.490 4.375 -71.320 4.545 ;
        RECT -64.255 4.815 -64.085 4.985 ;
        RECT -76.435 3.535 -76.265 3.705 ;
        RECT -69.200 3.975 -69.030 4.145 ;
        RECT -69.215 3.535 -69.045 3.705 ;
        RECT -64.240 4.375 -64.070 4.545 ;
        RECT -66.530 3.975 -66.360 4.145 ;
        RECT -61.555 4.815 -61.385 4.985 ;
        RECT -61.570 4.375 -61.400 4.545 ;
        RECT -54.335 4.815 -54.165 4.985 ;
        RECT -66.515 3.535 -66.345 3.705 ;
        RECT -59.280 3.975 -59.110 4.145 ;
        RECT -59.295 3.535 -59.125 3.705 ;
        RECT -54.320 4.375 -54.150 4.545 ;
        RECT -56.610 3.975 -56.440 4.145 ;
        RECT -51.635 4.815 -51.465 4.985 ;
        RECT -51.650 4.375 -51.480 4.545 ;
        RECT -44.415 4.815 -44.245 4.985 ;
        RECT -56.595 3.535 -56.425 3.705 ;
        RECT -49.360 3.975 -49.190 4.145 ;
        RECT -49.375 3.535 -49.205 3.705 ;
        RECT -44.400 4.375 -44.230 4.545 ;
        RECT -46.690 3.975 -46.520 4.145 ;
        RECT -41.715 4.815 -41.545 4.985 ;
        RECT -41.730 4.375 -41.560 4.545 ;
        RECT -34.495 4.815 -34.325 4.985 ;
        RECT -46.675 3.535 -46.505 3.705 ;
        RECT -39.440 3.975 -39.270 4.145 ;
        RECT -39.455 3.535 -39.285 3.705 ;
        RECT -34.480 4.375 -34.310 4.545 ;
        RECT -36.770 3.975 -36.600 4.145 ;
        RECT -31.795 4.815 -31.625 4.985 ;
        RECT -31.810 4.375 -31.640 4.545 ;
        RECT -24.575 4.815 -24.405 4.985 ;
        RECT -36.755 3.535 -36.585 3.705 ;
        RECT -29.520 3.975 -29.350 4.145 ;
        RECT -29.535 3.535 -29.365 3.705 ;
        RECT -24.560 4.375 -24.390 4.545 ;
        RECT -26.850 3.975 -26.680 4.145 ;
        RECT -21.875 4.815 -21.705 4.985 ;
        RECT -21.890 4.375 -21.720 4.545 ;
        RECT -14.655 4.815 -14.485 4.985 ;
        RECT -26.835 3.535 -26.665 3.705 ;
        RECT -19.600 3.975 -19.430 4.145 ;
        RECT -19.615 3.535 -19.445 3.705 ;
        RECT -14.640 4.375 -14.470 4.545 ;
        RECT -16.930 3.975 -16.760 4.145 ;
        RECT -11.955 4.815 -11.785 4.985 ;
        RECT -11.970 4.375 -11.800 4.545 ;
        RECT -4.735 4.815 -4.565 4.985 ;
        RECT -16.915 3.535 -16.745 3.705 ;
        RECT -9.680 3.975 -9.510 4.145 ;
        RECT -9.695 3.535 -9.525 3.705 ;
        RECT -4.720 4.375 -4.550 4.545 ;
        RECT -7.010 3.975 -6.840 4.145 ;
        RECT -2.035 4.815 -1.865 4.985 ;
        RECT -2.050 4.375 -1.880 4.545 ;
        RECT 5.185 4.815 5.355 4.985 ;
        RECT -6.995 3.535 -6.825 3.705 ;
        RECT 0.240 3.975 0.410 4.145 ;
        RECT 0.225 3.535 0.395 3.705 ;
        RECT 5.200 4.375 5.370 4.545 ;
        RECT 2.910 3.975 3.080 4.145 ;
        RECT 7.885 4.815 8.055 4.985 ;
        RECT 7.870 4.375 8.040 4.545 ;
        RECT 15.105 4.815 15.275 4.985 ;
        RECT 2.925 3.535 3.095 3.705 ;
        RECT 10.160 3.975 10.330 4.145 ;
        RECT 10.145 3.535 10.315 3.705 ;
        RECT 15.120 4.375 15.290 4.545 ;
        RECT 12.830 3.975 13.000 4.145 ;
        RECT 17.805 4.815 17.975 4.985 ;
        RECT 17.790 4.375 17.960 4.545 ;
        RECT 25.025 4.815 25.195 4.985 ;
        RECT 12.845 3.535 13.015 3.705 ;
        RECT 20.080 3.975 20.250 4.145 ;
        RECT 20.065 3.535 20.235 3.705 ;
        RECT 25.040 4.375 25.210 4.545 ;
        RECT 22.750 3.975 22.920 4.145 ;
        RECT 22.765 3.535 22.935 3.705 ;
        RECT -291.065 2.815 -290.895 2.985 ;
        RECT -290.605 2.815 -290.435 2.985 ;
        RECT -290.145 2.815 -289.975 2.985 ;
        RECT -289.685 2.815 -289.515 2.985 ;
        RECT -289.295 2.155 -289.125 2.325 ;
        RECT -289.295 1.695 -289.125 1.865 ;
        RECT -288.135 2.115 -287.965 2.285 ;
        RECT -284.075 2.115 -283.905 2.285 ;
        RECT -278.215 2.115 -278.045 2.285 ;
        RECT -274.155 2.115 -273.985 2.285 ;
        RECT -268.295 2.115 -268.125 2.285 ;
        RECT -264.235 2.115 -264.065 2.285 ;
        RECT -258.375 2.115 -258.205 2.285 ;
        RECT -254.315 2.115 -254.145 2.285 ;
        RECT -248.455 2.115 -248.285 2.285 ;
        RECT -244.395 2.115 -244.225 2.285 ;
        RECT -238.535 2.115 -238.365 2.285 ;
        RECT -234.475 2.115 -234.305 2.285 ;
        RECT -228.615 2.115 -228.445 2.285 ;
        RECT -224.555 2.115 -224.385 2.285 ;
        RECT -218.695 2.115 -218.525 2.285 ;
        RECT -214.635 2.115 -214.465 2.285 ;
        RECT -208.775 2.115 -208.605 2.285 ;
        RECT -204.715 2.115 -204.545 2.285 ;
        RECT -198.855 2.115 -198.685 2.285 ;
        RECT -194.795 2.115 -194.625 2.285 ;
        RECT -188.935 2.115 -188.765 2.285 ;
        RECT -184.875 2.115 -184.705 2.285 ;
        RECT -179.015 2.115 -178.845 2.285 ;
        RECT -174.955 2.115 -174.785 2.285 ;
        RECT -169.095 2.115 -168.925 2.285 ;
        RECT -165.035 2.115 -164.865 2.285 ;
        RECT -159.175 2.115 -159.005 2.285 ;
        RECT -155.115 2.115 -154.945 2.285 ;
        RECT -149.255 2.115 -149.085 2.285 ;
        RECT -145.195 2.115 -145.025 2.285 ;
        RECT -139.335 2.115 -139.165 2.285 ;
        RECT -135.275 2.115 -135.105 2.285 ;
        RECT -129.415 2.115 -129.245 2.285 ;
        RECT -125.355 2.115 -125.185 2.285 ;
        RECT -119.495 2.115 -119.325 2.285 ;
        RECT -115.435 2.115 -115.265 2.285 ;
        RECT -109.575 2.115 -109.405 2.285 ;
        RECT -105.515 2.115 -105.345 2.285 ;
        RECT -99.655 2.115 -99.485 2.285 ;
        RECT -95.595 2.115 -95.425 2.285 ;
        RECT -89.735 2.115 -89.565 2.285 ;
        RECT -85.675 2.115 -85.505 2.285 ;
        RECT -79.815 2.115 -79.645 2.285 ;
        RECT -75.755 2.115 -75.585 2.285 ;
        RECT -69.895 2.115 -69.725 2.285 ;
        RECT -65.835 2.115 -65.665 2.285 ;
        RECT -59.975 2.115 -59.805 2.285 ;
        RECT -55.915 2.115 -55.745 2.285 ;
        RECT -50.055 2.115 -49.885 2.285 ;
        RECT -45.995 2.115 -45.825 2.285 ;
        RECT -40.135 2.115 -39.965 2.285 ;
        RECT -36.075 2.115 -35.905 2.285 ;
        RECT -30.215 2.115 -30.045 2.285 ;
        RECT -26.155 2.115 -25.985 2.285 ;
        RECT -20.295 2.115 -20.125 2.285 ;
        RECT -16.235 2.115 -16.065 2.285 ;
        RECT -10.375 2.115 -10.205 2.285 ;
        RECT -6.315 2.115 -6.145 2.285 ;
        RECT -0.455 2.115 -0.285 2.285 ;
        RECT 3.605 2.115 3.775 2.285 ;
        RECT 9.465 2.115 9.635 2.285 ;
        RECT 13.525 2.115 13.695 2.285 ;
        RECT 19.385 2.115 19.555 2.285 ;
        RECT 23.445 2.115 23.615 2.285 ;
        RECT 24.605 2.155 24.775 2.325 ;
        RECT 24.605 1.695 24.775 1.865 ;
        RECT -289.765 1.245 -289.595 1.415 ;
        RECT -289.295 1.235 -289.125 1.405 ;
        RECT -284.810 1.265 -284.640 1.435 ;
        RECT -283.445 1.265 -283.275 1.435 ;
        RECT -274.890 1.265 -274.720 1.435 ;
        RECT -273.525 1.265 -273.355 1.435 ;
        RECT -264.970 1.265 -264.800 1.435 ;
        RECT -263.605 1.265 -263.435 1.435 ;
        RECT -255.050 1.265 -254.880 1.435 ;
        RECT -253.685 1.265 -253.515 1.435 ;
        RECT -245.130 1.265 -244.960 1.435 ;
        RECT -243.765 1.265 -243.595 1.435 ;
        RECT -235.210 1.265 -235.040 1.435 ;
        RECT -233.845 1.265 -233.675 1.435 ;
        RECT -225.290 1.265 -225.120 1.435 ;
        RECT -223.925 1.265 -223.755 1.435 ;
        RECT -215.370 1.265 -215.200 1.435 ;
        RECT -214.005 1.265 -213.835 1.435 ;
        RECT -205.450 1.265 -205.280 1.435 ;
        RECT -204.085 1.265 -203.915 1.435 ;
        RECT -195.530 1.265 -195.360 1.435 ;
        RECT -194.165 1.265 -193.995 1.435 ;
        RECT -185.610 1.265 -185.440 1.435 ;
        RECT -184.245 1.265 -184.075 1.435 ;
        RECT -175.690 1.265 -175.520 1.435 ;
        RECT -174.325 1.265 -174.155 1.435 ;
        RECT -165.770 1.265 -165.600 1.435 ;
        RECT -164.405 1.265 -164.235 1.435 ;
        RECT -155.850 1.265 -155.680 1.435 ;
        RECT -154.485 1.265 -154.315 1.435 ;
        RECT -145.930 1.265 -145.760 1.435 ;
        RECT -144.565 1.265 -144.395 1.435 ;
        RECT -136.010 1.265 -135.840 1.435 ;
        RECT -134.645 1.265 -134.475 1.435 ;
        RECT -126.090 1.265 -125.920 1.435 ;
        RECT -124.725 1.265 -124.555 1.435 ;
        RECT -116.170 1.265 -116.000 1.435 ;
        RECT -114.805 1.265 -114.635 1.435 ;
        RECT -106.250 1.265 -106.080 1.435 ;
        RECT -104.885 1.265 -104.715 1.435 ;
        RECT -96.330 1.265 -96.160 1.435 ;
        RECT -94.965 1.265 -94.795 1.435 ;
        RECT -86.410 1.265 -86.240 1.435 ;
        RECT -85.045 1.265 -84.875 1.435 ;
        RECT -76.490 1.265 -76.320 1.435 ;
        RECT -75.125 1.265 -74.955 1.435 ;
        RECT -66.570 1.265 -66.400 1.435 ;
        RECT -65.205 1.265 -65.035 1.435 ;
        RECT -56.650 1.265 -56.480 1.435 ;
        RECT -55.285 1.265 -55.115 1.435 ;
        RECT -46.730 1.265 -46.560 1.435 ;
        RECT -45.365 1.265 -45.195 1.435 ;
        RECT -36.810 1.265 -36.640 1.435 ;
        RECT -35.445 1.265 -35.275 1.435 ;
        RECT -26.890 1.265 -26.720 1.435 ;
        RECT -25.525 1.265 -25.355 1.435 ;
        RECT -16.970 1.265 -16.800 1.435 ;
        RECT -15.605 1.265 -15.435 1.435 ;
        RECT -7.050 1.265 -6.880 1.435 ;
        RECT -5.685 1.265 -5.515 1.435 ;
        RECT 2.870 1.265 3.040 1.435 ;
        RECT 4.235 1.265 4.405 1.435 ;
        RECT 12.790 1.265 12.960 1.435 ;
        RECT 14.155 1.265 14.325 1.435 ;
        RECT 22.710 1.265 22.880 1.435 ;
        RECT 24.075 1.265 24.245 1.435 ;
        RECT 24.605 1.235 24.775 1.405 ;
        RECT 25.075 1.245 25.245 1.415 ;
        RECT -289.305 -86.240 -289.135 -86.070 ;
        RECT -288.835 -86.235 -288.665 -86.065 ;
        RECT -288.010 -86.265 -287.840 -86.095 ;
        RECT -286.645 -86.265 -286.475 -86.095 ;
        RECT -278.090 -86.265 -277.920 -86.095 ;
        RECT -276.725 -86.265 -276.555 -86.095 ;
        RECT -268.170 -86.265 -268.000 -86.095 ;
        RECT -266.805 -86.265 -266.635 -86.095 ;
        RECT -258.250 -86.265 -258.080 -86.095 ;
        RECT -256.885 -86.265 -256.715 -86.095 ;
        RECT -248.330 -86.265 -248.160 -86.095 ;
        RECT -246.965 -86.265 -246.795 -86.095 ;
        RECT -238.410 -86.265 -238.240 -86.095 ;
        RECT -237.045 -86.265 -236.875 -86.095 ;
        RECT -228.490 -86.265 -228.320 -86.095 ;
        RECT -227.125 -86.265 -226.955 -86.095 ;
        RECT -218.570 -86.265 -218.400 -86.095 ;
        RECT -217.205 -86.265 -217.035 -86.095 ;
        RECT -208.650 -86.265 -208.480 -86.095 ;
        RECT -207.285 -86.265 -207.115 -86.095 ;
        RECT -198.730 -86.265 -198.560 -86.095 ;
        RECT -197.365 -86.265 -197.195 -86.095 ;
        RECT -188.810 -86.265 -188.640 -86.095 ;
        RECT -187.445 -86.265 -187.275 -86.095 ;
        RECT -178.890 -86.265 -178.720 -86.095 ;
        RECT -177.525 -86.265 -177.355 -86.095 ;
        RECT -168.970 -86.265 -168.800 -86.095 ;
        RECT -167.605 -86.265 -167.435 -86.095 ;
        RECT -159.050 -86.265 -158.880 -86.095 ;
        RECT -157.685 -86.265 -157.515 -86.095 ;
        RECT -149.130 -86.265 -148.960 -86.095 ;
        RECT -147.765 -86.265 -147.595 -86.095 ;
        RECT -139.210 -86.265 -139.040 -86.095 ;
        RECT -137.845 -86.265 -137.675 -86.095 ;
        RECT -129.290 -86.265 -129.120 -86.095 ;
        RECT -127.925 -86.265 -127.755 -86.095 ;
        RECT -119.370 -86.265 -119.200 -86.095 ;
        RECT -118.005 -86.265 -117.835 -86.095 ;
        RECT -109.450 -86.265 -109.280 -86.095 ;
        RECT -108.085 -86.265 -107.915 -86.095 ;
        RECT -99.530 -86.265 -99.360 -86.095 ;
        RECT -98.165 -86.265 -97.995 -86.095 ;
        RECT -89.610 -86.265 -89.440 -86.095 ;
        RECT -88.245 -86.265 -88.075 -86.095 ;
        RECT -79.690 -86.265 -79.520 -86.095 ;
        RECT -78.325 -86.265 -78.155 -86.095 ;
        RECT -69.770 -86.265 -69.600 -86.095 ;
        RECT -68.405 -86.265 -68.235 -86.095 ;
        RECT -59.850 -86.265 -59.680 -86.095 ;
        RECT -58.485 -86.265 -58.315 -86.095 ;
        RECT -49.930 -86.265 -49.760 -86.095 ;
        RECT -48.565 -86.265 -48.395 -86.095 ;
        RECT -40.010 -86.265 -39.840 -86.095 ;
        RECT -38.645 -86.265 -38.475 -86.095 ;
        RECT -30.090 -86.265 -29.920 -86.095 ;
        RECT -28.725 -86.265 -28.555 -86.095 ;
        RECT -20.170 -86.265 -20.000 -86.095 ;
        RECT -18.805 -86.265 -18.635 -86.095 ;
        RECT -10.250 -86.265 -10.080 -86.095 ;
        RECT -8.885 -86.265 -8.715 -86.095 ;
        RECT -0.330 -86.265 -0.160 -86.095 ;
        RECT 1.035 -86.265 1.205 -86.095 ;
        RECT 9.590 -86.265 9.760 -86.095 ;
        RECT 10.955 -86.265 11.125 -86.095 ;
        RECT 19.510 -86.265 19.680 -86.095 ;
        RECT 20.875 -86.265 21.045 -86.095 ;
        RECT -288.835 -86.695 -288.665 -86.525 ;
        RECT -288.835 -87.155 -288.665 -86.985 ;
        RECT -287.275 -87.115 -287.105 -86.945 ;
        RECT -281.415 -87.115 -281.245 -86.945 ;
        RECT -277.355 -87.115 -277.185 -86.945 ;
        RECT -271.495 -87.115 -271.325 -86.945 ;
        RECT -267.435 -87.115 -267.265 -86.945 ;
        RECT -261.575 -87.115 -261.405 -86.945 ;
        RECT -257.515 -87.115 -257.345 -86.945 ;
        RECT -251.655 -87.115 -251.485 -86.945 ;
        RECT -247.595 -87.115 -247.425 -86.945 ;
        RECT -241.735 -87.115 -241.565 -86.945 ;
        RECT -237.675 -87.115 -237.505 -86.945 ;
        RECT -231.815 -87.115 -231.645 -86.945 ;
        RECT -227.755 -87.115 -227.585 -86.945 ;
        RECT -221.895 -87.115 -221.725 -86.945 ;
        RECT -217.835 -87.115 -217.665 -86.945 ;
        RECT -211.975 -87.115 -211.805 -86.945 ;
        RECT -207.915 -87.115 -207.745 -86.945 ;
        RECT -202.055 -87.115 -201.885 -86.945 ;
        RECT -197.995 -87.115 -197.825 -86.945 ;
        RECT -192.135 -87.115 -191.965 -86.945 ;
        RECT -188.075 -87.115 -187.905 -86.945 ;
        RECT -182.215 -87.115 -182.045 -86.945 ;
        RECT -178.155 -87.115 -177.985 -86.945 ;
        RECT -172.295 -87.115 -172.125 -86.945 ;
        RECT -168.235 -87.115 -168.065 -86.945 ;
        RECT -162.375 -87.115 -162.205 -86.945 ;
        RECT -158.315 -87.115 -158.145 -86.945 ;
        RECT -152.455 -87.115 -152.285 -86.945 ;
        RECT -148.395 -87.115 -148.225 -86.945 ;
        RECT -142.535 -87.115 -142.365 -86.945 ;
        RECT -138.475 -87.115 -138.305 -86.945 ;
        RECT -132.615 -87.115 -132.445 -86.945 ;
        RECT -128.555 -87.115 -128.385 -86.945 ;
        RECT -122.695 -87.115 -122.525 -86.945 ;
        RECT -118.635 -87.115 -118.465 -86.945 ;
        RECT -112.775 -87.115 -112.605 -86.945 ;
        RECT -108.715 -87.115 -108.545 -86.945 ;
        RECT -102.855 -87.115 -102.685 -86.945 ;
        RECT -98.795 -87.115 -98.625 -86.945 ;
        RECT -92.935 -87.115 -92.765 -86.945 ;
        RECT -88.875 -87.115 -88.705 -86.945 ;
        RECT -83.015 -87.115 -82.845 -86.945 ;
        RECT -78.955 -87.115 -78.785 -86.945 ;
        RECT -73.095 -87.115 -72.925 -86.945 ;
        RECT -69.035 -87.115 -68.865 -86.945 ;
        RECT -63.175 -87.115 -63.005 -86.945 ;
        RECT -59.115 -87.115 -58.945 -86.945 ;
        RECT -53.255 -87.115 -53.085 -86.945 ;
        RECT -49.195 -87.115 -49.025 -86.945 ;
        RECT -43.335 -87.115 -43.165 -86.945 ;
        RECT -39.275 -87.115 -39.105 -86.945 ;
        RECT -33.415 -87.115 -33.245 -86.945 ;
        RECT -29.355 -87.115 -29.185 -86.945 ;
        RECT -23.495 -87.115 -23.325 -86.945 ;
        RECT -19.435 -87.115 -19.265 -86.945 ;
        RECT -13.575 -87.115 -13.405 -86.945 ;
        RECT -9.515 -87.115 -9.345 -86.945 ;
        RECT -3.655 -87.115 -3.485 -86.945 ;
        RECT 0.405 -87.115 0.575 -86.945 ;
        RECT 6.265 -87.115 6.435 -86.945 ;
        RECT 10.325 -87.115 10.495 -86.945 ;
        RECT 16.185 -87.115 16.355 -86.945 ;
        RECT 20.245 -87.115 20.415 -86.945 ;
        RECT 26.105 -87.115 26.275 -86.945 ;
        RECT -289.305 -87.815 -289.135 -87.645 ;
        RECT -288.845 -87.815 -288.675 -87.645 ;
        RECT -288.385 -87.815 -288.215 -87.645 ;
        RECT -287.925 -87.815 -287.755 -87.645 ;
        RECT 26.755 -87.815 26.925 -87.645 ;
        RECT 27.215 -87.815 27.385 -87.645 ;
        RECT 27.675 -87.815 27.845 -87.645 ;
        RECT 28.135 -87.815 28.305 -87.645 ;
        RECT -287.955 -88.535 -287.785 -88.365 ;
        RECT -287.970 -88.975 -287.800 -88.805 ;
        RECT -280.735 -88.535 -280.565 -88.365 ;
        RECT -285.680 -89.375 -285.510 -89.205 ;
        RECT -285.695 -89.815 -285.525 -89.645 ;
        RECT -280.720 -88.975 -280.550 -88.805 ;
        RECT -283.010 -89.375 -282.840 -89.205 ;
        RECT -278.035 -88.535 -277.865 -88.365 ;
        RECT -278.050 -88.975 -277.880 -88.805 ;
        RECT -270.815 -88.535 -270.645 -88.365 ;
        RECT -282.995 -89.815 -282.825 -89.645 ;
        RECT -275.760 -89.375 -275.590 -89.205 ;
        RECT -275.775 -89.815 -275.605 -89.645 ;
        RECT -270.800 -88.975 -270.630 -88.805 ;
        RECT -273.090 -89.375 -272.920 -89.205 ;
        RECT -268.115 -88.535 -267.945 -88.365 ;
        RECT -268.130 -88.975 -267.960 -88.805 ;
        RECT -260.895 -88.535 -260.725 -88.365 ;
        RECT -273.075 -89.815 -272.905 -89.645 ;
        RECT -265.840 -89.375 -265.670 -89.205 ;
        RECT -265.855 -89.815 -265.685 -89.645 ;
        RECT -260.880 -88.975 -260.710 -88.805 ;
        RECT -263.170 -89.375 -263.000 -89.205 ;
        RECT -258.195 -88.535 -258.025 -88.365 ;
        RECT -258.210 -88.975 -258.040 -88.805 ;
        RECT -250.975 -88.535 -250.805 -88.365 ;
        RECT -263.155 -89.815 -262.985 -89.645 ;
        RECT -255.920 -89.375 -255.750 -89.205 ;
        RECT -255.935 -89.815 -255.765 -89.645 ;
        RECT -250.960 -88.975 -250.790 -88.805 ;
        RECT -253.250 -89.375 -253.080 -89.205 ;
        RECT -248.275 -88.535 -248.105 -88.365 ;
        RECT -248.290 -88.975 -248.120 -88.805 ;
        RECT -241.055 -88.535 -240.885 -88.365 ;
        RECT -253.235 -89.815 -253.065 -89.645 ;
        RECT -246.000 -89.375 -245.830 -89.205 ;
        RECT -246.015 -89.815 -245.845 -89.645 ;
        RECT -241.040 -88.975 -240.870 -88.805 ;
        RECT -243.330 -89.375 -243.160 -89.205 ;
        RECT -238.355 -88.535 -238.185 -88.365 ;
        RECT -238.370 -88.975 -238.200 -88.805 ;
        RECT -231.135 -88.535 -230.965 -88.365 ;
        RECT -243.315 -89.815 -243.145 -89.645 ;
        RECT -236.080 -89.375 -235.910 -89.205 ;
        RECT -236.095 -89.815 -235.925 -89.645 ;
        RECT -231.120 -88.975 -230.950 -88.805 ;
        RECT -233.410 -89.375 -233.240 -89.205 ;
        RECT -228.435 -88.535 -228.265 -88.365 ;
        RECT -228.450 -88.975 -228.280 -88.805 ;
        RECT -221.215 -88.535 -221.045 -88.365 ;
        RECT -233.395 -89.815 -233.225 -89.645 ;
        RECT -226.160 -89.375 -225.990 -89.205 ;
        RECT -226.175 -89.815 -226.005 -89.645 ;
        RECT -221.200 -88.975 -221.030 -88.805 ;
        RECT -223.490 -89.375 -223.320 -89.205 ;
        RECT -218.515 -88.535 -218.345 -88.365 ;
        RECT -218.530 -88.975 -218.360 -88.805 ;
        RECT -211.295 -88.535 -211.125 -88.365 ;
        RECT -223.475 -89.815 -223.305 -89.645 ;
        RECT -216.240 -89.375 -216.070 -89.205 ;
        RECT -216.255 -89.815 -216.085 -89.645 ;
        RECT -211.280 -88.975 -211.110 -88.805 ;
        RECT -213.570 -89.375 -213.400 -89.205 ;
        RECT -208.595 -88.535 -208.425 -88.365 ;
        RECT -208.610 -88.975 -208.440 -88.805 ;
        RECT -201.375 -88.535 -201.205 -88.365 ;
        RECT -213.555 -89.815 -213.385 -89.645 ;
        RECT -206.320 -89.375 -206.150 -89.205 ;
        RECT -206.335 -89.815 -206.165 -89.645 ;
        RECT -201.360 -88.975 -201.190 -88.805 ;
        RECT -203.650 -89.375 -203.480 -89.205 ;
        RECT -198.675 -88.535 -198.505 -88.365 ;
        RECT -198.690 -88.975 -198.520 -88.805 ;
        RECT -191.455 -88.535 -191.285 -88.365 ;
        RECT -203.635 -89.815 -203.465 -89.645 ;
        RECT -196.400 -89.375 -196.230 -89.205 ;
        RECT -196.415 -89.815 -196.245 -89.645 ;
        RECT -191.440 -88.975 -191.270 -88.805 ;
        RECT -193.730 -89.375 -193.560 -89.205 ;
        RECT -188.755 -88.535 -188.585 -88.365 ;
        RECT -188.770 -88.975 -188.600 -88.805 ;
        RECT -181.535 -88.535 -181.365 -88.365 ;
        RECT -193.715 -89.815 -193.545 -89.645 ;
        RECT -186.480 -89.375 -186.310 -89.205 ;
        RECT -186.495 -89.815 -186.325 -89.645 ;
        RECT -181.520 -88.975 -181.350 -88.805 ;
        RECT -183.810 -89.375 -183.640 -89.205 ;
        RECT -178.835 -88.535 -178.665 -88.365 ;
        RECT -178.850 -88.975 -178.680 -88.805 ;
        RECT -171.615 -88.535 -171.445 -88.365 ;
        RECT -183.795 -89.815 -183.625 -89.645 ;
        RECT -176.560 -89.375 -176.390 -89.205 ;
        RECT -176.575 -89.815 -176.405 -89.645 ;
        RECT -171.600 -88.975 -171.430 -88.805 ;
        RECT -173.890 -89.375 -173.720 -89.205 ;
        RECT -168.915 -88.535 -168.745 -88.365 ;
        RECT -168.930 -88.975 -168.760 -88.805 ;
        RECT -161.695 -88.535 -161.525 -88.365 ;
        RECT -173.875 -89.815 -173.705 -89.645 ;
        RECT -166.640 -89.375 -166.470 -89.205 ;
        RECT -166.655 -89.815 -166.485 -89.645 ;
        RECT -161.680 -88.975 -161.510 -88.805 ;
        RECT -163.970 -89.375 -163.800 -89.205 ;
        RECT -158.995 -88.535 -158.825 -88.365 ;
        RECT -159.010 -88.975 -158.840 -88.805 ;
        RECT -151.775 -88.535 -151.605 -88.365 ;
        RECT -163.955 -89.815 -163.785 -89.645 ;
        RECT -156.720 -89.375 -156.550 -89.205 ;
        RECT -156.735 -89.815 -156.565 -89.645 ;
        RECT -151.760 -88.975 -151.590 -88.805 ;
        RECT -154.050 -89.375 -153.880 -89.205 ;
        RECT -149.075 -88.535 -148.905 -88.365 ;
        RECT -149.090 -88.975 -148.920 -88.805 ;
        RECT -141.855 -88.535 -141.685 -88.365 ;
        RECT -154.035 -89.815 -153.865 -89.645 ;
        RECT -146.800 -89.375 -146.630 -89.205 ;
        RECT -146.815 -89.815 -146.645 -89.645 ;
        RECT -141.840 -88.975 -141.670 -88.805 ;
        RECT -144.130 -89.375 -143.960 -89.205 ;
        RECT -139.155 -88.535 -138.985 -88.365 ;
        RECT -139.170 -88.975 -139.000 -88.805 ;
        RECT -131.935 -88.535 -131.765 -88.365 ;
        RECT -144.115 -89.815 -143.945 -89.645 ;
        RECT -136.880 -89.375 -136.710 -89.205 ;
        RECT -136.895 -89.815 -136.725 -89.645 ;
        RECT -131.920 -88.975 -131.750 -88.805 ;
        RECT -134.210 -89.375 -134.040 -89.205 ;
        RECT -129.235 -88.535 -129.065 -88.365 ;
        RECT -129.250 -88.975 -129.080 -88.805 ;
        RECT -122.015 -88.535 -121.845 -88.365 ;
        RECT -134.195 -89.815 -134.025 -89.645 ;
        RECT -126.960 -89.375 -126.790 -89.205 ;
        RECT -126.975 -89.815 -126.805 -89.645 ;
        RECT -122.000 -88.975 -121.830 -88.805 ;
        RECT -124.290 -89.375 -124.120 -89.205 ;
        RECT -119.315 -88.535 -119.145 -88.365 ;
        RECT -119.330 -88.975 -119.160 -88.805 ;
        RECT -112.095 -88.535 -111.925 -88.365 ;
        RECT -124.275 -89.815 -124.105 -89.645 ;
        RECT -117.040 -89.375 -116.870 -89.205 ;
        RECT -117.055 -89.815 -116.885 -89.645 ;
        RECT -112.080 -88.975 -111.910 -88.805 ;
        RECT -114.370 -89.375 -114.200 -89.205 ;
        RECT -109.395 -88.535 -109.225 -88.365 ;
        RECT -109.410 -88.975 -109.240 -88.805 ;
        RECT -102.175 -88.535 -102.005 -88.365 ;
        RECT -114.355 -89.815 -114.185 -89.645 ;
        RECT -107.120 -89.375 -106.950 -89.205 ;
        RECT -107.135 -89.815 -106.965 -89.645 ;
        RECT -102.160 -88.975 -101.990 -88.805 ;
        RECT -104.450 -89.375 -104.280 -89.205 ;
        RECT -99.475 -88.535 -99.305 -88.365 ;
        RECT -99.490 -88.975 -99.320 -88.805 ;
        RECT -92.255 -88.535 -92.085 -88.365 ;
        RECT -104.435 -89.815 -104.265 -89.645 ;
        RECT -97.200 -89.375 -97.030 -89.205 ;
        RECT -97.215 -89.815 -97.045 -89.645 ;
        RECT -92.240 -88.975 -92.070 -88.805 ;
        RECT -94.530 -89.375 -94.360 -89.205 ;
        RECT -89.555 -88.535 -89.385 -88.365 ;
        RECT -89.570 -88.975 -89.400 -88.805 ;
        RECT -82.335 -88.535 -82.165 -88.365 ;
        RECT -94.515 -89.815 -94.345 -89.645 ;
        RECT -87.280 -89.375 -87.110 -89.205 ;
        RECT -87.295 -89.815 -87.125 -89.645 ;
        RECT -82.320 -88.975 -82.150 -88.805 ;
        RECT -84.610 -89.375 -84.440 -89.205 ;
        RECT -79.635 -88.535 -79.465 -88.365 ;
        RECT -79.650 -88.975 -79.480 -88.805 ;
        RECT -72.415 -88.535 -72.245 -88.365 ;
        RECT -84.595 -89.815 -84.425 -89.645 ;
        RECT -77.360 -89.375 -77.190 -89.205 ;
        RECT -77.375 -89.815 -77.205 -89.645 ;
        RECT -72.400 -88.975 -72.230 -88.805 ;
        RECT -74.690 -89.375 -74.520 -89.205 ;
        RECT -69.715 -88.535 -69.545 -88.365 ;
        RECT -69.730 -88.975 -69.560 -88.805 ;
        RECT -62.495 -88.535 -62.325 -88.365 ;
        RECT -74.675 -89.815 -74.505 -89.645 ;
        RECT -67.440 -89.375 -67.270 -89.205 ;
        RECT -67.455 -89.815 -67.285 -89.645 ;
        RECT -62.480 -88.975 -62.310 -88.805 ;
        RECT -64.770 -89.375 -64.600 -89.205 ;
        RECT -59.795 -88.535 -59.625 -88.365 ;
        RECT -59.810 -88.975 -59.640 -88.805 ;
        RECT -52.575 -88.535 -52.405 -88.365 ;
        RECT -64.755 -89.815 -64.585 -89.645 ;
        RECT -57.520 -89.375 -57.350 -89.205 ;
        RECT -57.535 -89.815 -57.365 -89.645 ;
        RECT -52.560 -88.975 -52.390 -88.805 ;
        RECT -54.850 -89.375 -54.680 -89.205 ;
        RECT -49.875 -88.535 -49.705 -88.365 ;
        RECT -49.890 -88.975 -49.720 -88.805 ;
        RECT -42.655 -88.535 -42.485 -88.365 ;
        RECT -54.835 -89.815 -54.665 -89.645 ;
        RECT -47.600 -89.375 -47.430 -89.205 ;
        RECT -47.615 -89.815 -47.445 -89.645 ;
        RECT -42.640 -88.975 -42.470 -88.805 ;
        RECT -44.930 -89.375 -44.760 -89.205 ;
        RECT -39.955 -88.535 -39.785 -88.365 ;
        RECT -39.970 -88.975 -39.800 -88.805 ;
        RECT -32.735 -88.535 -32.565 -88.365 ;
        RECT -44.915 -89.815 -44.745 -89.645 ;
        RECT -37.680 -89.375 -37.510 -89.205 ;
        RECT -37.695 -89.815 -37.525 -89.645 ;
        RECT -32.720 -88.975 -32.550 -88.805 ;
        RECT -35.010 -89.375 -34.840 -89.205 ;
        RECT -30.035 -88.535 -29.865 -88.365 ;
        RECT -30.050 -88.975 -29.880 -88.805 ;
        RECT -22.815 -88.535 -22.645 -88.365 ;
        RECT -34.995 -89.815 -34.825 -89.645 ;
        RECT -27.760 -89.375 -27.590 -89.205 ;
        RECT -27.775 -89.815 -27.605 -89.645 ;
        RECT -22.800 -88.975 -22.630 -88.805 ;
        RECT -25.090 -89.375 -24.920 -89.205 ;
        RECT -20.115 -88.535 -19.945 -88.365 ;
        RECT -20.130 -88.975 -19.960 -88.805 ;
        RECT -12.895 -88.535 -12.725 -88.365 ;
        RECT -25.075 -89.815 -24.905 -89.645 ;
        RECT -17.840 -89.375 -17.670 -89.205 ;
        RECT -17.855 -89.815 -17.685 -89.645 ;
        RECT -12.880 -88.975 -12.710 -88.805 ;
        RECT -15.170 -89.375 -15.000 -89.205 ;
        RECT -10.195 -88.535 -10.025 -88.365 ;
        RECT -10.210 -88.975 -10.040 -88.805 ;
        RECT -2.975 -88.535 -2.805 -88.365 ;
        RECT -15.155 -89.815 -14.985 -89.645 ;
        RECT -7.920 -89.375 -7.750 -89.205 ;
        RECT -7.935 -89.815 -7.765 -89.645 ;
        RECT -2.960 -88.975 -2.790 -88.805 ;
        RECT -5.250 -89.375 -5.080 -89.205 ;
        RECT -0.275 -88.535 -0.105 -88.365 ;
        RECT -0.290 -88.975 -0.120 -88.805 ;
        RECT 6.945 -88.535 7.115 -88.365 ;
        RECT -5.235 -89.815 -5.065 -89.645 ;
        RECT 2.000 -89.375 2.170 -89.205 ;
        RECT 1.985 -89.815 2.155 -89.645 ;
        RECT 6.960 -88.975 7.130 -88.805 ;
        RECT 4.670 -89.375 4.840 -89.205 ;
        RECT 9.645 -88.535 9.815 -88.365 ;
        RECT 9.630 -88.975 9.800 -88.805 ;
        RECT 16.865 -88.535 17.035 -88.365 ;
        RECT 4.685 -89.815 4.855 -89.645 ;
        RECT 11.920 -89.375 12.090 -89.205 ;
        RECT 11.905 -89.815 12.075 -89.645 ;
        RECT 16.880 -88.975 17.050 -88.805 ;
        RECT 14.590 -89.375 14.760 -89.205 ;
        RECT 19.565 -88.535 19.735 -88.365 ;
        RECT 19.550 -88.975 19.720 -88.805 ;
        RECT 26.785 -88.535 26.955 -88.365 ;
        RECT 14.605 -89.815 14.775 -89.645 ;
        RECT 21.840 -89.375 22.010 -89.205 ;
        RECT 21.825 -89.815 21.995 -89.645 ;
        RECT 26.800 -88.975 26.970 -88.805 ;
        RECT 24.510 -89.375 24.680 -89.205 ;
        RECT 24.525 -89.815 24.695 -89.645 ;
        RECT -289.305 -90.535 -289.135 -90.365 ;
        RECT -288.845 -90.535 -288.675 -90.365 ;
        RECT -288.385 -90.535 -288.215 -90.365 ;
        RECT -287.925 -90.535 -287.755 -90.365 ;
        RECT -287.535 -91.195 -287.365 -91.025 ;
        RECT -287.535 -91.655 -287.365 -91.485 ;
        RECT -286.375 -91.235 -286.205 -91.065 ;
        RECT -282.315 -91.235 -282.145 -91.065 ;
        RECT -276.455 -91.235 -276.285 -91.065 ;
        RECT -272.395 -91.235 -272.225 -91.065 ;
        RECT -266.535 -91.235 -266.365 -91.065 ;
        RECT -262.475 -91.235 -262.305 -91.065 ;
        RECT -256.615 -91.235 -256.445 -91.065 ;
        RECT -252.555 -91.235 -252.385 -91.065 ;
        RECT -246.695 -91.235 -246.525 -91.065 ;
        RECT -242.635 -91.235 -242.465 -91.065 ;
        RECT -236.775 -91.235 -236.605 -91.065 ;
        RECT -232.715 -91.235 -232.545 -91.065 ;
        RECT -226.855 -91.235 -226.685 -91.065 ;
        RECT -222.795 -91.235 -222.625 -91.065 ;
        RECT -216.935 -91.235 -216.765 -91.065 ;
        RECT -212.875 -91.235 -212.705 -91.065 ;
        RECT -207.015 -91.235 -206.845 -91.065 ;
        RECT -202.955 -91.235 -202.785 -91.065 ;
        RECT -197.095 -91.235 -196.925 -91.065 ;
        RECT -193.035 -91.235 -192.865 -91.065 ;
        RECT -187.175 -91.235 -187.005 -91.065 ;
        RECT -183.115 -91.235 -182.945 -91.065 ;
        RECT -177.255 -91.235 -177.085 -91.065 ;
        RECT -173.195 -91.235 -173.025 -91.065 ;
        RECT -167.335 -91.235 -167.165 -91.065 ;
        RECT -163.275 -91.235 -163.105 -91.065 ;
        RECT -157.415 -91.235 -157.245 -91.065 ;
        RECT -153.355 -91.235 -153.185 -91.065 ;
        RECT -147.495 -91.235 -147.325 -91.065 ;
        RECT -143.435 -91.235 -143.265 -91.065 ;
        RECT -137.575 -91.235 -137.405 -91.065 ;
        RECT -133.515 -91.235 -133.345 -91.065 ;
        RECT -127.655 -91.235 -127.485 -91.065 ;
        RECT -123.595 -91.235 -123.425 -91.065 ;
        RECT -117.735 -91.235 -117.565 -91.065 ;
        RECT -113.675 -91.235 -113.505 -91.065 ;
        RECT -107.815 -91.235 -107.645 -91.065 ;
        RECT -103.755 -91.235 -103.585 -91.065 ;
        RECT -97.895 -91.235 -97.725 -91.065 ;
        RECT -93.835 -91.235 -93.665 -91.065 ;
        RECT -87.975 -91.235 -87.805 -91.065 ;
        RECT -83.915 -91.235 -83.745 -91.065 ;
        RECT -78.055 -91.235 -77.885 -91.065 ;
        RECT -73.995 -91.235 -73.825 -91.065 ;
        RECT -68.135 -91.235 -67.965 -91.065 ;
        RECT -64.075 -91.235 -63.905 -91.065 ;
        RECT -58.215 -91.235 -58.045 -91.065 ;
        RECT -54.155 -91.235 -53.985 -91.065 ;
        RECT -48.295 -91.235 -48.125 -91.065 ;
        RECT -44.235 -91.235 -44.065 -91.065 ;
        RECT -38.375 -91.235 -38.205 -91.065 ;
        RECT -34.315 -91.235 -34.145 -91.065 ;
        RECT -28.455 -91.235 -28.285 -91.065 ;
        RECT -24.395 -91.235 -24.225 -91.065 ;
        RECT -18.535 -91.235 -18.365 -91.065 ;
        RECT -14.475 -91.235 -14.305 -91.065 ;
        RECT -8.615 -91.235 -8.445 -91.065 ;
        RECT -4.555 -91.235 -4.385 -91.065 ;
        RECT 1.305 -91.235 1.475 -91.065 ;
        RECT 5.365 -91.235 5.535 -91.065 ;
        RECT 11.225 -91.235 11.395 -91.065 ;
        RECT 15.285 -91.235 15.455 -91.065 ;
        RECT 21.145 -91.235 21.315 -91.065 ;
        RECT 25.205 -91.235 25.375 -91.065 ;
        RECT 26.365 -91.195 26.535 -91.025 ;
        RECT 26.365 -91.655 26.535 -91.485 ;
        RECT -288.005 -92.105 -287.835 -91.935 ;
        RECT -287.535 -92.115 -287.365 -91.945 ;
        RECT -283.050 -92.085 -282.880 -91.915 ;
        RECT -281.685 -92.085 -281.515 -91.915 ;
        RECT -273.130 -92.085 -272.960 -91.915 ;
        RECT -271.765 -92.085 -271.595 -91.915 ;
        RECT -263.210 -92.085 -263.040 -91.915 ;
        RECT -261.845 -92.085 -261.675 -91.915 ;
        RECT -253.290 -92.085 -253.120 -91.915 ;
        RECT -251.925 -92.085 -251.755 -91.915 ;
        RECT -243.370 -92.085 -243.200 -91.915 ;
        RECT -242.005 -92.085 -241.835 -91.915 ;
        RECT -233.450 -92.085 -233.280 -91.915 ;
        RECT -232.085 -92.085 -231.915 -91.915 ;
        RECT -223.530 -92.085 -223.360 -91.915 ;
        RECT -222.165 -92.085 -221.995 -91.915 ;
        RECT -213.610 -92.085 -213.440 -91.915 ;
        RECT -212.245 -92.085 -212.075 -91.915 ;
        RECT -203.690 -92.085 -203.520 -91.915 ;
        RECT -202.325 -92.085 -202.155 -91.915 ;
        RECT -193.770 -92.085 -193.600 -91.915 ;
        RECT -192.405 -92.085 -192.235 -91.915 ;
        RECT -183.850 -92.085 -183.680 -91.915 ;
        RECT -182.485 -92.085 -182.315 -91.915 ;
        RECT -173.930 -92.085 -173.760 -91.915 ;
        RECT -172.565 -92.085 -172.395 -91.915 ;
        RECT -164.010 -92.085 -163.840 -91.915 ;
        RECT -162.645 -92.085 -162.475 -91.915 ;
        RECT -154.090 -92.085 -153.920 -91.915 ;
        RECT -152.725 -92.085 -152.555 -91.915 ;
        RECT -144.170 -92.085 -144.000 -91.915 ;
        RECT -142.805 -92.085 -142.635 -91.915 ;
        RECT -134.250 -92.085 -134.080 -91.915 ;
        RECT -132.885 -92.085 -132.715 -91.915 ;
        RECT -124.330 -92.085 -124.160 -91.915 ;
        RECT -122.965 -92.085 -122.795 -91.915 ;
        RECT -114.410 -92.085 -114.240 -91.915 ;
        RECT -113.045 -92.085 -112.875 -91.915 ;
        RECT -104.490 -92.085 -104.320 -91.915 ;
        RECT -103.125 -92.085 -102.955 -91.915 ;
        RECT -94.570 -92.085 -94.400 -91.915 ;
        RECT -93.205 -92.085 -93.035 -91.915 ;
        RECT -84.650 -92.085 -84.480 -91.915 ;
        RECT -83.285 -92.085 -83.115 -91.915 ;
        RECT -74.730 -92.085 -74.560 -91.915 ;
        RECT -73.365 -92.085 -73.195 -91.915 ;
        RECT -64.810 -92.085 -64.640 -91.915 ;
        RECT -63.445 -92.085 -63.275 -91.915 ;
        RECT -54.890 -92.085 -54.720 -91.915 ;
        RECT -53.525 -92.085 -53.355 -91.915 ;
        RECT -44.970 -92.085 -44.800 -91.915 ;
        RECT -43.605 -92.085 -43.435 -91.915 ;
        RECT -35.050 -92.085 -34.880 -91.915 ;
        RECT -33.685 -92.085 -33.515 -91.915 ;
        RECT -25.130 -92.085 -24.960 -91.915 ;
        RECT -23.765 -92.085 -23.595 -91.915 ;
        RECT -15.210 -92.085 -15.040 -91.915 ;
        RECT -13.845 -92.085 -13.675 -91.915 ;
        RECT -5.290 -92.085 -5.120 -91.915 ;
        RECT -3.925 -92.085 -3.755 -91.915 ;
        RECT 4.630 -92.085 4.800 -91.915 ;
        RECT 5.995 -92.085 6.165 -91.915 ;
        RECT 14.550 -92.085 14.720 -91.915 ;
        RECT 15.915 -92.085 16.085 -91.915 ;
        RECT 24.470 -92.085 24.640 -91.915 ;
        RECT 25.835 -92.085 26.005 -91.915 ;
        RECT 26.365 -92.115 26.535 -91.945 ;
        RECT 26.835 -92.105 27.005 -91.935 ;
        RECT -289.055 -173.950 -288.885 -173.780 ;
        RECT -288.585 -173.945 -288.415 -173.775 ;
        RECT -287.760 -173.975 -287.590 -173.805 ;
        RECT -286.395 -173.975 -286.225 -173.805 ;
        RECT -277.840 -173.975 -277.670 -173.805 ;
        RECT -276.475 -173.975 -276.305 -173.805 ;
        RECT -267.920 -173.975 -267.750 -173.805 ;
        RECT -266.555 -173.975 -266.385 -173.805 ;
        RECT -258.000 -173.975 -257.830 -173.805 ;
        RECT -256.635 -173.975 -256.465 -173.805 ;
        RECT -248.080 -173.975 -247.910 -173.805 ;
        RECT -246.715 -173.975 -246.545 -173.805 ;
        RECT -238.160 -173.975 -237.990 -173.805 ;
        RECT -236.795 -173.975 -236.625 -173.805 ;
        RECT -228.240 -173.975 -228.070 -173.805 ;
        RECT -226.875 -173.975 -226.705 -173.805 ;
        RECT -218.320 -173.975 -218.150 -173.805 ;
        RECT -216.955 -173.975 -216.785 -173.805 ;
        RECT -208.400 -173.975 -208.230 -173.805 ;
        RECT -207.035 -173.975 -206.865 -173.805 ;
        RECT -198.480 -173.975 -198.310 -173.805 ;
        RECT -197.115 -173.975 -196.945 -173.805 ;
        RECT -188.560 -173.975 -188.390 -173.805 ;
        RECT -187.195 -173.975 -187.025 -173.805 ;
        RECT -178.640 -173.975 -178.470 -173.805 ;
        RECT -177.275 -173.975 -177.105 -173.805 ;
        RECT -168.720 -173.975 -168.550 -173.805 ;
        RECT -167.355 -173.975 -167.185 -173.805 ;
        RECT -158.800 -173.975 -158.630 -173.805 ;
        RECT -157.435 -173.975 -157.265 -173.805 ;
        RECT -148.880 -173.975 -148.710 -173.805 ;
        RECT -147.515 -173.975 -147.345 -173.805 ;
        RECT -138.960 -173.975 -138.790 -173.805 ;
        RECT -137.595 -173.975 -137.425 -173.805 ;
        RECT -129.040 -173.975 -128.870 -173.805 ;
        RECT -127.675 -173.975 -127.505 -173.805 ;
        RECT -119.120 -173.975 -118.950 -173.805 ;
        RECT -117.755 -173.975 -117.585 -173.805 ;
        RECT -109.200 -173.975 -109.030 -173.805 ;
        RECT -107.835 -173.975 -107.665 -173.805 ;
        RECT -99.280 -173.975 -99.110 -173.805 ;
        RECT -97.915 -173.975 -97.745 -173.805 ;
        RECT -89.360 -173.975 -89.190 -173.805 ;
        RECT -87.995 -173.975 -87.825 -173.805 ;
        RECT -79.440 -173.975 -79.270 -173.805 ;
        RECT -78.075 -173.975 -77.905 -173.805 ;
        RECT -69.520 -173.975 -69.350 -173.805 ;
        RECT -68.155 -173.975 -67.985 -173.805 ;
        RECT -59.600 -173.975 -59.430 -173.805 ;
        RECT -58.235 -173.975 -58.065 -173.805 ;
        RECT -49.680 -173.975 -49.510 -173.805 ;
        RECT -48.315 -173.975 -48.145 -173.805 ;
        RECT -39.760 -173.975 -39.590 -173.805 ;
        RECT -38.395 -173.975 -38.225 -173.805 ;
        RECT -29.840 -173.975 -29.670 -173.805 ;
        RECT -28.475 -173.975 -28.305 -173.805 ;
        RECT -19.920 -173.975 -19.750 -173.805 ;
        RECT -18.555 -173.975 -18.385 -173.805 ;
        RECT -10.000 -173.975 -9.830 -173.805 ;
        RECT -8.635 -173.975 -8.465 -173.805 ;
        RECT -0.080 -173.975 0.090 -173.805 ;
        RECT 1.285 -173.975 1.455 -173.805 ;
        RECT 9.840 -173.975 10.010 -173.805 ;
        RECT 11.205 -173.975 11.375 -173.805 ;
        RECT 19.760 -173.975 19.930 -173.805 ;
        RECT 21.125 -173.975 21.295 -173.805 ;
        RECT -288.585 -174.405 -288.415 -174.235 ;
        RECT -288.585 -174.865 -288.415 -174.695 ;
        RECT -287.025 -174.825 -286.855 -174.655 ;
        RECT -281.165 -174.825 -280.995 -174.655 ;
        RECT -277.105 -174.825 -276.935 -174.655 ;
        RECT -271.245 -174.825 -271.075 -174.655 ;
        RECT -267.185 -174.825 -267.015 -174.655 ;
        RECT -261.325 -174.825 -261.155 -174.655 ;
        RECT -257.265 -174.825 -257.095 -174.655 ;
        RECT -251.405 -174.825 -251.235 -174.655 ;
        RECT -247.345 -174.825 -247.175 -174.655 ;
        RECT -241.485 -174.825 -241.315 -174.655 ;
        RECT -237.425 -174.825 -237.255 -174.655 ;
        RECT -231.565 -174.825 -231.395 -174.655 ;
        RECT -227.505 -174.825 -227.335 -174.655 ;
        RECT -221.645 -174.825 -221.475 -174.655 ;
        RECT -217.585 -174.825 -217.415 -174.655 ;
        RECT -211.725 -174.825 -211.555 -174.655 ;
        RECT -207.665 -174.825 -207.495 -174.655 ;
        RECT -201.805 -174.825 -201.635 -174.655 ;
        RECT -197.745 -174.825 -197.575 -174.655 ;
        RECT -191.885 -174.825 -191.715 -174.655 ;
        RECT -187.825 -174.825 -187.655 -174.655 ;
        RECT -181.965 -174.825 -181.795 -174.655 ;
        RECT -177.905 -174.825 -177.735 -174.655 ;
        RECT -172.045 -174.825 -171.875 -174.655 ;
        RECT -167.985 -174.825 -167.815 -174.655 ;
        RECT -162.125 -174.825 -161.955 -174.655 ;
        RECT -158.065 -174.825 -157.895 -174.655 ;
        RECT -152.205 -174.825 -152.035 -174.655 ;
        RECT -148.145 -174.825 -147.975 -174.655 ;
        RECT -142.285 -174.825 -142.115 -174.655 ;
        RECT -138.225 -174.825 -138.055 -174.655 ;
        RECT -132.365 -174.825 -132.195 -174.655 ;
        RECT -128.305 -174.825 -128.135 -174.655 ;
        RECT -122.445 -174.825 -122.275 -174.655 ;
        RECT -118.385 -174.825 -118.215 -174.655 ;
        RECT -112.525 -174.825 -112.355 -174.655 ;
        RECT -108.465 -174.825 -108.295 -174.655 ;
        RECT -102.605 -174.825 -102.435 -174.655 ;
        RECT -98.545 -174.825 -98.375 -174.655 ;
        RECT -92.685 -174.825 -92.515 -174.655 ;
        RECT -88.625 -174.825 -88.455 -174.655 ;
        RECT -82.765 -174.825 -82.595 -174.655 ;
        RECT -78.705 -174.825 -78.535 -174.655 ;
        RECT -72.845 -174.825 -72.675 -174.655 ;
        RECT -68.785 -174.825 -68.615 -174.655 ;
        RECT -62.925 -174.825 -62.755 -174.655 ;
        RECT -58.865 -174.825 -58.695 -174.655 ;
        RECT -53.005 -174.825 -52.835 -174.655 ;
        RECT -48.945 -174.825 -48.775 -174.655 ;
        RECT -43.085 -174.825 -42.915 -174.655 ;
        RECT -39.025 -174.825 -38.855 -174.655 ;
        RECT -33.165 -174.825 -32.995 -174.655 ;
        RECT -29.105 -174.825 -28.935 -174.655 ;
        RECT -23.245 -174.825 -23.075 -174.655 ;
        RECT -19.185 -174.825 -19.015 -174.655 ;
        RECT -13.325 -174.825 -13.155 -174.655 ;
        RECT -9.265 -174.825 -9.095 -174.655 ;
        RECT -3.405 -174.825 -3.235 -174.655 ;
        RECT 0.655 -174.825 0.825 -174.655 ;
        RECT 6.515 -174.825 6.685 -174.655 ;
        RECT 10.575 -174.825 10.745 -174.655 ;
        RECT 16.435 -174.825 16.605 -174.655 ;
        RECT 20.495 -174.825 20.665 -174.655 ;
        RECT 26.355 -174.825 26.525 -174.655 ;
        RECT -289.055 -175.525 -288.885 -175.355 ;
        RECT -288.595 -175.525 -288.425 -175.355 ;
        RECT -288.135 -175.525 -287.965 -175.355 ;
        RECT -287.675 -175.525 -287.505 -175.355 ;
        RECT 27.005 -175.525 27.175 -175.355 ;
        RECT 27.465 -175.525 27.635 -175.355 ;
        RECT 27.925 -175.525 28.095 -175.355 ;
        RECT 28.385 -175.525 28.555 -175.355 ;
        RECT -287.705 -176.245 -287.535 -176.075 ;
        RECT -287.720 -176.685 -287.550 -176.515 ;
        RECT -280.485 -176.245 -280.315 -176.075 ;
        RECT -285.430 -177.085 -285.260 -176.915 ;
        RECT -285.445 -177.525 -285.275 -177.355 ;
        RECT -280.470 -176.685 -280.300 -176.515 ;
        RECT -282.760 -177.085 -282.590 -176.915 ;
        RECT -277.785 -176.245 -277.615 -176.075 ;
        RECT -277.800 -176.685 -277.630 -176.515 ;
        RECT -270.565 -176.245 -270.395 -176.075 ;
        RECT -282.745 -177.525 -282.575 -177.355 ;
        RECT -275.510 -177.085 -275.340 -176.915 ;
        RECT -275.525 -177.525 -275.355 -177.355 ;
        RECT -270.550 -176.685 -270.380 -176.515 ;
        RECT -272.840 -177.085 -272.670 -176.915 ;
        RECT -267.865 -176.245 -267.695 -176.075 ;
        RECT -267.880 -176.685 -267.710 -176.515 ;
        RECT -260.645 -176.245 -260.475 -176.075 ;
        RECT -272.825 -177.525 -272.655 -177.355 ;
        RECT -265.590 -177.085 -265.420 -176.915 ;
        RECT -265.605 -177.525 -265.435 -177.355 ;
        RECT -260.630 -176.685 -260.460 -176.515 ;
        RECT -262.920 -177.085 -262.750 -176.915 ;
        RECT -257.945 -176.245 -257.775 -176.075 ;
        RECT -257.960 -176.685 -257.790 -176.515 ;
        RECT -250.725 -176.245 -250.555 -176.075 ;
        RECT -262.905 -177.525 -262.735 -177.355 ;
        RECT -255.670 -177.085 -255.500 -176.915 ;
        RECT -255.685 -177.525 -255.515 -177.355 ;
        RECT -250.710 -176.685 -250.540 -176.515 ;
        RECT -253.000 -177.085 -252.830 -176.915 ;
        RECT -248.025 -176.245 -247.855 -176.075 ;
        RECT -248.040 -176.685 -247.870 -176.515 ;
        RECT -240.805 -176.245 -240.635 -176.075 ;
        RECT -252.985 -177.525 -252.815 -177.355 ;
        RECT -245.750 -177.085 -245.580 -176.915 ;
        RECT -245.765 -177.525 -245.595 -177.355 ;
        RECT -240.790 -176.685 -240.620 -176.515 ;
        RECT -243.080 -177.085 -242.910 -176.915 ;
        RECT -238.105 -176.245 -237.935 -176.075 ;
        RECT -238.120 -176.685 -237.950 -176.515 ;
        RECT -230.885 -176.245 -230.715 -176.075 ;
        RECT -243.065 -177.525 -242.895 -177.355 ;
        RECT -235.830 -177.085 -235.660 -176.915 ;
        RECT -235.845 -177.525 -235.675 -177.355 ;
        RECT -230.870 -176.685 -230.700 -176.515 ;
        RECT -233.160 -177.085 -232.990 -176.915 ;
        RECT -228.185 -176.245 -228.015 -176.075 ;
        RECT -228.200 -176.685 -228.030 -176.515 ;
        RECT -220.965 -176.245 -220.795 -176.075 ;
        RECT -233.145 -177.525 -232.975 -177.355 ;
        RECT -225.910 -177.085 -225.740 -176.915 ;
        RECT -225.925 -177.525 -225.755 -177.355 ;
        RECT -220.950 -176.685 -220.780 -176.515 ;
        RECT -223.240 -177.085 -223.070 -176.915 ;
        RECT -218.265 -176.245 -218.095 -176.075 ;
        RECT -218.280 -176.685 -218.110 -176.515 ;
        RECT -211.045 -176.245 -210.875 -176.075 ;
        RECT -223.225 -177.525 -223.055 -177.355 ;
        RECT -215.990 -177.085 -215.820 -176.915 ;
        RECT -216.005 -177.525 -215.835 -177.355 ;
        RECT -211.030 -176.685 -210.860 -176.515 ;
        RECT -213.320 -177.085 -213.150 -176.915 ;
        RECT -208.345 -176.245 -208.175 -176.075 ;
        RECT -208.360 -176.685 -208.190 -176.515 ;
        RECT -201.125 -176.245 -200.955 -176.075 ;
        RECT -213.305 -177.525 -213.135 -177.355 ;
        RECT -206.070 -177.085 -205.900 -176.915 ;
        RECT -206.085 -177.525 -205.915 -177.355 ;
        RECT -201.110 -176.685 -200.940 -176.515 ;
        RECT -203.400 -177.085 -203.230 -176.915 ;
        RECT -198.425 -176.245 -198.255 -176.075 ;
        RECT -198.440 -176.685 -198.270 -176.515 ;
        RECT -191.205 -176.245 -191.035 -176.075 ;
        RECT -203.385 -177.525 -203.215 -177.355 ;
        RECT -196.150 -177.085 -195.980 -176.915 ;
        RECT -196.165 -177.525 -195.995 -177.355 ;
        RECT -191.190 -176.685 -191.020 -176.515 ;
        RECT -193.480 -177.085 -193.310 -176.915 ;
        RECT -188.505 -176.245 -188.335 -176.075 ;
        RECT -188.520 -176.685 -188.350 -176.515 ;
        RECT -181.285 -176.245 -181.115 -176.075 ;
        RECT -193.465 -177.525 -193.295 -177.355 ;
        RECT -186.230 -177.085 -186.060 -176.915 ;
        RECT -186.245 -177.525 -186.075 -177.355 ;
        RECT -181.270 -176.685 -181.100 -176.515 ;
        RECT -183.560 -177.085 -183.390 -176.915 ;
        RECT -178.585 -176.245 -178.415 -176.075 ;
        RECT -178.600 -176.685 -178.430 -176.515 ;
        RECT -171.365 -176.245 -171.195 -176.075 ;
        RECT -183.545 -177.525 -183.375 -177.355 ;
        RECT -176.310 -177.085 -176.140 -176.915 ;
        RECT -176.325 -177.525 -176.155 -177.355 ;
        RECT -171.350 -176.685 -171.180 -176.515 ;
        RECT -173.640 -177.085 -173.470 -176.915 ;
        RECT -168.665 -176.245 -168.495 -176.075 ;
        RECT -168.680 -176.685 -168.510 -176.515 ;
        RECT -161.445 -176.245 -161.275 -176.075 ;
        RECT -173.625 -177.525 -173.455 -177.355 ;
        RECT -166.390 -177.085 -166.220 -176.915 ;
        RECT -166.405 -177.525 -166.235 -177.355 ;
        RECT -161.430 -176.685 -161.260 -176.515 ;
        RECT -163.720 -177.085 -163.550 -176.915 ;
        RECT -158.745 -176.245 -158.575 -176.075 ;
        RECT -158.760 -176.685 -158.590 -176.515 ;
        RECT -151.525 -176.245 -151.355 -176.075 ;
        RECT -163.705 -177.525 -163.535 -177.355 ;
        RECT -156.470 -177.085 -156.300 -176.915 ;
        RECT -156.485 -177.525 -156.315 -177.355 ;
        RECT -151.510 -176.685 -151.340 -176.515 ;
        RECT -153.800 -177.085 -153.630 -176.915 ;
        RECT -148.825 -176.245 -148.655 -176.075 ;
        RECT -148.840 -176.685 -148.670 -176.515 ;
        RECT -141.605 -176.245 -141.435 -176.075 ;
        RECT -153.785 -177.525 -153.615 -177.355 ;
        RECT -146.550 -177.085 -146.380 -176.915 ;
        RECT -146.565 -177.525 -146.395 -177.355 ;
        RECT -141.590 -176.685 -141.420 -176.515 ;
        RECT -143.880 -177.085 -143.710 -176.915 ;
        RECT -138.905 -176.245 -138.735 -176.075 ;
        RECT -138.920 -176.685 -138.750 -176.515 ;
        RECT -131.685 -176.245 -131.515 -176.075 ;
        RECT -143.865 -177.525 -143.695 -177.355 ;
        RECT -136.630 -177.085 -136.460 -176.915 ;
        RECT -136.645 -177.525 -136.475 -177.355 ;
        RECT -131.670 -176.685 -131.500 -176.515 ;
        RECT -133.960 -177.085 -133.790 -176.915 ;
        RECT -128.985 -176.245 -128.815 -176.075 ;
        RECT -129.000 -176.685 -128.830 -176.515 ;
        RECT -121.765 -176.245 -121.595 -176.075 ;
        RECT -133.945 -177.525 -133.775 -177.355 ;
        RECT -126.710 -177.085 -126.540 -176.915 ;
        RECT -126.725 -177.525 -126.555 -177.355 ;
        RECT -121.750 -176.685 -121.580 -176.515 ;
        RECT -124.040 -177.085 -123.870 -176.915 ;
        RECT -119.065 -176.245 -118.895 -176.075 ;
        RECT -119.080 -176.685 -118.910 -176.515 ;
        RECT -111.845 -176.245 -111.675 -176.075 ;
        RECT -124.025 -177.525 -123.855 -177.355 ;
        RECT -116.790 -177.085 -116.620 -176.915 ;
        RECT -116.805 -177.525 -116.635 -177.355 ;
        RECT -111.830 -176.685 -111.660 -176.515 ;
        RECT -114.120 -177.085 -113.950 -176.915 ;
        RECT -109.145 -176.245 -108.975 -176.075 ;
        RECT -109.160 -176.685 -108.990 -176.515 ;
        RECT -101.925 -176.245 -101.755 -176.075 ;
        RECT -114.105 -177.525 -113.935 -177.355 ;
        RECT -106.870 -177.085 -106.700 -176.915 ;
        RECT -106.885 -177.525 -106.715 -177.355 ;
        RECT -101.910 -176.685 -101.740 -176.515 ;
        RECT -104.200 -177.085 -104.030 -176.915 ;
        RECT -99.225 -176.245 -99.055 -176.075 ;
        RECT -99.240 -176.685 -99.070 -176.515 ;
        RECT -92.005 -176.245 -91.835 -176.075 ;
        RECT -104.185 -177.525 -104.015 -177.355 ;
        RECT -96.950 -177.085 -96.780 -176.915 ;
        RECT -96.965 -177.525 -96.795 -177.355 ;
        RECT -91.990 -176.685 -91.820 -176.515 ;
        RECT -94.280 -177.085 -94.110 -176.915 ;
        RECT -89.305 -176.245 -89.135 -176.075 ;
        RECT -89.320 -176.685 -89.150 -176.515 ;
        RECT -82.085 -176.245 -81.915 -176.075 ;
        RECT -94.265 -177.525 -94.095 -177.355 ;
        RECT -87.030 -177.085 -86.860 -176.915 ;
        RECT -87.045 -177.525 -86.875 -177.355 ;
        RECT -82.070 -176.685 -81.900 -176.515 ;
        RECT -84.360 -177.085 -84.190 -176.915 ;
        RECT -79.385 -176.245 -79.215 -176.075 ;
        RECT -79.400 -176.685 -79.230 -176.515 ;
        RECT -72.165 -176.245 -71.995 -176.075 ;
        RECT -84.345 -177.525 -84.175 -177.355 ;
        RECT -77.110 -177.085 -76.940 -176.915 ;
        RECT -77.125 -177.525 -76.955 -177.355 ;
        RECT -72.150 -176.685 -71.980 -176.515 ;
        RECT -74.440 -177.085 -74.270 -176.915 ;
        RECT -69.465 -176.245 -69.295 -176.075 ;
        RECT -69.480 -176.685 -69.310 -176.515 ;
        RECT -62.245 -176.245 -62.075 -176.075 ;
        RECT -74.425 -177.525 -74.255 -177.355 ;
        RECT -67.190 -177.085 -67.020 -176.915 ;
        RECT -67.205 -177.525 -67.035 -177.355 ;
        RECT -62.230 -176.685 -62.060 -176.515 ;
        RECT -64.520 -177.085 -64.350 -176.915 ;
        RECT -59.545 -176.245 -59.375 -176.075 ;
        RECT -59.560 -176.685 -59.390 -176.515 ;
        RECT -52.325 -176.245 -52.155 -176.075 ;
        RECT -64.505 -177.525 -64.335 -177.355 ;
        RECT -57.270 -177.085 -57.100 -176.915 ;
        RECT -57.285 -177.525 -57.115 -177.355 ;
        RECT -52.310 -176.685 -52.140 -176.515 ;
        RECT -54.600 -177.085 -54.430 -176.915 ;
        RECT -49.625 -176.245 -49.455 -176.075 ;
        RECT -49.640 -176.685 -49.470 -176.515 ;
        RECT -42.405 -176.245 -42.235 -176.075 ;
        RECT -54.585 -177.525 -54.415 -177.355 ;
        RECT -47.350 -177.085 -47.180 -176.915 ;
        RECT -47.365 -177.525 -47.195 -177.355 ;
        RECT -42.390 -176.685 -42.220 -176.515 ;
        RECT -44.680 -177.085 -44.510 -176.915 ;
        RECT -39.705 -176.245 -39.535 -176.075 ;
        RECT -39.720 -176.685 -39.550 -176.515 ;
        RECT -32.485 -176.245 -32.315 -176.075 ;
        RECT -44.665 -177.525 -44.495 -177.355 ;
        RECT -37.430 -177.085 -37.260 -176.915 ;
        RECT -37.445 -177.525 -37.275 -177.355 ;
        RECT -32.470 -176.685 -32.300 -176.515 ;
        RECT -34.760 -177.085 -34.590 -176.915 ;
        RECT -29.785 -176.245 -29.615 -176.075 ;
        RECT -29.800 -176.685 -29.630 -176.515 ;
        RECT -22.565 -176.245 -22.395 -176.075 ;
        RECT -34.745 -177.525 -34.575 -177.355 ;
        RECT -27.510 -177.085 -27.340 -176.915 ;
        RECT -27.525 -177.525 -27.355 -177.355 ;
        RECT -22.550 -176.685 -22.380 -176.515 ;
        RECT -24.840 -177.085 -24.670 -176.915 ;
        RECT -19.865 -176.245 -19.695 -176.075 ;
        RECT -19.880 -176.685 -19.710 -176.515 ;
        RECT -12.645 -176.245 -12.475 -176.075 ;
        RECT -24.825 -177.525 -24.655 -177.355 ;
        RECT -17.590 -177.085 -17.420 -176.915 ;
        RECT -17.605 -177.525 -17.435 -177.355 ;
        RECT -12.630 -176.685 -12.460 -176.515 ;
        RECT -14.920 -177.085 -14.750 -176.915 ;
        RECT -9.945 -176.245 -9.775 -176.075 ;
        RECT -9.960 -176.685 -9.790 -176.515 ;
        RECT -2.725 -176.245 -2.555 -176.075 ;
        RECT -14.905 -177.525 -14.735 -177.355 ;
        RECT -7.670 -177.085 -7.500 -176.915 ;
        RECT -7.685 -177.525 -7.515 -177.355 ;
        RECT -2.710 -176.685 -2.540 -176.515 ;
        RECT -5.000 -177.085 -4.830 -176.915 ;
        RECT -0.025 -176.245 0.145 -176.075 ;
        RECT -0.040 -176.685 0.130 -176.515 ;
        RECT 7.195 -176.245 7.365 -176.075 ;
        RECT -4.985 -177.525 -4.815 -177.355 ;
        RECT 2.250 -177.085 2.420 -176.915 ;
        RECT 2.235 -177.525 2.405 -177.355 ;
        RECT 7.210 -176.685 7.380 -176.515 ;
        RECT 4.920 -177.085 5.090 -176.915 ;
        RECT 9.895 -176.245 10.065 -176.075 ;
        RECT 9.880 -176.685 10.050 -176.515 ;
        RECT 17.115 -176.245 17.285 -176.075 ;
        RECT 4.935 -177.525 5.105 -177.355 ;
        RECT 12.170 -177.085 12.340 -176.915 ;
        RECT 12.155 -177.525 12.325 -177.355 ;
        RECT 17.130 -176.685 17.300 -176.515 ;
        RECT 14.840 -177.085 15.010 -176.915 ;
        RECT 19.815 -176.245 19.985 -176.075 ;
        RECT 19.800 -176.685 19.970 -176.515 ;
        RECT 27.035 -176.245 27.205 -176.075 ;
        RECT 14.855 -177.525 15.025 -177.355 ;
        RECT 22.090 -177.085 22.260 -176.915 ;
        RECT 22.075 -177.525 22.245 -177.355 ;
        RECT 27.050 -176.685 27.220 -176.515 ;
        RECT 24.760 -177.085 24.930 -176.915 ;
        RECT 24.775 -177.525 24.945 -177.355 ;
        RECT -289.055 -178.245 -288.885 -178.075 ;
        RECT -288.595 -178.245 -288.425 -178.075 ;
        RECT -288.135 -178.245 -287.965 -178.075 ;
        RECT -287.675 -178.245 -287.505 -178.075 ;
        RECT -287.285 -178.905 -287.115 -178.735 ;
        RECT -287.285 -179.365 -287.115 -179.195 ;
        RECT -286.125 -178.945 -285.955 -178.775 ;
        RECT -282.065 -178.945 -281.895 -178.775 ;
        RECT -276.205 -178.945 -276.035 -178.775 ;
        RECT -272.145 -178.945 -271.975 -178.775 ;
        RECT -266.285 -178.945 -266.115 -178.775 ;
        RECT -262.225 -178.945 -262.055 -178.775 ;
        RECT -256.365 -178.945 -256.195 -178.775 ;
        RECT -252.305 -178.945 -252.135 -178.775 ;
        RECT -246.445 -178.945 -246.275 -178.775 ;
        RECT -242.385 -178.945 -242.215 -178.775 ;
        RECT -236.525 -178.945 -236.355 -178.775 ;
        RECT -232.465 -178.945 -232.295 -178.775 ;
        RECT -226.605 -178.945 -226.435 -178.775 ;
        RECT -222.545 -178.945 -222.375 -178.775 ;
        RECT -216.685 -178.945 -216.515 -178.775 ;
        RECT -212.625 -178.945 -212.455 -178.775 ;
        RECT -206.765 -178.945 -206.595 -178.775 ;
        RECT -202.705 -178.945 -202.535 -178.775 ;
        RECT -196.845 -178.945 -196.675 -178.775 ;
        RECT -192.785 -178.945 -192.615 -178.775 ;
        RECT -186.925 -178.945 -186.755 -178.775 ;
        RECT -182.865 -178.945 -182.695 -178.775 ;
        RECT -177.005 -178.945 -176.835 -178.775 ;
        RECT -172.945 -178.945 -172.775 -178.775 ;
        RECT -167.085 -178.945 -166.915 -178.775 ;
        RECT -163.025 -178.945 -162.855 -178.775 ;
        RECT -157.165 -178.945 -156.995 -178.775 ;
        RECT -153.105 -178.945 -152.935 -178.775 ;
        RECT -147.245 -178.945 -147.075 -178.775 ;
        RECT -143.185 -178.945 -143.015 -178.775 ;
        RECT -137.325 -178.945 -137.155 -178.775 ;
        RECT -133.265 -178.945 -133.095 -178.775 ;
        RECT -127.405 -178.945 -127.235 -178.775 ;
        RECT -123.345 -178.945 -123.175 -178.775 ;
        RECT -117.485 -178.945 -117.315 -178.775 ;
        RECT -113.425 -178.945 -113.255 -178.775 ;
        RECT -107.565 -178.945 -107.395 -178.775 ;
        RECT -103.505 -178.945 -103.335 -178.775 ;
        RECT -97.645 -178.945 -97.475 -178.775 ;
        RECT -93.585 -178.945 -93.415 -178.775 ;
        RECT -87.725 -178.945 -87.555 -178.775 ;
        RECT -83.665 -178.945 -83.495 -178.775 ;
        RECT -77.805 -178.945 -77.635 -178.775 ;
        RECT -73.745 -178.945 -73.575 -178.775 ;
        RECT -67.885 -178.945 -67.715 -178.775 ;
        RECT -63.825 -178.945 -63.655 -178.775 ;
        RECT -57.965 -178.945 -57.795 -178.775 ;
        RECT -53.905 -178.945 -53.735 -178.775 ;
        RECT -48.045 -178.945 -47.875 -178.775 ;
        RECT -43.985 -178.945 -43.815 -178.775 ;
        RECT -38.125 -178.945 -37.955 -178.775 ;
        RECT -34.065 -178.945 -33.895 -178.775 ;
        RECT -28.205 -178.945 -28.035 -178.775 ;
        RECT -24.145 -178.945 -23.975 -178.775 ;
        RECT -18.285 -178.945 -18.115 -178.775 ;
        RECT -14.225 -178.945 -14.055 -178.775 ;
        RECT -8.365 -178.945 -8.195 -178.775 ;
        RECT -4.305 -178.945 -4.135 -178.775 ;
        RECT 1.555 -178.945 1.725 -178.775 ;
        RECT 5.615 -178.945 5.785 -178.775 ;
        RECT 11.475 -178.945 11.645 -178.775 ;
        RECT 15.535 -178.945 15.705 -178.775 ;
        RECT 21.395 -178.945 21.565 -178.775 ;
        RECT 25.455 -178.945 25.625 -178.775 ;
        RECT 26.615 -178.905 26.785 -178.735 ;
        RECT 26.615 -179.365 26.785 -179.195 ;
        RECT -287.755 -179.815 -287.585 -179.645 ;
        RECT -287.285 -179.825 -287.115 -179.655 ;
        RECT -282.800 -179.795 -282.630 -179.625 ;
        RECT -281.435 -179.795 -281.265 -179.625 ;
        RECT -272.880 -179.795 -272.710 -179.625 ;
        RECT -271.515 -179.795 -271.345 -179.625 ;
        RECT -262.960 -179.795 -262.790 -179.625 ;
        RECT -261.595 -179.795 -261.425 -179.625 ;
        RECT -253.040 -179.795 -252.870 -179.625 ;
        RECT -251.675 -179.795 -251.505 -179.625 ;
        RECT -243.120 -179.795 -242.950 -179.625 ;
        RECT -241.755 -179.795 -241.585 -179.625 ;
        RECT -233.200 -179.795 -233.030 -179.625 ;
        RECT -231.835 -179.795 -231.665 -179.625 ;
        RECT -223.280 -179.795 -223.110 -179.625 ;
        RECT -221.915 -179.795 -221.745 -179.625 ;
        RECT -213.360 -179.795 -213.190 -179.625 ;
        RECT -211.995 -179.795 -211.825 -179.625 ;
        RECT -203.440 -179.795 -203.270 -179.625 ;
        RECT -202.075 -179.795 -201.905 -179.625 ;
        RECT -193.520 -179.795 -193.350 -179.625 ;
        RECT -192.155 -179.795 -191.985 -179.625 ;
        RECT -183.600 -179.795 -183.430 -179.625 ;
        RECT -182.235 -179.795 -182.065 -179.625 ;
        RECT -173.680 -179.795 -173.510 -179.625 ;
        RECT -172.315 -179.795 -172.145 -179.625 ;
        RECT -163.760 -179.795 -163.590 -179.625 ;
        RECT -162.395 -179.795 -162.225 -179.625 ;
        RECT -153.840 -179.795 -153.670 -179.625 ;
        RECT -152.475 -179.795 -152.305 -179.625 ;
        RECT -143.920 -179.795 -143.750 -179.625 ;
        RECT -142.555 -179.795 -142.385 -179.625 ;
        RECT -134.000 -179.795 -133.830 -179.625 ;
        RECT -132.635 -179.795 -132.465 -179.625 ;
        RECT -124.080 -179.795 -123.910 -179.625 ;
        RECT -122.715 -179.795 -122.545 -179.625 ;
        RECT -114.160 -179.795 -113.990 -179.625 ;
        RECT -112.795 -179.795 -112.625 -179.625 ;
        RECT -104.240 -179.795 -104.070 -179.625 ;
        RECT -102.875 -179.795 -102.705 -179.625 ;
        RECT -94.320 -179.795 -94.150 -179.625 ;
        RECT -92.955 -179.795 -92.785 -179.625 ;
        RECT -84.400 -179.795 -84.230 -179.625 ;
        RECT -83.035 -179.795 -82.865 -179.625 ;
        RECT -74.480 -179.795 -74.310 -179.625 ;
        RECT -73.115 -179.795 -72.945 -179.625 ;
        RECT -64.560 -179.795 -64.390 -179.625 ;
        RECT -63.195 -179.795 -63.025 -179.625 ;
        RECT -54.640 -179.795 -54.470 -179.625 ;
        RECT -53.275 -179.795 -53.105 -179.625 ;
        RECT -44.720 -179.795 -44.550 -179.625 ;
        RECT -43.355 -179.795 -43.185 -179.625 ;
        RECT -34.800 -179.795 -34.630 -179.625 ;
        RECT -33.435 -179.795 -33.265 -179.625 ;
        RECT -24.880 -179.795 -24.710 -179.625 ;
        RECT -23.515 -179.795 -23.345 -179.625 ;
        RECT -14.960 -179.795 -14.790 -179.625 ;
        RECT -13.595 -179.795 -13.425 -179.625 ;
        RECT -5.040 -179.795 -4.870 -179.625 ;
        RECT -3.675 -179.795 -3.505 -179.625 ;
        RECT 4.880 -179.795 5.050 -179.625 ;
        RECT 6.245 -179.795 6.415 -179.625 ;
        RECT 14.800 -179.795 14.970 -179.625 ;
        RECT 16.165 -179.795 16.335 -179.625 ;
        RECT 24.720 -179.795 24.890 -179.625 ;
        RECT 26.085 -179.795 26.255 -179.625 ;
        RECT 26.615 -179.825 26.785 -179.655 ;
        RECT 27.085 -179.815 27.255 -179.645 ;
      LAYER met1 ;
        RECT -291.460 95.140 -291.000 95.145 ;
        RECT -291.460 94.665 -290.520 95.140 ;
        RECT -289.600 95.060 -288.600 95.760 ;
        RECT -279.680 95.060 -278.680 95.760 ;
        RECT -269.760 95.060 -268.760 95.760 ;
        RECT -259.840 95.060 -258.840 95.760 ;
        RECT -249.920 95.060 -248.920 95.760 ;
        RECT -240.000 95.060 -239.000 95.760 ;
        RECT -230.080 95.060 -229.080 95.760 ;
        RECT -220.160 95.060 -219.160 95.760 ;
        RECT -210.240 95.060 -209.240 95.760 ;
        RECT -200.320 95.060 -199.320 95.760 ;
        RECT -190.400 95.060 -189.400 95.760 ;
        RECT -180.480 95.060 -179.480 95.760 ;
        RECT -170.560 95.060 -169.560 95.760 ;
        RECT -160.640 95.060 -159.640 95.760 ;
        RECT -150.720 95.060 -149.720 95.760 ;
        RECT -140.800 95.060 -139.800 95.760 ;
        RECT -130.880 95.060 -129.880 95.760 ;
        RECT -120.960 95.060 -119.960 95.760 ;
        RECT -111.040 95.060 -110.040 95.760 ;
        RECT -101.120 95.060 -100.120 95.760 ;
        RECT -91.200 95.060 -90.200 95.760 ;
        RECT -81.280 95.060 -80.280 95.760 ;
        RECT -71.360 95.060 -70.360 95.760 ;
        RECT -61.440 95.060 -60.440 95.760 ;
        RECT -51.520 95.060 -50.520 95.760 ;
        RECT -41.600 95.060 -40.600 95.760 ;
        RECT -31.680 95.060 -30.680 95.760 ;
        RECT -21.760 95.060 -20.760 95.760 ;
        RECT -11.840 95.060 -10.840 95.760 ;
        RECT -1.920 95.060 -0.920 95.760 ;
        RECT 8.000 95.060 9.000 95.760 ;
        RECT 17.920 95.060 18.920 95.760 ;
        RECT -290.110 94.760 -288.420 95.060 ;
        RECT -280.190 94.760 -278.500 95.060 ;
        RECT -270.270 94.760 -268.580 95.060 ;
        RECT -260.350 94.760 -258.660 95.060 ;
        RECT -250.430 94.760 -248.740 95.060 ;
        RECT -240.510 94.760 -238.820 95.060 ;
        RECT -230.590 94.760 -228.900 95.060 ;
        RECT -220.670 94.760 -218.980 95.060 ;
        RECT -210.750 94.760 -209.060 95.060 ;
        RECT -200.830 94.760 -199.140 95.060 ;
        RECT -190.910 94.760 -189.220 95.060 ;
        RECT -180.990 94.760 -179.300 95.060 ;
        RECT -171.070 94.760 -169.380 95.060 ;
        RECT -161.150 94.760 -159.460 95.060 ;
        RECT -151.230 94.760 -149.540 95.060 ;
        RECT -141.310 94.760 -139.620 95.060 ;
        RECT -131.390 94.760 -129.700 95.060 ;
        RECT -121.470 94.760 -119.780 95.060 ;
        RECT -111.550 94.760 -109.860 95.060 ;
        RECT -101.630 94.760 -99.940 95.060 ;
        RECT -91.710 94.760 -90.020 95.060 ;
        RECT -81.790 94.760 -80.100 95.060 ;
        RECT -71.870 94.760 -70.180 95.060 ;
        RECT -61.950 94.760 -60.260 95.060 ;
        RECT -52.030 94.760 -50.340 95.060 ;
        RECT -42.110 94.760 -40.420 95.060 ;
        RECT -32.190 94.760 -30.500 95.060 ;
        RECT -22.270 94.760 -20.580 95.060 ;
        RECT -12.350 94.760 -10.660 95.060 ;
        RECT -2.430 94.760 -0.740 95.060 ;
        RECT 7.490 94.760 9.180 95.060 ;
        RECT 17.410 94.760 19.100 95.060 ;
        RECT -291.000 93.760 -290.520 94.665 ;
        RECT -289.370 93.890 -289.050 94.180 ;
        RECT -283.490 93.890 -283.170 94.180 ;
        RECT -279.450 93.890 -279.130 94.180 ;
        RECT -273.570 93.890 -273.250 94.180 ;
        RECT -269.530 93.890 -269.210 94.180 ;
        RECT -263.650 93.890 -263.330 94.180 ;
        RECT -259.610 93.890 -259.290 94.180 ;
        RECT -253.730 93.890 -253.410 94.180 ;
        RECT -249.690 93.890 -249.370 94.180 ;
        RECT -243.810 93.890 -243.490 94.180 ;
        RECT -239.770 93.890 -239.450 94.180 ;
        RECT -233.890 93.890 -233.570 94.180 ;
        RECT -229.850 93.890 -229.530 94.180 ;
        RECT -223.970 93.890 -223.650 94.180 ;
        RECT -219.930 93.890 -219.610 94.180 ;
        RECT -214.050 93.890 -213.730 94.180 ;
        RECT -210.010 93.890 -209.690 94.180 ;
        RECT -204.130 93.890 -203.810 94.180 ;
        RECT -200.090 93.890 -199.770 94.180 ;
        RECT -194.210 93.890 -193.890 94.180 ;
        RECT -190.170 93.890 -189.850 94.180 ;
        RECT -184.290 93.890 -183.970 94.180 ;
        RECT -180.250 93.890 -179.930 94.180 ;
        RECT -174.370 93.890 -174.050 94.180 ;
        RECT -170.330 93.890 -170.010 94.180 ;
        RECT -164.450 93.890 -164.130 94.180 ;
        RECT -160.410 93.890 -160.090 94.180 ;
        RECT -154.530 93.890 -154.210 94.180 ;
        RECT -150.490 93.890 -150.170 94.180 ;
        RECT -144.610 93.890 -144.290 94.180 ;
        RECT -140.570 93.890 -140.250 94.180 ;
        RECT -134.690 93.890 -134.370 94.180 ;
        RECT -130.650 93.890 -130.330 94.180 ;
        RECT -124.770 93.890 -124.450 94.180 ;
        RECT -120.730 93.890 -120.410 94.180 ;
        RECT -114.850 93.890 -114.530 94.180 ;
        RECT -110.810 93.890 -110.490 94.180 ;
        RECT -104.930 93.890 -104.610 94.180 ;
        RECT -100.890 93.890 -100.570 94.180 ;
        RECT -95.010 93.890 -94.690 94.180 ;
        RECT -90.970 93.890 -90.650 94.180 ;
        RECT -85.090 93.890 -84.770 94.180 ;
        RECT -81.050 93.890 -80.730 94.180 ;
        RECT -75.170 93.890 -74.850 94.180 ;
        RECT -71.130 93.890 -70.810 94.180 ;
        RECT -65.250 93.890 -64.930 94.180 ;
        RECT -61.210 93.890 -60.890 94.180 ;
        RECT -55.330 93.890 -55.010 94.180 ;
        RECT -51.290 93.890 -50.970 94.180 ;
        RECT -45.410 93.890 -45.090 94.180 ;
        RECT -41.370 93.890 -41.050 94.180 ;
        RECT -35.490 93.890 -35.170 94.180 ;
        RECT -31.450 93.890 -31.130 94.180 ;
        RECT -25.570 93.890 -25.250 94.180 ;
        RECT -21.530 93.890 -21.210 94.180 ;
        RECT -15.650 93.890 -15.330 94.180 ;
        RECT -11.610 93.890 -11.290 94.180 ;
        RECT -5.730 93.890 -5.410 94.180 ;
        RECT -1.690 93.890 -1.370 94.180 ;
        RECT 4.190 93.890 4.510 94.180 ;
        RECT 8.230 93.890 8.550 94.180 ;
        RECT 14.110 93.890 14.430 94.180 ;
        RECT 18.150 93.890 18.470 94.180 ;
        RECT 24.030 93.890 24.350 94.180 ;
        RECT -291.460 93.090 -289.620 93.570 ;
        RECT -289.290 92.760 -289.100 93.890 ;
        RECT -283.440 92.760 -283.250 93.890 ;
        RECT -279.370 92.760 -279.180 93.890 ;
        RECT -273.520 92.760 -273.330 93.890 ;
        RECT -269.450 92.760 -269.260 93.890 ;
        RECT -263.600 92.760 -263.410 93.890 ;
        RECT -259.530 92.760 -259.340 93.890 ;
        RECT -253.680 92.760 -253.490 93.890 ;
        RECT -249.610 92.760 -249.420 93.890 ;
        RECT -243.760 92.760 -243.570 93.890 ;
        RECT -239.690 92.760 -239.500 93.890 ;
        RECT -233.840 92.760 -233.650 93.890 ;
        RECT -229.770 92.760 -229.580 93.890 ;
        RECT -223.920 92.760 -223.730 93.890 ;
        RECT -219.850 92.760 -219.660 93.890 ;
        RECT -214.000 92.760 -213.810 93.890 ;
        RECT -209.930 92.760 -209.740 93.890 ;
        RECT -204.080 92.760 -203.890 93.890 ;
        RECT -200.010 92.760 -199.820 93.890 ;
        RECT -194.160 92.760 -193.970 93.890 ;
        RECT -190.090 92.760 -189.900 93.890 ;
        RECT -184.240 92.760 -184.050 93.890 ;
        RECT -180.170 92.760 -179.980 93.890 ;
        RECT -174.320 92.760 -174.130 93.890 ;
        RECT -170.250 92.760 -170.060 93.890 ;
        RECT -164.400 92.760 -164.210 93.890 ;
        RECT -160.330 92.760 -160.140 93.890 ;
        RECT -154.480 92.760 -154.290 93.890 ;
        RECT -150.410 92.760 -150.220 93.890 ;
        RECT -144.560 92.760 -144.370 93.890 ;
        RECT -140.490 92.760 -140.300 93.890 ;
        RECT -134.640 92.760 -134.450 93.890 ;
        RECT -130.570 92.760 -130.380 93.890 ;
        RECT -124.720 92.760 -124.530 93.890 ;
        RECT -120.650 92.760 -120.460 93.890 ;
        RECT -114.800 92.760 -114.610 93.890 ;
        RECT -110.730 92.760 -110.540 93.890 ;
        RECT -104.880 92.760 -104.690 93.890 ;
        RECT -100.810 92.760 -100.620 93.890 ;
        RECT -94.960 92.760 -94.770 93.890 ;
        RECT -90.890 92.760 -90.700 93.890 ;
        RECT -85.040 92.760 -84.850 93.890 ;
        RECT -80.970 92.760 -80.780 93.890 ;
        RECT -75.120 92.760 -74.930 93.890 ;
        RECT -71.050 92.760 -70.860 93.890 ;
        RECT -65.200 92.760 -65.010 93.890 ;
        RECT -61.130 92.760 -60.940 93.890 ;
        RECT -55.280 92.760 -55.090 93.890 ;
        RECT -51.210 92.760 -51.020 93.890 ;
        RECT -45.360 92.760 -45.170 93.890 ;
        RECT -41.290 92.760 -41.100 93.890 ;
        RECT -35.440 92.760 -35.250 93.890 ;
        RECT -31.370 92.760 -31.180 93.890 ;
        RECT -25.520 92.760 -25.330 93.890 ;
        RECT -21.450 92.760 -21.260 93.890 ;
        RECT -15.600 92.760 -15.410 93.890 ;
        RECT -11.530 92.760 -11.340 93.890 ;
        RECT -5.680 92.760 -5.490 93.890 ;
        RECT -1.610 92.760 -1.420 93.890 ;
        RECT 4.240 92.760 4.430 93.890 ;
        RECT 8.310 92.760 8.500 93.890 ;
        RECT 14.160 92.760 14.350 93.890 ;
        RECT 18.230 92.760 18.420 93.890 ;
        RECT 24.080 92.760 24.270 93.890 ;
        RECT 24.600 93.090 26.440 93.570 ;
        RECT -290.050 92.610 -288.110 92.760 ;
        RECT -290.050 92.460 -289.710 92.610 ;
        RECT -290.050 92.260 -289.730 92.290 ;
        RECT -290.050 92.120 -289.230 92.260 ;
        RECT -290.050 92.010 -289.730 92.120 ;
        RECT -289.390 91.330 -289.230 92.120 ;
        RECT -288.270 91.820 -288.110 92.610 ;
        RECT -284.430 92.610 -282.490 92.760 ;
        RECT -287.770 91.820 -287.450 91.930 ;
        RECT -288.270 91.680 -287.450 91.820 ;
        RECT -287.770 91.650 -287.450 91.680 ;
        RECT -285.090 91.820 -284.770 91.930 ;
        RECT -284.430 91.820 -284.270 92.610 ;
        RECT -282.830 92.460 -282.490 92.610 ;
        RECT -280.130 92.610 -278.190 92.760 ;
        RECT -280.130 92.460 -279.790 92.610 ;
        RECT -282.810 92.260 -282.490 92.290 ;
        RECT -285.090 91.680 -284.270 91.820 ;
        RECT -283.310 92.120 -282.490 92.260 ;
        RECT -285.090 91.650 -284.770 91.680 ;
        RECT -287.790 91.330 -287.450 91.480 ;
        RECT -289.390 91.180 -287.450 91.330 ;
        RECT -285.090 91.330 -284.750 91.480 ;
        RECT -283.310 91.330 -283.150 92.120 ;
        RECT -282.810 92.010 -282.490 92.120 ;
        RECT -280.130 92.260 -279.810 92.290 ;
        RECT -280.130 92.120 -279.310 92.260 ;
        RECT -280.130 92.010 -279.810 92.120 ;
        RECT -285.090 91.180 -283.150 91.330 ;
        RECT -279.470 91.330 -279.310 92.120 ;
        RECT -278.350 91.820 -278.190 92.610 ;
        RECT -274.510 92.610 -272.570 92.760 ;
        RECT -277.850 91.820 -277.530 91.930 ;
        RECT -278.350 91.680 -277.530 91.820 ;
        RECT -277.850 91.650 -277.530 91.680 ;
        RECT -275.170 91.820 -274.850 91.930 ;
        RECT -274.510 91.820 -274.350 92.610 ;
        RECT -272.910 92.460 -272.570 92.610 ;
        RECT -270.210 92.610 -268.270 92.760 ;
        RECT -270.210 92.460 -269.870 92.610 ;
        RECT -272.890 92.260 -272.570 92.290 ;
        RECT -275.170 91.680 -274.350 91.820 ;
        RECT -273.390 92.120 -272.570 92.260 ;
        RECT -275.170 91.650 -274.850 91.680 ;
        RECT -277.870 91.330 -277.530 91.480 ;
        RECT -279.470 91.180 -277.530 91.330 ;
        RECT -275.170 91.330 -274.830 91.480 ;
        RECT -273.390 91.330 -273.230 92.120 ;
        RECT -272.890 92.010 -272.570 92.120 ;
        RECT -270.210 92.260 -269.890 92.290 ;
        RECT -270.210 92.120 -269.390 92.260 ;
        RECT -270.210 92.010 -269.890 92.120 ;
        RECT -275.170 91.180 -273.230 91.330 ;
        RECT -269.550 91.330 -269.390 92.120 ;
        RECT -268.430 91.820 -268.270 92.610 ;
        RECT -264.590 92.610 -262.650 92.760 ;
        RECT -267.930 91.820 -267.610 91.930 ;
        RECT -268.430 91.680 -267.610 91.820 ;
        RECT -267.930 91.650 -267.610 91.680 ;
        RECT -265.250 91.820 -264.930 91.930 ;
        RECT -264.590 91.820 -264.430 92.610 ;
        RECT -262.990 92.460 -262.650 92.610 ;
        RECT -260.290 92.610 -258.350 92.760 ;
        RECT -260.290 92.460 -259.950 92.610 ;
        RECT -262.970 92.260 -262.650 92.290 ;
        RECT -265.250 91.680 -264.430 91.820 ;
        RECT -263.470 92.120 -262.650 92.260 ;
        RECT -265.250 91.650 -264.930 91.680 ;
        RECT -267.950 91.330 -267.610 91.480 ;
        RECT -269.550 91.180 -267.610 91.330 ;
        RECT -265.250 91.330 -264.910 91.480 ;
        RECT -263.470 91.330 -263.310 92.120 ;
        RECT -262.970 92.010 -262.650 92.120 ;
        RECT -260.290 92.260 -259.970 92.290 ;
        RECT -260.290 92.120 -259.470 92.260 ;
        RECT -260.290 92.010 -259.970 92.120 ;
        RECT -265.250 91.180 -263.310 91.330 ;
        RECT -259.630 91.330 -259.470 92.120 ;
        RECT -258.510 91.820 -258.350 92.610 ;
        RECT -254.670 92.610 -252.730 92.760 ;
        RECT -258.010 91.820 -257.690 91.930 ;
        RECT -258.510 91.680 -257.690 91.820 ;
        RECT -258.010 91.650 -257.690 91.680 ;
        RECT -255.330 91.820 -255.010 91.930 ;
        RECT -254.670 91.820 -254.510 92.610 ;
        RECT -253.070 92.460 -252.730 92.610 ;
        RECT -250.370 92.610 -248.430 92.760 ;
        RECT -250.370 92.460 -250.030 92.610 ;
        RECT -253.050 92.260 -252.730 92.290 ;
        RECT -255.330 91.680 -254.510 91.820 ;
        RECT -253.550 92.120 -252.730 92.260 ;
        RECT -255.330 91.650 -255.010 91.680 ;
        RECT -258.030 91.330 -257.690 91.480 ;
        RECT -259.630 91.180 -257.690 91.330 ;
        RECT -255.330 91.330 -254.990 91.480 ;
        RECT -253.550 91.330 -253.390 92.120 ;
        RECT -253.050 92.010 -252.730 92.120 ;
        RECT -250.370 92.260 -250.050 92.290 ;
        RECT -250.370 92.120 -249.550 92.260 ;
        RECT -250.370 92.010 -250.050 92.120 ;
        RECT -255.330 91.180 -253.390 91.330 ;
        RECT -249.710 91.330 -249.550 92.120 ;
        RECT -248.590 91.820 -248.430 92.610 ;
        RECT -244.750 92.610 -242.810 92.760 ;
        RECT -248.090 91.820 -247.770 91.930 ;
        RECT -248.590 91.680 -247.770 91.820 ;
        RECT -248.090 91.650 -247.770 91.680 ;
        RECT -245.410 91.820 -245.090 91.930 ;
        RECT -244.750 91.820 -244.590 92.610 ;
        RECT -243.150 92.460 -242.810 92.610 ;
        RECT -240.450 92.610 -238.510 92.760 ;
        RECT -240.450 92.460 -240.110 92.610 ;
        RECT -243.130 92.260 -242.810 92.290 ;
        RECT -245.410 91.680 -244.590 91.820 ;
        RECT -243.630 92.120 -242.810 92.260 ;
        RECT -245.410 91.650 -245.090 91.680 ;
        RECT -248.110 91.330 -247.770 91.480 ;
        RECT -249.710 91.180 -247.770 91.330 ;
        RECT -245.410 91.330 -245.070 91.480 ;
        RECT -243.630 91.330 -243.470 92.120 ;
        RECT -243.130 92.010 -242.810 92.120 ;
        RECT -240.450 92.260 -240.130 92.290 ;
        RECT -240.450 92.120 -239.630 92.260 ;
        RECT -240.450 92.010 -240.130 92.120 ;
        RECT -245.410 91.180 -243.470 91.330 ;
        RECT -239.790 91.330 -239.630 92.120 ;
        RECT -238.670 91.820 -238.510 92.610 ;
        RECT -234.830 92.610 -232.890 92.760 ;
        RECT -238.170 91.820 -237.850 91.930 ;
        RECT -238.670 91.680 -237.850 91.820 ;
        RECT -238.170 91.650 -237.850 91.680 ;
        RECT -235.490 91.820 -235.170 91.930 ;
        RECT -234.830 91.820 -234.670 92.610 ;
        RECT -233.230 92.460 -232.890 92.610 ;
        RECT -230.530 92.610 -228.590 92.760 ;
        RECT -230.530 92.460 -230.190 92.610 ;
        RECT -233.210 92.260 -232.890 92.290 ;
        RECT -235.490 91.680 -234.670 91.820 ;
        RECT -233.710 92.120 -232.890 92.260 ;
        RECT -235.490 91.650 -235.170 91.680 ;
        RECT -238.190 91.330 -237.850 91.480 ;
        RECT -239.790 91.180 -237.850 91.330 ;
        RECT -235.490 91.330 -235.150 91.480 ;
        RECT -233.710 91.330 -233.550 92.120 ;
        RECT -233.210 92.010 -232.890 92.120 ;
        RECT -230.530 92.260 -230.210 92.290 ;
        RECT -230.530 92.120 -229.710 92.260 ;
        RECT -230.530 92.010 -230.210 92.120 ;
        RECT -235.490 91.180 -233.550 91.330 ;
        RECT -229.870 91.330 -229.710 92.120 ;
        RECT -228.750 91.820 -228.590 92.610 ;
        RECT -224.910 92.610 -222.970 92.760 ;
        RECT -228.250 91.820 -227.930 91.930 ;
        RECT -228.750 91.680 -227.930 91.820 ;
        RECT -228.250 91.650 -227.930 91.680 ;
        RECT -225.570 91.820 -225.250 91.930 ;
        RECT -224.910 91.820 -224.750 92.610 ;
        RECT -223.310 92.460 -222.970 92.610 ;
        RECT -220.610 92.610 -218.670 92.760 ;
        RECT -220.610 92.460 -220.270 92.610 ;
        RECT -223.290 92.260 -222.970 92.290 ;
        RECT -225.570 91.680 -224.750 91.820 ;
        RECT -223.790 92.120 -222.970 92.260 ;
        RECT -225.570 91.650 -225.250 91.680 ;
        RECT -228.270 91.330 -227.930 91.480 ;
        RECT -229.870 91.180 -227.930 91.330 ;
        RECT -225.570 91.330 -225.230 91.480 ;
        RECT -223.790 91.330 -223.630 92.120 ;
        RECT -223.290 92.010 -222.970 92.120 ;
        RECT -220.610 92.260 -220.290 92.290 ;
        RECT -220.610 92.120 -219.790 92.260 ;
        RECT -220.610 92.010 -220.290 92.120 ;
        RECT -225.570 91.180 -223.630 91.330 ;
        RECT -219.950 91.330 -219.790 92.120 ;
        RECT -218.830 91.820 -218.670 92.610 ;
        RECT -214.990 92.610 -213.050 92.760 ;
        RECT -218.330 91.820 -218.010 91.930 ;
        RECT -218.830 91.680 -218.010 91.820 ;
        RECT -218.330 91.650 -218.010 91.680 ;
        RECT -215.650 91.820 -215.330 91.930 ;
        RECT -214.990 91.820 -214.830 92.610 ;
        RECT -213.390 92.460 -213.050 92.610 ;
        RECT -210.690 92.610 -208.750 92.760 ;
        RECT -210.690 92.460 -210.350 92.610 ;
        RECT -213.370 92.260 -213.050 92.290 ;
        RECT -215.650 91.680 -214.830 91.820 ;
        RECT -213.870 92.120 -213.050 92.260 ;
        RECT -215.650 91.650 -215.330 91.680 ;
        RECT -218.350 91.330 -218.010 91.480 ;
        RECT -219.950 91.180 -218.010 91.330 ;
        RECT -215.650 91.330 -215.310 91.480 ;
        RECT -213.870 91.330 -213.710 92.120 ;
        RECT -213.370 92.010 -213.050 92.120 ;
        RECT -210.690 92.260 -210.370 92.290 ;
        RECT -210.690 92.120 -209.870 92.260 ;
        RECT -210.690 92.010 -210.370 92.120 ;
        RECT -215.650 91.180 -213.710 91.330 ;
        RECT -210.030 91.330 -209.870 92.120 ;
        RECT -208.910 91.820 -208.750 92.610 ;
        RECT -205.070 92.610 -203.130 92.760 ;
        RECT -208.410 91.820 -208.090 91.930 ;
        RECT -208.910 91.680 -208.090 91.820 ;
        RECT -208.410 91.650 -208.090 91.680 ;
        RECT -205.730 91.820 -205.410 91.930 ;
        RECT -205.070 91.820 -204.910 92.610 ;
        RECT -203.470 92.460 -203.130 92.610 ;
        RECT -200.770 92.610 -198.830 92.760 ;
        RECT -200.770 92.460 -200.430 92.610 ;
        RECT -203.450 92.260 -203.130 92.290 ;
        RECT -205.730 91.680 -204.910 91.820 ;
        RECT -203.950 92.120 -203.130 92.260 ;
        RECT -205.730 91.650 -205.410 91.680 ;
        RECT -208.430 91.330 -208.090 91.480 ;
        RECT -210.030 91.180 -208.090 91.330 ;
        RECT -205.730 91.330 -205.390 91.480 ;
        RECT -203.950 91.330 -203.790 92.120 ;
        RECT -203.450 92.010 -203.130 92.120 ;
        RECT -200.770 92.260 -200.450 92.290 ;
        RECT -200.770 92.120 -199.950 92.260 ;
        RECT -200.770 92.010 -200.450 92.120 ;
        RECT -205.730 91.180 -203.790 91.330 ;
        RECT -200.110 91.330 -199.950 92.120 ;
        RECT -198.990 91.820 -198.830 92.610 ;
        RECT -195.150 92.610 -193.210 92.760 ;
        RECT -198.490 91.820 -198.170 91.930 ;
        RECT -198.990 91.680 -198.170 91.820 ;
        RECT -198.490 91.650 -198.170 91.680 ;
        RECT -195.810 91.820 -195.490 91.930 ;
        RECT -195.150 91.820 -194.990 92.610 ;
        RECT -193.550 92.460 -193.210 92.610 ;
        RECT -190.850 92.610 -188.910 92.760 ;
        RECT -190.850 92.460 -190.510 92.610 ;
        RECT -193.530 92.260 -193.210 92.290 ;
        RECT -195.810 91.680 -194.990 91.820 ;
        RECT -194.030 92.120 -193.210 92.260 ;
        RECT -195.810 91.650 -195.490 91.680 ;
        RECT -198.510 91.330 -198.170 91.480 ;
        RECT -200.110 91.180 -198.170 91.330 ;
        RECT -195.810 91.330 -195.470 91.480 ;
        RECT -194.030 91.330 -193.870 92.120 ;
        RECT -193.530 92.010 -193.210 92.120 ;
        RECT -190.850 92.260 -190.530 92.290 ;
        RECT -190.850 92.120 -190.030 92.260 ;
        RECT -190.850 92.010 -190.530 92.120 ;
        RECT -195.810 91.180 -193.870 91.330 ;
        RECT -190.190 91.330 -190.030 92.120 ;
        RECT -189.070 91.820 -188.910 92.610 ;
        RECT -185.230 92.610 -183.290 92.760 ;
        RECT -188.570 91.820 -188.250 91.930 ;
        RECT -189.070 91.680 -188.250 91.820 ;
        RECT -188.570 91.650 -188.250 91.680 ;
        RECT -185.890 91.820 -185.570 91.930 ;
        RECT -185.230 91.820 -185.070 92.610 ;
        RECT -183.630 92.460 -183.290 92.610 ;
        RECT -180.930 92.610 -178.990 92.760 ;
        RECT -180.930 92.460 -180.590 92.610 ;
        RECT -183.610 92.260 -183.290 92.290 ;
        RECT -185.890 91.680 -185.070 91.820 ;
        RECT -184.110 92.120 -183.290 92.260 ;
        RECT -185.890 91.650 -185.570 91.680 ;
        RECT -188.590 91.330 -188.250 91.480 ;
        RECT -190.190 91.180 -188.250 91.330 ;
        RECT -185.890 91.330 -185.550 91.480 ;
        RECT -184.110 91.330 -183.950 92.120 ;
        RECT -183.610 92.010 -183.290 92.120 ;
        RECT -180.930 92.260 -180.610 92.290 ;
        RECT -180.930 92.120 -180.110 92.260 ;
        RECT -180.930 92.010 -180.610 92.120 ;
        RECT -185.890 91.180 -183.950 91.330 ;
        RECT -180.270 91.330 -180.110 92.120 ;
        RECT -179.150 91.820 -178.990 92.610 ;
        RECT -175.310 92.610 -173.370 92.760 ;
        RECT -178.650 91.820 -178.330 91.930 ;
        RECT -179.150 91.680 -178.330 91.820 ;
        RECT -178.650 91.650 -178.330 91.680 ;
        RECT -175.970 91.820 -175.650 91.930 ;
        RECT -175.310 91.820 -175.150 92.610 ;
        RECT -173.710 92.460 -173.370 92.610 ;
        RECT -171.010 92.610 -169.070 92.760 ;
        RECT -171.010 92.460 -170.670 92.610 ;
        RECT -173.690 92.260 -173.370 92.290 ;
        RECT -175.970 91.680 -175.150 91.820 ;
        RECT -174.190 92.120 -173.370 92.260 ;
        RECT -175.970 91.650 -175.650 91.680 ;
        RECT -178.670 91.330 -178.330 91.480 ;
        RECT -180.270 91.180 -178.330 91.330 ;
        RECT -175.970 91.330 -175.630 91.480 ;
        RECT -174.190 91.330 -174.030 92.120 ;
        RECT -173.690 92.010 -173.370 92.120 ;
        RECT -171.010 92.260 -170.690 92.290 ;
        RECT -171.010 92.120 -170.190 92.260 ;
        RECT -171.010 92.010 -170.690 92.120 ;
        RECT -175.970 91.180 -174.030 91.330 ;
        RECT -170.350 91.330 -170.190 92.120 ;
        RECT -169.230 91.820 -169.070 92.610 ;
        RECT -165.390 92.610 -163.450 92.760 ;
        RECT -168.730 91.820 -168.410 91.930 ;
        RECT -169.230 91.680 -168.410 91.820 ;
        RECT -168.730 91.650 -168.410 91.680 ;
        RECT -166.050 91.820 -165.730 91.930 ;
        RECT -165.390 91.820 -165.230 92.610 ;
        RECT -163.790 92.460 -163.450 92.610 ;
        RECT -161.090 92.610 -159.150 92.760 ;
        RECT -161.090 92.460 -160.750 92.610 ;
        RECT -163.770 92.260 -163.450 92.290 ;
        RECT -166.050 91.680 -165.230 91.820 ;
        RECT -164.270 92.120 -163.450 92.260 ;
        RECT -166.050 91.650 -165.730 91.680 ;
        RECT -168.750 91.330 -168.410 91.480 ;
        RECT -170.350 91.180 -168.410 91.330 ;
        RECT -166.050 91.330 -165.710 91.480 ;
        RECT -164.270 91.330 -164.110 92.120 ;
        RECT -163.770 92.010 -163.450 92.120 ;
        RECT -161.090 92.260 -160.770 92.290 ;
        RECT -161.090 92.120 -160.270 92.260 ;
        RECT -161.090 92.010 -160.770 92.120 ;
        RECT -166.050 91.180 -164.110 91.330 ;
        RECT -160.430 91.330 -160.270 92.120 ;
        RECT -159.310 91.820 -159.150 92.610 ;
        RECT -155.470 92.610 -153.530 92.760 ;
        RECT -158.810 91.820 -158.490 91.930 ;
        RECT -159.310 91.680 -158.490 91.820 ;
        RECT -158.810 91.650 -158.490 91.680 ;
        RECT -156.130 91.820 -155.810 91.930 ;
        RECT -155.470 91.820 -155.310 92.610 ;
        RECT -153.870 92.460 -153.530 92.610 ;
        RECT -151.170 92.610 -149.230 92.760 ;
        RECT -151.170 92.460 -150.830 92.610 ;
        RECT -153.850 92.260 -153.530 92.290 ;
        RECT -156.130 91.680 -155.310 91.820 ;
        RECT -154.350 92.120 -153.530 92.260 ;
        RECT -156.130 91.650 -155.810 91.680 ;
        RECT -158.830 91.330 -158.490 91.480 ;
        RECT -160.430 91.180 -158.490 91.330 ;
        RECT -156.130 91.330 -155.790 91.480 ;
        RECT -154.350 91.330 -154.190 92.120 ;
        RECT -153.850 92.010 -153.530 92.120 ;
        RECT -151.170 92.260 -150.850 92.290 ;
        RECT -151.170 92.120 -150.350 92.260 ;
        RECT -151.170 92.010 -150.850 92.120 ;
        RECT -156.130 91.180 -154.190 91.330 ;
        RECT -150.510 91.330 -150.350 92.120 ;
        RECT -149.390 91.820 -149.230 92.610 ;
        RECT -145.550 92.610 -143.610 92.760 ;
        RECT -148.890 91.820 -148.570 91.930 ;
        RECT -149.390 91.680 -148.570 91.820 ;
        RECT -148.890 91.650 -148.570 91.680 ;
        RECT -146.210 91.820 -145.890 91.930 ;
        RECT -145.550 91.820 -145.390 92.610 ;
        RECT -143.950 92.460 -143.610 92.610 ;
        RECT -141.250 92.610 -139.310 92.760 ;
        RECT -141.250 92.460 -140.910 92.610 ;
        RECT -143.930 92.260 -143.610 92.290 ;
        RECT -146.210 91.680 -145.390 91.820 ;
        RECT -144.430 92.120 -143.610 92.260 ;
        RECT -146.210 91.650 -145.890 91.680 ;
        RECT -148.910 91.330 -148.570 91.480 ;
        RECT -150.510 91.180 -148.570 91.330 ;
        RECT -146.210 91.330 -145.870 91.480 ;
        RECT -144.430 91.330 -144.270 92.120 ;
        RECT -143.930 92.010 -143.610 92.120 ;
        RECT -141.250 92.260 -140.930 92.290 ;
        RECT -141.250 92.120 -140.430 92.260 ;
        RECT -141.250 92.010 -140.930 92.120 ;
        RECT -146.210 91.180 -144.270 91.330 ;
        RECT -140.590 91.330 -140.430 92.120 ;
        RECT -139.470 91.820 -139.310 92.610 ;
        RECT -135.630 92.610 -133.690 92.760 ;
        RECT -138.970 91.820 -138.650 91.930 ;
        RECT -139.470 91.680 -138.650 91.820 ;
        RECT -138.970 91.650 -138.650 91.680 ;
        RECT -136.290 91.820 -135.970 91.930 ;
        RECT -135.630 91.820 -135.470 92.610 ;
        RECT -134.030 92.460 -133.690 92.610 ;
        RECT -131.330 92.610 -129.390 92.760 ;
        RECT -131.330 92.460 -130.990 92.610 ;
        RECT -134.010 92.260 -133.690 92.290 ;
        RECT -136.290 91.680 -135.470 91.820 ;
        RECT -134.510 92.120 -133.690 92.260 ;
        RECT -136.290 91.650 -135.970 91.680 ;
        RECT -138.990 91.330 -138.650 91.480 ;
        RECT -140.590 91.180 -138.650 91.330 ;
        RECT -136.290 91.330 -135.950 91.480 ;
        RECT -134.510 91.330 -134.350 92.120 ;
        RECT -134.010 92.010 -133.690 92.120 ;
        RECT -131.330 92.260 -131.010 92.290 ;
        RECT -131.330 92.120 -130.510 92.260 ;
        RECT -131.330 92.010 -131.010 92.120 ;
        RECT -136.290 91.180 -134.350 91.330 ;
        RECT -130.670 91.330 -130.510 92.120 ;
        RECT -129.550 91.820 -129.390 92.610 ;
        RECT -125.710 92.610 -123.770 92.760 ;
        RECT -129.050 91.820 -128.730 91.930 ;
        RECT -129.550 91.680 -128.730 91.820 ;
        RECT -129.050 91.650 -128.730 91.680 ;
        RECT -126.370 91.820 -126.050 91.930 ;
        RECT -125.710 91.820 -125.550 92.610 ;
        RECT -124.110 92.460 -123.770 92.610 ;
        RECT -121.410 92.610 -119.470 92.760 ;
        RECT -121.410 92.460 -121.070 92.610 ;
        RECT -124.090 92.260 -123.770 92.290 ;
        RECT -126.370 91.680 -125.550 91.820 ;
        RECT -124.590 92.120 -123.770 92.260 ;
        RECT -126.370 91.650 -126.050 91.680 ;
        RECT -129.070 91.330 -128.730 91.480 ;
        RECT -130.670 91.180 -128.730 91.330 ;
        RECT -126.370 91.330 -126.030 91.480 ;
        RECT -124.590 91.330 -124.430 92.120 ;
        RECT -124.090 92.010 -123.770 92.120 ;
        RECT -121.410 92.260 -121.090 92.290 ;
        RECT -121.410 92.120 -120.590 92.260 ;
        RECT -121.410 92.010 -121.090 92.120 ;
        RECT -126.370 91.180 -124.430 91.330 ;
        RECT -120.750 91.330 -120.590 92.120 ;
        RECT -119.630 91.820 -119.470 92.610 ;
        RECT -115.790 92.610 -113.850 92.760 ;
        RECT -119.130 91.820 -118.810 91.930 ;
        RECT -119.630 91.680 -118.810 91.820 ;
        RECT -119.130 91.650 -118.810 91.680 ;
        RECT -116.450 91.820 -116.130 91.930 ;
        RECT -115.790 91.820 -115.630 92.610 ;
        RECT -114.190 92.460 -113.850 92.610 ;
        RECT -111.490 92.610 -109.550 92.760 ;
        RECT -111.490 92.460 -111.150 92.610 ;
        RECT -114.170 92.260 -113.850 92.290 ;
        RECT -116.450 91.680 -115.630 91.820 ;
        RECT -114.670 92.120 -113.850 92.260 ;
        RECT -116.450 91.650 -116.130 91.680 ;
        RECT -119.150 91.330 -118.810 91.480 ;
        RECT -120.750 91.180 -118.810 91.330 ;
        RECT -116.450 91.330 -116.110 91.480 ;
        RECT -114.670 91.330 -114.510 92.120 ;
        RECT -114.170 92.010 -113.850 92.120 ;
        RECT -111.490 92.260 -111.170 92.290 ;
        RECT -111.490 92.120 -110.670 92.260 ;
        RECT -111.490 92.010 -111.170 92.120 ;
        RECT -116.450 91.180 -114.510 91.330 ;
        RECT -110.830 91.330 -110.670 92.120 ;
        RECT -109.710 91.820 -109.550 92.610 ;
        RECT -105.870 92.610 -103.930 92.760 ;
        RECT -109.210 91.820 -108.890 91.930 ;
        RECT -109.710 91.680 -108.890 91.820 ;
        RECT -109.210 91.650 -108.890 91.680 ;
        RECT -106.530 91.820 -106.210 91.930 ;
        RECT -105.870 91.820 -105.710 92.610 ;
        RECT -104.270 92.460 -103.930 92.610 ;
        RECT -101.570 92.610 -99.630 92.760 ;
        RECT -101.570 92.460 -101.230 92.610 ;
        RECT -104.250 92.260 -103.930 92.290 ;
        RECT -106.530 91.680 -105.710 91.820 ;
        RECT -104.750 92.120 -103.930 92.260 ;
        RECT -106.530 91.650 -106.210 91.680 ;
        RECT -109.230 91.330 -108.890 91.480 ;
        RECT -110.830 91.180 -108.890 91.330 ;
        RECT -106.530 91.330 -106.190 91.480 ;
        RECT -104.750 91.330 -104.590 92.120 ;
        RECT -104.250 92.010 -103.930 92.120 ;
        RECT -101.570 92.260 -101.250 92.290 ;
        RECT -101.570 92.120 -100.750 92.260 ;
        RECT -101.570 92.010 -101.250 92.120 ;
        RECT -106.530 91.180 -104.590 91.330 ;
        RECT -100.910 91.330 -100.750 92.120 ;
        RECT -99.790 91.820 -99.630 92.610 ;
        RECT -95.950 92.610 -94.010 92.760 ;
        RECT -99.290 91.820 -98.970 91.930 ;
        RECT -99.790 91.680 -98.970 91.820 ;
        RECT -99.290 91.650 -98.970 91.680 ;
        RECT -96.610 91.820 -96.290 91.930 ;
        RECT -95.950 91.820 -95.790 92.610 ;
        RECT -94.350 92.460 -94.010 92.610 ;
        RECT -91.650 92.610 -89.710 92.760 ;
        RECT -91.650 92.460 -91.310 92.610 ;
        RECT -94.330 92.260 -94.010 92.290 ;
        RECT -96.610 91.680 -95.790 91.820 ;
        RECT -94.830 92.120 -94.010 92.260 ;
        RECT -96.610 91.650 -96.290 91.680 ;
        RECT -99.310 91.330 -98.970 91.480 ;
        RECT -100.910 91.180 -98.970 91.330 ;
        RECT -96.610 91.330 -96.270 91.480 ;
        RECT -94.830 91.330 -94.670 92.120 ;
        RECT -94.330 92.010 -94.010 92.120 ;
        RECT -91.650 92.260 -91.330 92.290 ;
        RECT -91.650 92.120 -90.830 92.260 ;
        RECT -91.650 92.010 -91.330 92.120 ;
        RECT -96.610 91.180 -94.670 91.330 ;
        RECT -90.990 91.330 -90.830 92.120 ;
        RECT -89.870 91.820 -89.710 92.610 ;
        RECT -86.030 92.610 -84.090 92.760 ;
        RECT -89.370 91.820 -89.050 91.930 ;
        RECT -89.870 91.680 -89.050 91.820 ;
        RECT -89.370 91.650 -89.050 91.680 ;
        RECT -86.690 91.820 -86.370 91.930 ;
        RECT -86.030 91.820 -85.870 92.610 ;
        RECT -84.430 92.460 -84.090 92.610 ;
        RECT -81.730 92.610 -79.790 92.760 ;
        RECT -81.730 92.460 -81.390 92.610 ;
        RECT -84.410 92.260 -84.090 92.290 ;
        RECT -86.690 91.680 -85.870 91.820 ;
        RECT -84.910 92.120 -84.090 92.260 ;
        RECT -86.690 91.650 -86.370 91.680 ;
        RECT -89.390 91.330 -89.050 91.480 ;
        RECT -90.990 91.180 -89.050 91.330 ;
        RECT -86.690 91.330 -86.350 91.480 ;
        RECT -84.910 91.330 -84.750 92.120 ;
        RECT -84.410 92.010 -84.090 92.120 ;
        RECT -81.730 92.260 -81.410 92.290 ;
        RECT -81.730 92.120 -80.910 92.260 ;
        RECT -81.730 92.010 -81.410 92.120 ;
        RECT -86.690 91.180 -84.750 91.330 ;
        RECT -81.070 91.330 -80.910 92.120 ;
        RECT -79.950 91.820 -79.790 92.610 ;
        RECT -76.110 92.610 -74.170 92.760 ;
        RECT -79.450 91.820 -79.130 91.930 ;
        RECT -79.950 91.680 -79.130 91.820 ;
        RECT -79.450 91.650 -79.130 91.680 ;
        RECT -76.770 91.820 -76.450 91.930 ;
        RECT -76.110 91.820 -75.950 92.610 ;
        RECT -74.510 92.460 -74.170 92.610 ;
        RECT -71.810 92.610 -69.870 92.760 ;
        RECT -71.810 92.460 -71.470 92.610 ;
        RECT -74.490 92.260 -74.170 92.290 ;
        RECT -76.770 91.680 -75.950 91.820 ;
        RECT -74.990 92.120 -74.170 92.260 ;
        RECT -76.770 91.650 -76.450 91.680 ;
        RECT -79.470 91.330 -79.130 91.480 ;
        RECT -81.070 91.180 -79.130 91.330 ;
        RECT -76.770 91.330 -76.430 91.480 ;
        RECT -74.990 91.330 -74.830 92.120 ;
        RECT -74.490 92.010 -74.170 92.120 ;
        RECT -71.810 92.260 -71.490 92.290 ;
        RECT -71.810 92.120 -70.990 92.260 ;
        RECT -71.810 92.010 -71.490 92.120 ;
        RECT -76.770 91.180 -74.830 91.330 ;
        RECT -71.150 91.330 -70.990 92.120 ;
        RECT -70.030 91.820 -69.870 92.610 ;
        RECT -66.190 92.610 -64.250 92.760 ;
        RECT -69.530 91.820 -69.210 91.930 ;
        RECT -70.030 91.680 -69.210 91.820 ;
        RECT -69.530 91.650 -69.210 91.680 ;
        RECT -66.850 91.820 -66.530 91.930 ;
        RECT -66.190 91.820 -66.030 92.610 ;
        RECT -64.590 92.460 -64.250 92.610 ;
        RECT -61.890 92.610 -59.950 92.760 ;
        RECT -61.890 92.460 -61.550 92.610 ;
        RECT -64.570 92.260 -64.250 92.290 ;
        RECT -66.850 91.680 -66.030 91.820 ;
        RECT -65.070 92.120 -64.250 92.260 ;
        RECT -66.850 91.650 -66.530 91.680 ;
        RECT -69.550 91.330 -69.210 91.480 ;
        RECT -71.150 91.180 -69.210 91.330 ;
        RECT -66.850 91.330 -66.510 91.480 ;
        RECT -65.070 91.330 -64.910 92.120 ;
        RECT -64.570 92.010 -64.250 92.120 ;
        RECT -61.890 92.260 -61.570 92.290 ;
        RECT -61.890 92.120 -61.070 92.260 ;
        RECT -61.890 92.010 -61.570 92.120 ;
        RECT -66.850 91.180 -64.910 91.330 ;
        RECT -61.230 91.330 -61.070 92.120 ;
        RECT -60.110 91.820 -59.950 92.610 ;
        RECT -56.270 92.610 -54.330 92.760 ;
        RECT -59.610 91.820 -59.290 91.930 ;
        RECT -60.110 91.680 -59.290 91.820 ;
        RECT -59.610 91.650 -59.290 91.680 ;
        RECT -56.930 91.820 -56.610 91.930 ;
        RECT -56.270 91.820 -56.110 92.610 ;
        RECT -54.670 92.460 -54.330 92.610 ;
        RECT -51.970 92.610 -50.030 92.760 ;
        RECT -51.970 92.460 -51.630 92.610 ;
        RECT -54.650 92.260 -54.330 92.290 ;
        RECT -56.930 91.680 -56.110 91.820 ;
        RECT -55.150 92.120 -54.330 92.260 ;
        RECT -56.930 91.650 -56.610 91.680 ;
        RECT -59.630 91.330 -59.290 91.480 ;
        RECT -61.230 91.180 -59.290 91.330 ;
        RECT -56.930 91.330 -56.590 91.480 ;
        RECT -55.150 91.330 -54.990 92.120 ;
        RECT -54.650 92.010 -54.330 92.120 ;
        RECT -51.970 92.260 -51.650 92.290 ;
        RECT -51.970 92.120 -51.150 92.260 ;
        RECT -51.970 92.010 -51.650 92.120 ;
        RECT -56.930 91.180 -54.990 91.330 ;
        RECT -51.310 91.330 -51.150 92.120 ;
        RECT -50.190 91.820 -50.030 92.610 ;
        RECT -46.350 92.610 -44.410 92.760 ;
        RECT -49.690 91.820 -49.370 91.930 ;
        RECT -50.190 91.680 -49.370 91.820 ;
        RECT -49.690 91.650 -49.370 91.680 ;
        RECT -47.010 91.820 -46.690 91.930 ;
        RECT -46.350 91.820 -46.190 92.610 ;
        RECT -44.750 92.460 -44.410 92.610 ;
        RECT -42.050 92.610 -40.110 92.760 ;
        RECT -42.050 92.460 -41.710 92.610 ;
        RECT -44.730 92.260 -44.410 92.290 ;
        RECT -47.010 91.680 -46.190 91.820 ;
        RECT -45.230 92.120 -44.410 92.260 ;
        RECT -47.010 91.650 -46.690 91.680 ;
        RECT -49.710 91.330 -49.370 91.480 ;
        RECT -51.310 91.180 -49.370 91.330 ;
        RECT -47.010 91.330 -46.670 91.480 ;
        RECT -45.230 91.330 -45.070 92.120 ;
        RECT -44.730 92.010 -44.410 92.120 ;
        RECT -42.050 92.260 -41.730 92.290 ;
        RECT -42.050 92.120 -41.230 92.260 ;
        RECT -42.050 92.010 -41.730 92.120 ;
        RECT -47.010 91.180 -45.070 91.330 ;
        RECT -41.390 91.330 -41.230 92.120 ;
        RECT -40.270 91.820 -40.110 92.610 ;
        RECT -36.430 92.610 -34.490 92.760 ;
        RECT -39.770 91.820 -39.450 91.930 ;
        RECT -40.270 91.680 -39.450 91.820 ;
        RECT -39.770 91.650 -39.450 91.680 ;
        RECT -37.090 91.820 -36.770 91.930 ;
        RECT -36.430 91.820 -36.270 92.610 ;
        RECT -34.830 92.460 -34.490 92.610 ;
        RECT -32.130 92.610 -30.190 92.760 ;
        RECT -32.130 92.460 -31.790 92.610 ;
        RECT -34.810 92.260 -34.490 92.290 ;
        RECT -37.090 91.680 -36.270 91.820 ;
        RECT -35.310 92.120 -34.490 92.260 ;
        RECT -37.090 91.650 -36.770 91.680 ;
        RECT -39.790 91.330 -39.450 91.480 ;
        RECT -41.390 91.180 -39.450 91.330 ;
        RECT -37.090 91.330 -36.750 91.480 ;
        RECT -35.310 91.330 -35.150 92.120 ;
        RECT -34.810 92.010 -34.490 92.120 ;
        RECT -32.130 92.260 -31.810 92.290 ;
        RECT -32.130 92.120 -31.310 92.260 ;
        RECT -32.130 92.010 -31.810 92.120 ;
        RECT -37.090 91.180 -35.150 91.330 ;
        RECT -31.470 91.330 -31.310 92.120 ;
        RECT -30.350 91.820 -30.190 92.610 ;
        RECT -26.510 92.610 -24.570 92.760 ;
        RECT -29.850 91.820 -29.530 91.930 ;
        RECT -30.350 91.680 -29.530 91.820 ;
        RECT -29.850 91.650 -29.530 91.680 ;
        RECT -27.170 91.820 -26.850 91.930 ;
        RECT -26.510 91.820 -26.350 92.610 ;
        RECT -24.910 92.460 -24.570 92.610 ;
        RECT -22.210 92.610 -20.270 92.760 ;
        RECT -22.210 92.460 -21.870 92.610 ;
        RECT -24.890 92.260 -24.570 92.290 ;
        RECT -27.170 91.680 -26.350 91.820 ;
        RECT -25.390 92.120 -24.570 92.260 ;
        RECT -27.170 91.650 -26.850 91.680 ;
        RECT -29.870 91.330 -29.530 91.480 ;
        RECT -31.470 91.180 -29.530 91.330 ;
        RECT -27.170 91.330 -26.830 91.480 ;
        RECT -25.390 91.330 -25.230 92.120 ;
        RECT -24.890 92.010 -24.570 92.120 ;
        RECT -22.210 92.260 -21.890 92.290 ;
        RECT -22.210 92.120 -21.390 92.260 ;
        RECT -22.210 92.010 -21.890 92.120 ;
        RECT -27.170 91.180 -25.230 91.330 ;
        RECT -21.550 91.330 -21.390 92.120 ;
        RECT -20.430 91.820 -20.270 92.610 ;
        RECT -16.590 92.610 -14.650 92.760 ;
        RECT -19.930 91.820 -19.610 91.930 ;
        RECT -20.430 91.680 -19.610 91.820 ;
        RECT -19.930 91.650 -19.610 91.680 ;
        RECT -17.250 91.820 -16.930 91.930 ;
        RECT -16.590 91.820 -16.430 92.610 ;
        RECT -14.990 92.460 -14.650 92.610 ;
        RECT -12.290 92.610 -10.350 92.760 ;
        RECT -12.290 92.460 -11.950 92.610 ;
        RECT -14.970 92.260 -14.650 92.290 ;
        RECT -17.250 91.680 -16.430 91.820 ;
        RECT -15.470 92.120 -14.650 92.260 ;
        RECT -17.250 91.650 -16.930 91.680 ;
        RECT -19.950 91.330 -19.610 91.480 ;
        RECT -21.550 91.180 -19.610 91.330 ;
        RECT -17.250 91.330 -16.910 91.480 ;
        RECT -15.470 91.330 -15.310 92.120 ;
        RECT -14.970 92.010 -14.650 92.120 ;
        RECT -12.290 92.260 -11.970 92.290 ;
        RECT -12.290 92.120 -11.470 92.260 ;
        RECT -12.290 92.010 -11.970 92.120 ;
        RECT -17.250 91.180 -15.310 91.330 ;
        RECT -11.630 91.330 -11.470 92.120 ;
        RECT -10.510 91.820 -10.350 92.610 ;
        RECT -6.670 92.610 -4.730 92.760 ;
        RECT -10.010 91.820 -9.690 91.930 ;
        RECT -10.510 91.680 -9.690 91.820 ;
        RECT -10.010 91.650 -9.690 91.680 ;
        RECT -7.330 91.820 -7.010 91.930 ;
        RECT -6.670 91.820 -6.510 92.610 ;
        RECT -5.070 92.460 -4.730 92.610 ;
        RECT -2.370 92.610 -0.430 92.760 ;
        RECT -2.370 92.460 -2.030 92.610 ;
        RECT -5.050 92.260 -4.730 92.290 ;
        RECT -7.330 91.680 -6.510 91.820 ;
        RECT -5.550 92.120 -4.730 92.260 ;
        RECT -7.330 91.650 -7.010 91.680 ;
        RECT -10.030 91.330 -9.690 91.480 ;
        RECT -11.630 91.180 -9.690 91.330 ;
        RECT -7.330 91.330 -6.990 91.480 ;
        RECT -5.550 91.330 -5.390 92.120 ;
        RECT -5.050 92.010 -4.730 92.120 ;
        RECT -2.370 92.260 -2.050 92.290 ;
        RECT -2.370 92.120 -1.550 92.260 ;
        RECT -2.370 92.010 -2.050 92.120 ;
        RECT -7.330 91.180 -5.390 91.330 ;
        RECT -1.710 91.330 -1.550 92.120 ;
        RECT -0.590 91.820 -0.430 92.610 ;
        RECT 3.250 92.610 5.190 92.760 ;
        RECT -0.090 91.820 0.230 91.930 ;
        RECT -0.590 91.680 0.230 91.820 ;
        RECT -0.090 91.650 0.230 91.680 ;
        RECT 2.590 91.820 2.910 91.930 ;
        RECT 3.250 91.820 3.410 92.610 ;
        RECT 4.850 92.460 5.190 92.610 ;
        RECT 7.550 92.610 9.490 92.760 ;
        RECT 7.550 92.460 7.890 92.610 ;
        RECT 4.870 92.260 5.190 92.290 ;
        RECT 2.590 91.680 3.410 91.820 ;
        RECT 4.370 92.120 5.190 92.260 ;
        RECT 2.590 91.650 2.910 91.680 ;
        RECT -0.110 91.330 0.230 91.480 ;
        RECT -1.710 91.180 0.230 91.330 ;
        RECT 2.590 91.330 2.930 91.480 ;
        RECT 4.370 91.330 4.530 92.120 ;
        RECT 4.870 92.010 5.190 92.120 ;
        RECT 7.550 92.260 7.870 92.290 ;
        RECT 7.550 92.120 8.370 92.260 ;
        RECT 7.550 92.010 7.870 92.120 ;
        RECT 2.590 91.180 4.530 91.330 ;
        RECT 8.210 91.330 8.370 92.120 ;
        RECT 9.330 91.820 9.490 92.610 ;
        RECT 13.170 92.610 15.110 92.760 ;
        RECT 9.830 91.820 10.150 91.930 ;
        RECT 9.330 91.680 10.150 91.820 ;
        RECT 9.830 91.650 10.150 91.680 ;
        RECT 12.510 91.820 12.830 91.930 ;
        RECT 13.170 91.820 13.330 92.610 ;
        RECT 14.770 92.460 15.110 92.610 ;
        RECT 17.470 92.610 19.410 92.760 ;
        RECT 17.470 92.460 17.810 92.610 ;
        RECT 14.790 92.260 15.110 92.290 ;
        RECT 12.510 91.680 13.330 91.820 ;
        RECT 14.290 92.120 15.110 92.260 ;
        RECT 12.510 91.650 12.830 91.680 ;
        RECT 9.810 91.330 10.150 91.480 ;
        RECT 8.210 91.180 10.150 91.330 ;
        RECT 12.510 91.330 12.850 91.480 ;
        RECT 14.290 91.330 14.450 92.120 ;
        RECT 14.790 92.010 15.110 92.120 ;
        RECT 17.470 92.260 17.790 92.290 ;
        RECT 17.470 92.120 18.290 92.260 ;
        RECT 17.470 92.010 17.790 92.120 ;
        RECT 12.510 91.180 14.450 91.330 ;
        RECT 18.130 91.330 18.290 92.120 ;
        RECT 19.250 91.820 19.410 92.610 ;
        RECT 23.090 92.610 25.030 92.760 ;
        RECT 19.750 91.820 20.070 91.930 ;
        RECT 19.250 91.680 20.070 91.820 ;
        RECT 19.750 91.650 20.070 91.680 ;
        RECT 22.430 91.820 22.750 91.930 ;
        RECT 23.090 91.820 23.250 92.610 ;
        RECT 24.690 92.460 25.030 92.610 ;
        RECT 24.710 92.260 25.030 92.290 ;
        RECT 22.430 91.680 23.250 91.820 ;
        RECT 24.210 92.120 25.030 92.260 ;
        RECT 22.430 91.650 22.750 91.680 ;
        RECT 19.730 91.330 20.070 91.480 ;
        RECT 18.130 91.180 20.070 91.330 ;
        RECT 22.430 91.330 22.770 91.480 ;
        RECT 24.210 91.330 24.370 92.120 ;
        RECT 24.710 92.010 25.030 92.120 ;
        RECT 22.430 91.180 24.370 91.330 ;
        RECT -291.460 90.370 -289.620 90.850 ;
        RECT -289.700 89.280 -289.220 90.180 ;
        RECT -288.400 90.050 -288.210 91.180 ;
        RECT -284.330 90.050 -284.140 91.180 ;
        RECT -278.480 90.050 -278.290 91.180 ;
        RECT -274.410 90.050 -274.220 91.180 ;
        RECT -268.560 90.050 -268.370 91.180 ;
        RECT -264.490 90.050 -264.300 91.180 ;
        RECT -258.640 90.050 -258.450 91.180 ;
        RECT -254.570 90.050 -254.380 91.180 ;
        RECT -248.720 90.050 -248.530 91.180 ;
        RECT -244.650 90.050 -244.460 91.180 ;
        RECT -238.800 90.050 -238.610 91.180 ;
        RECT -234.730 90.050 -234.540 91.180 ;
        RECT -228.880 90.050 -228.690 91.180 ;
        RECT -224.810 90.050 -224.620 91.180 ;
        RECT -218.960 90.050 -218.770 91.180 ;
        RECT -214.890 90.050 -214.700 91.180 ;
        RECT -209.040 90.050 -208.850 91.180 ;
        RECT -204.970 90.050 -204.780 91.180 ;
        RECT -199.120 90.050 -198.930 91.180 ;
        RECT -195.050 90.050 -194.860 91.180 ;
        RECT -189.200 90.050 -189.010 91.180 ;
        RECT -185.130 90.050 -184.940 91.180 ;
        RECT -179.280 90.050 -179.090 91.180 ;
        RECT -175.210 90.050 -175.020 91.180 ;
        RECT -169.360 90.050 -169.170 91.180 ;
        RECT -165.290 90.050 -165.100 91.180 ;
        RECT -159.440 90.050 -159.250 91.180 ;
        RECT -155.370 90.050 -155.180 91.180 ;
        RECT -149.520 90.050 -149.330 91.180 ;
        RECT -145.450 90.050 -145.260 91.180 ;
        RECT -139.600 90.050 -139.410 91.180 ;
        RECT -135.530 90.050 -135.340 91.180 ;
        RECT -129.680 90.050 -129.490 91.180 ;
        RECT -125.610 90.050 -125.420 91.180 ;
        RECT -119.760 90.050 -119.570 91.180 ;
        RECT -115.690 90.050 -115.500 91.180 ;
        RECT -109.840 90.050 -109.650 91.180 ;
        RECT -105.770 90.050 -105.580 91.180 ;
        RECT -99.920 90.050 -99.730 91.180 ;
        RECT -95.850 90.050 -95.660 91.180 ;
        RECT -90.000 90.050 -89.810 91.180 ;
        RECT -85.930 90.050 -85.740 91.180 ;
        RECT -80.080 90.050 -79.890 91.180 ;
        RECT -76.010 90.050 -75.820 91.180 ;
        RECT -70.160 90.050 -69.970 91.180 ;
        RECT -66.090 90.050 -65.900 91.180 ;
        RECT -60.240 90.050 -60.050 91.180 ;
        RECT -56.170 90.050 -55.980 91.180 ;
        RECT -50.320 90.050 -50.130 91.180 ;
        RECT -46.250 90.050 -46.060 91.180 ;
        RECT -40.400 90.050 -40.210 91.180 ;
        RECT -36.330 90.050 -36.140 91.180 ;
        RECT -30.480 90.050 -30.290 91.180 ;
        RECT -26.410 90.050 -26.220 91.180 ;
        RECT -20.560 90.050 -20.370 91.180 ;
        RECT -16.490 90.050 -16.300 91.180 ;
        RECT -10.640 90.050 -10.450 91.180 ;
        RECT -6.570 90.050 -6.380 91.180 ;
        RECT -0.720 90.050 -0.530 91.180 ;
        RECT 3.350 90.050 3.540 91.180 ;
        RECT 9.200 90.050 9.390 91.180 ;
        RECT 13.270 90.050 13.460 91.180 ;
        RECT 19.120 90.050 19.310 91.180 ;
        RECT 23.190 90.050 23.380 91.180 ;
        RECT -288.450 89.760 -288.130 90.050 ;
        RECT -284.410 89.760 -284.090 90.050 ;
        RECT -278.530 89.760 -278.210 90.050 ;
        RECT -274.490 89.760 -274.170 90.050 ;
        RECT -268.610 89.760 -268.290 90.050 ;
        RECT -264.570 89.760 -264.250 90.050 ;
        RECT -258.690 89.760 -258.370 90.050 ;
        RECT -254.650 89.760 -254.330 90.050 ;
        RECT -248.770 89.760 -248.450 90.050 ;
        RECT -244.730 89.760 -244.410 90.050 ;
        RECT -238.850 89.760 -238.530 90.050 ;
        RECT -234.810 89.760 -234.490 90.050 ;
        RECT -228.930 89.760 -228.610 90.050 ;
        RECT -224.890 89.760 -224.570 90.050 ;
        RECT -219.010 89.760 -218.690 90.050 ;
        RECT -214.970 89.760 -214.650 90.050 ;
        RECT -209.090 89.760 -208.770 90.050 ;
        RECT -205.050 89.760 -204.730 90.050 ;
        RECT -199.170 89.760 -198.850 90.050 ;
        RECT -195.130 89.760 -194.810 90.050 ;
        RECT -189.250 89.760 -188.930 90.050 ;
        RECT -185.210 89.760 -184.890 90.050 ;
        RECT -179.330 89.760 -179.010 90.050 ;
        RECT -175.290 89.760 -174.970 90.050 ;
        RECT -169.410 89.760 -169.090 90.050 ;
        RECT -165.370 89.760 -165.050 90.050 ;
        RECT -159.490 89.760 -159.170 90.050 ;
        RECT -155.450 89.760 -155.130 90.050 ;
        RECT -149.570 89.760 -149.250 90.050 ;
        RECT -145.530 89.760 -145.210 90.050 ;
        RECT -139.650 89.760 -139.330 90.050 ;
        RECT -135.610 89.760 -135.290 90.050 ;
        RECT -129.730 89.760 -129.410 90.050 ;
        RECT -125.690 89.760 -125.370 90.050 ;
        RECT -119.810 89.760 -119.490 90.050 ;
        RECT -115.770 89.760 -115.450 90.050 ;
        RECT -109.890 89.760 -109.570 90.050 ;
        RECT -105.850 89.760 -105.530 90.050 ;
        RECT -99.970 89.760 -99.650 90.050 ;
        RECT -95.930 89.760 -95.610 90.050 ;
        RECT -90.050 89.760 -89.730 90.050 ;
        RECT -86.010 89.760 -85.690 90.050 ;
        RECT -80.130 89.760 -79.810 90.050 ;
        RECT -76.090 89.760 -75.770 90.050 ;
        RECT -70.210 89.760 -69.890 90.050 ;
        RECT -66.170 89.760 -65.850 90.050 ;
        RECT -60.290 89.760 -59.970 90.050 ;
        RECT -56.250 89.760 -55.930 90.050 ;
        RECT -50.370 89.760 -50.050 90.050 ;
        RECT -46.330 89.760 -46.010 90.050 ;
        RECT -40.450 89.760 -40.130 90.050 ;
        RECT -36.410 89.760 -36.090 90.050 ;
        RECT -30.530 89.760 -30.210 90.050 ;
        RECT -26.490 89.760 -26.170 90.050 ;
        RECT -20.610 89.760 -20.290 90.050 ;
        RECT -16.570 89.760 -16.250 90.050 ;
        RECT -10.690 89.760 -10.370 90.050 ;
        RECT -6.650 89.760 -6.330 90.050 ;
        RECT -0.770 89.760 -0.450 90.050 ;
        RECT 3.270 89.760 3.590 90.050 ;
        RECT 9.150 89.760 9.470 90.050 ;
        RECT 13.190 89.760 13.510 90.050 ;
        RECT 19.070 89.760 19.390 90.050 ;
        RECT 23.110 89.760 23.430 90.050 ;
        RECT -290.160 88.800 -289.220 89.280 ;
        RECT 24.200 89.280 24.680 90.180 ;
        RECT -285.150 88.880 -283.460 89.180 ;
        RECT -275.230 88.880 -273.540 89.180 ;
        RECT -265.310 88.880 -263.620 89.180 ;
        RECT -255.390 88.880 -253.700 89.180 ;
        RECT -245.470 88.880 -243.780 89.180 ;
        RECT -235.550 88.880 -233.860 89.180 ;
        RECT -225.630 88.880 -223.940 89.180 ;
        RECT -215.710 88.880 -214.020 89.180 ;
        RECT -205.790 88.880 -204.100 89.180 ;
        RECT -195.870 88.880 -194.180 89.180 ;
        RECT -185.950 88.880 -184.260 89.180 ;
        RECT -176.030 88.880 -174.340 89.180 ;
        RECT -166.110 88.880 -164.420 89.180 ;
        RECT -156.190 88.880 -154.500 89.180 ;
        RECT -146.270 88.880 -144.580 89.180 ;
        RECT -136.350 88.880 -134.660 89.180 ;
        RECT -126.430 88.880 -124.740 89.180 ;
        RECT -116.510 88.880 -114.820 89.180 ;
        RECT -106.590 88.880 -104.900 89.180 ;
        RECT -96.670 88.880 -94.980 89.180 ;
        RECT -86.750 88.880 -85.060 89.180 ;
        RECT -76.830 88.880 -75.140 89.180 ;
        RECT -66.910 88.880 -65.220 89.180 ;
        RECT -56.990 88.880 -55.300 89.180 ;
        RECT -47.070 88.880 -45.380 89.180 ;
        RECT -37.150 88.880 -35.460 89.180 ;
        RECT -27.230 88.880 -25.540 89.180 ;
        RECT -17.310 88.880 -15.620 89.180 ;
        RECT -7.390 88.880 -5.700 89.180 ;
        RECT 2.530 88.880 4.220 89.180 ;
        RECT 12.450 88.880 14.140 89.180 ;
        RECT 22.370 88.880 24.060 89.180 ;
        RECT -284.640 88.180 -283.640 88.880 ;
        RECT -274.720 88.180 -273.720 88.880 ;
        RECT -264.800 88.180 -263.800 88.880 ;
        RECT -254.880 88.180 -253.880 88.880 ;
        RECT -244.960 88.180 -243.960 88.880 ;
        RECT -235.040 88.180 -234.040 88.880 ;
        RECT -225.120 88.180 -224.120 88.880 ;
        RECT -215.200 88.180 -214.200 88.880 ;
        RECT -205.280 88.180 -204.280 88.880 ;
        RECT -195.360 88.180 -194.360 88.880 ;
        RECT -185.440 88.180 -184.440 88.880 ;
        RECT -175.520 88.180 -174.520 88.880 ;
        RECT -165.600 88.180 -164.600 88.880 ;
        RECT -155.680 88.180 -154.680 88.880 ;
        RECT -145.760 88.180 -144.760 88.880 ;
        RECT -135.840 88.180 -134.840 88.880 ;
        RECT -125.920 88.180 -124.920 88.880 ;
        RECT -116.000 88.180 -115.000 88.880 ;
        RECT -106.080 88.180 -105.080 88.880 ;
        RECT -96.160 88.180 -95.160 88.880 ;
        RECT -86.240 88.180 -85.240 88.880 ;
        RECT -76.320 88.180 -75.320 88.880 ;
        RECT -66.400 88.180 -65.400 88.880 ;
        RECT -56.480 88.180 -55.480 88.880 ;
        RECT -46.560 88.180 -45.560 88.880 ;
        RECT -36.640 88.180 -35.640 88.880 ;
        RECT -26.720 88.180 -25.720 88.880 ;
        RECT -16.800 88.180 -15.800 88.880 ;
        RECT -6.880 88.180 -5.880 88.880 ;
        RECT 3.040 88.180 4.040 88.880 ;
        RECT 12.960 88.180 13.960 88.880 ;
        RECT 22.880 88.180 23.880 88.880 ;
        RECT 24.200 88.800 25.140 89.280 ;
        RECT -291.210 7.430 -290.750 7.435 ;
        RECT -291.210 6.955 -290.270 7.430 ;
        RECT -289.350 7.350 -288.350 8.050 ;
        RECT -279.430 7.350 -278.430 8.050 ;
        RECT -269.510 7.350 -268.510 8.050 ;
        RECT -259.590 7.350 -258.590 8.050 ;
        RECT -249.670 7.350 -248.670 8.050 ;
        RECT -239.750 7.350 -238.750 8.050 ;
        RECT -229.830 7.350 -228.830 8.050 ;
        RECT -219.910 7.350 -218.910 8.050 ;
        RECT -209.990 7.350 -208.990 8.050 ;
        RECT -200.070 7.350 -199.070 8.050 ;
        RECT -190.150 7.350 -189.150 8.050 ;
        RECT -180.230 7.350 -179.230 8.050 ;
        RECT -170.310 7.350 -169.310 8.050 ;
        RECT -160.390 7.350 -159.390 8.050 ;
        RECT -150.470 7.350 -149.470 8.050 ;
        RECT -140.550 7.350 -139.550 8.050 ;
        RECT -130.630 7.350 -129.630 8.050 ;
        RECT -120.710 7.350 -119.710 8.050 ;
        RECT -110.790 7.350 -109.790 8.050 ;
        RECT -100.870 7.350 -99.870 8.050 ;
        RECT -90.950 7.350 -89.950 8.050 ;
        RECT -81.030 7.350 -80.030 8.050 ;
        RECT -71.110 7.350 -70.110 8.050 ;
        RECT -61.190 7.350 -60.190 8.050 ;
        RECT -51.270 7.350 -50.270 8.050 ;
        RECT -41.350 7.350 -40.350 8.050 ;
        RECT -31.430 7.350 -30.430 8.050 ;
        RECT -21.510 7.350 -20.510 8.050 ;
        RECT -11.590 7.350 -10.590 8.050 ;
        RECT -1.670 7.350 -0.670 8.050 ;
        RECT 8.250 7.350 9.250 8.050 ;
        RECT 18.170 7.350 19.170 8.050 ;
        RECT -289.860 7.050 -288.170 7.350 ;
        RECT -279.940 7.050 -278.250 7.350 ;
        RECT -270.020 7.050 -268.330 7.350 ;
        RECT -260.100 7.050 -258.410 7.350 ;
        RECT -250.180 7.050 -248.490 7.350 ;
        RECT -240.260 7.050 -238.570 7.350 ;
        RECT -230.340 7.050 -228.650 7.350 ;
        RECT -220.420 7.050 -218.730 7.350 ;
        RECT -210.500 7.050 -208.810 7.350 ;
        RECT -200.580 7.050 -198.890 7.350 ;
        RECT -190.660 7.050 -188.970 7.350 ;
        RECT -180.740 7.050 -179.050 7.350 ;
        RECT -170.820 7.050 -169.130 7.350 ;
        RECT -160.900 7.050 -159.210 7.350 ;
        RECT -150.980 7.050 -149.290 7.350 ;
        RECT -141.060 7.050 -139.370 7.350 ;
        RECT -131.140 7.050 -129.450 7.350 ;
        RECT -121.220 7.050 -119.530 7.350 ;
        RECT -111.300 7.050 -109.610 7.350 ;
        RECT -101.380 7.050 -99.690 7.350 ;
        RECT -91.460 7.050 -89.770 7.350 ;
        RECT -81.540 7.050 -79.850 7.350 ;
        RECT -71.620 7.050 -69.930 7.350 ;
        RECT -61.700 7.050 -60.010 7.350 ;
        RECT -51.780 7.050 -50.090 7.350 ;
        RECT -41.860 7.050 -40.170 7.350 ;
        RECT -31.940 7.050 -30.250 7.350 ;
        RECT -22.020 7.050 -20.330 7.350 ;
        RECT -12.100 7.050 -10.410 7.350 ;
        RECT -2.180 7.050 -0.490 7.350 ;
        RECT 7.740 7.050 9.430 7.350 ;
        RECT 17.660 7.050 19.350 7.350 ;
        RECT -290.750 6.050 -290.270 6.955 ;
        RECT -289.120 6.180 -288.800 6.470 ;
        RECT -283.240 6.180 -282.920 6.470 ;
        RECT -279.200 6.180 -278.880 6.470 ;
        RECT -273.320 6.180 -273.000 6.470 ;
        RECT -269.280 6.180 -268.960 6.470 ;
        RECT -263.400 6.180 -263.080 6.470 ;
        RECT -259.360 6.180 -259.040 6.470 ;
        RECT -253.480 6.180 -253.160 6.470 ;
        RECT -249.440 6.180 -249.120 6.470 ;
        RECT -243.560 6.180 -243.240 6.470 ;
        RECT -239.520 6.180 -239.200 6.470 ;
        RECT -233.640 6.180 -233.320 6.470 ;
        RECT -229.600 6.180 -229.280 6.470 ;
        RECT -223.720 6.180 -223.400 6.470 ;
        RECT -219.680 6.180 -219.360 6.470 ;
        RECT -213.800 6.180 -213.480 6.470 ;
        RECT -209.760 6.180 -209.440 6.470 ;
        RECT -203.880 6.180 -203.560 6.470 ;
        RECT -199.840 6.180 -199.520 6.470 ;
        RECT -193.960 6.180 -193.640 6.470 ;
        RECT -189.920 6.180 -189.600 6.470 ;
        RECT -184.040 6.180 -183.720 6.470 ;
        RECT -180.000 6.180 -179.680 6.470 ;
        RECT -174.120 6.180 -173.800 6.470 ;
        RECT -170.080 6.180 -169.760 6.470 ;
        RECT -164.200 6.180 -163.880 6.470 ;
        RECT -160.160 6.180 -159.840 6.470 ;
        RECT -154.280 6.180 -153.960 6.470 ;
        RECT -150.240 6.180 -149.920 6.470 ;
        RECT -144.360 6.180 -144.040 6.470 ;
        RECT -140.320 6.180 -140.000 6.470 ;
        RECT -134.440 6.180 -134.120 6.470 ;
        RECT -130.400 6.180 -130.080 6.470 ;
        RECT -124.520 6.180 -124.200 6.470 ;
        RECT -120.480 6.180 -120.160 6.470 ;
        RECT -114.600 6.180 -114.280 6.470 ;
        RECT -110.560 6.180 -110.240 6.470 ;
        RECT -104.680 6.180 -104.360 6.470 ;
        RECT -100.640 6.180 -100.320 6.470 ;
        RECT -94.760 6.180 -94.440 6.470 ;
        RECT -90.720 6.180 -90.400 6.470 ;
        RECT -84.840 6.180 -84.520 6.470 ;
        RECT -80.800 6.180 -80.480 6.470 ;
        RECT -74.920 6.180 -74.600 6.470 ;
        RECT -70.880 6.180 -70.560 6.470 ;
        RECT -65.000 6.180 -64.680 6.470 ;
        RECT -60.960 6.180 -60.640 6.470 ;
        RECT -55.080 6.180 -54.760 6.470 ;
        RECT -51.040 6.180 -50.720 6.470 ;
        RECT -45.160 6.180 -44.840 6.470 ;
        RECT -41.120 6.180 -40.800 6.470 ;
        RECT -35.240 6.180 -34.920 6.470 ;
        RECT -31.200 6.180 -30.880 6.470 ;
        RECT -25.320 6.180 -25.000 6.470 ;
        RECT -21.280 6.180 -20.960 6.470 ;
        RECT -15.400 6.180 -15.080 6.470 ;
        RECT -11.360 6.180 -11.040 6.470 ;
        RECT -5.480 6.180 -5.160 6.470 ;
        RECT -1.440 6.180 -1.120 6.470 ;
        RECT 4.440 6.180 4.760 6.470 ;
        RECT 8.480 6.180 8.800 6.470 ;
        RECT 14.360 6.180 14.680 6.470 ;
        RECT 18.400 6.180 18.720 6.470 ;
        RECT 24.280 6.180 24.600 6.470 ;
        RECT -291.210 5.380 -289.370 5.860 ;
        RECT -289.040 5.050 -288.850 6.180 ;
        RECT -283.190 5.050 -283.000 6.180 ;
        RECT -279.120 5.050 -278.930 6.180 ;
        RECT -273.270 5.050 -273.080 6.180 ;
        RECT -269.200 5.050 -269.010 6.180 ;
        RECT -263.350 5.050 -263.160 6.180 ;
        RECT -259.280 5.050 -259.090 6.180 ;
        RECT -253.430 5.050 -253.240 6.180 ;
        RECT -249.360 5.050 -249.170 6.180 ;
        RECT -243.510 5.050 -243.320 6.180 ;
        RECT -239.440 5.050 -239.250 6.180 ;
        RECT -233.590 5.050 -233.400 6.180 ;
        RECT -229.520 5.050 -229.330 6.180 ;
        RECT -223.670 5.050 -223.480 6.180 ;
        RECT -219.600 5.050 -219.410 6.180 ;
        RECT -213.750 5.050 -213.560 6.180 ;
        RECT -209.680 5.050 -209.490 6.180 ;
        RECT -203.830 5.050 -203.640 6.180 ;
        RECT -199.760 5.050 -199.570 6.180 ;
        RECT -193.910 5.050 -193.720 6.180 ;
        RECT -189.840 5.050 -189.650 6.180 ;
        RECT -183.990 5.050 -183.800 6.180 ;
        RECT -179.920 5.050 -179.730 6.180 ;
        RECT -174.070 5.050 -173.880 6.180 ;
        RECT -170.000 5.050 -169.810 6.180 ;
        RECT -164.150 5.050 -163.960 6.180 ;
        RECT -160.080 5.050 -159.890 6.180 ;
        RECT -154.230 5.050 -154.040 6.180 ;
        RECT -150.160 5.050 -149.970 6.180 ;
        RECT -144.310 5.050 -144.120 6.180 ;
        RECT -140.240 5.050 -140.050 6.180 ;
        RECT -134.390 5.050 -134.200 6.180 ;
        RECT -130.320 5.050 -130.130 6.180 ;
        RECT -124.470 5.050 -124.280 6.180 ;
        RECT -120.400 5.050 -120.210 6.180 ;
        RECT -114.550 5.050 -114.360 6.180 ;
        RECT -110.480 5.050 -110.290 6.180 ;
        RECT -104.630 5.050 -104.440 6.180 ;
        RECT -100.560 5.050 -100.370 6.180 ;
        RECT -94.710 5.050 -94.520 6.180 ;
        RECT -90.640 5.050 -90.450 6.180 ;
        RECT -84.790 5.050 -84.600 6.180 ;
        RECT -80.720 5.050 -80.530 6.180 ;
        RECT -74.870 5.050 -74.680 6.180 ;
        RECT -70.800 5.050 -70.610 6.180 ;
        RECT -64.950 5.050 -64.760 6.180 ;
        RECT -60.880 5.050 -60.690 6.180 ;
        RECT -55.030 5.050 -54.840 6.180 ;
        RECT -50.960 5.050 -50.770 6.180 ;
        RECT -45.110 5.050 -44.920 6.180 ;
        RECT -41.040 5.050 -40.850 6.180 ;
        RECT -35.190 5.050 -35.000 6.180 ;
        RECT -31.120 5.050 -30.930 6.180 ;
        RECT -25.270 5.050 -25.080 6.180 ;
        RECT -21.200 5.050 -21.010 6.180 ;
        RECT -15.350 5.050 -15.160 6.180 ;
        RECT -11.280 5.050 -11.090 6.180 ;
        RECT -5.430 5.050 -5.240 6.180 ;
        RECT -1.360 5.050 -1.170 6.180 ;
        RECT 4.490 5.050 4.680 6.180 ;
        RECT 8.560 5.050 8.750 6.180 ;
        RECT 14.410 5.050 14.600 6.180 ;
        RECT 18.480 5.050 18.670 6.180 ;
        RECT 24.330 5.050 24.520 6.180 ;
        RECT 24.850 5.380 26.690 5.860 ;
        RECT -289.800 4.900 -287.860 5.050 ;
        RECT -289.800 4.750 -289.460 4.900 ;
        RECT -289.800 4.550 -289.480 4.580 ;
        RECT -289.800 4.410 -288.980 4.550 ;
        RECT -289.800 4.300 -289.480 4.410 ;
        RECT -289.140 3.620 -288.980 4.410 ;
        RECT -288.020 4.110 -287.860 4.900 ;
        RECT -284.180 4.900 -282.240 5.050 ;
        RECT -287.520 4.110 -287.200 4.220 ;
        RECT -288.020 3.970 -287.200 4.110 ;
        RECT -287.520 3.940 -287.200 3.970 ;
        RECT -284.840 4.110 -284.520 4.220 ;
        RECT -284.180 4.110 -284.020 4.900 ;
        RECT -282.580 4.750 -282.240 4.900 ;
        RECT -279.880 4.900 -277.940 5.050 ;
        RECT -279.880 4.750 -279.540 4.900 ;
        RECT -282.560 4.550 -282.240 4.580 ;
        RECT -284.840 3.970 -284.020 4.110 ;
        RECT -283.060 4.410 -282.240 4.550 ;
        RECT -284.840 3.940 -284.520 3.970 ;
        RECT -287.540 3.620 -287.200 3.770 ;
        RECT -289.140 3.470 -287.200 3.620 ;
        RECT -284.840 3.620 -284.500 3.770 ;
        RECT -283.060 3.620 -282.900 4.410 ;
        RECT -282.560 4.300 -282.240 4.410 ;
        RECT -279.880 4.550 -279.560 4.580 ;
        RECT -279.880 4.410 -279.060 4.550 ;
        RECT -279.880 4.300 -279.560 4.410 ;
        RECT -284.840 3.470 -282.900 3.620 ;
        RECT -279.220 3.620 -279.060 4.410 ;
        RECT -278.100 4.110 -277.940 4.900 ;
        RECT -274.260 4.900 -272.320 5.050 ;
        RECT -277.600 4.110 -277.280 4.220 ;
        RECT -278.100 3.970 -277.280 4.110 ;
        RECT -277.600 3.940 -277.280 3.970 ;
        RECT -274.920 4.110 -274.600 4.220 ;
        RECT -274.260 4.110 -274.100 4.900 ;
        RECT -272.660 4.750 -272.320 4.900 ;
        RECT -269.960 4.900 -268.020 5.050 ;
        RECT -269.960 4.750 -269.620 4.900 ;
        RECT -272.640 4.550 -272.320 4.580 ;
        RECT -274.920 3.970 -274.100 4.110 ;
        RECT -273.140 4.410 -272.320 4.550 ;
        RECT -274.920 3.940 -274.600 3.970 ;
        RECT -277.620 3.620 -277.280 3.770 ;
        RECT -279.220 3.470 -277.280 3.620 ;
        RECT -274.920 3.620 -274.580 3.770 ;
        RECT -273.140 3.620 -272.980 4.410 ;
        RECT -272.640 4.300 -272.320 4.410 ;
        RECT -269.960 4.550 -269.640 4.580 ;
        RECT -269.960 4.410 -269.140 4.550 ;
        RECT -269.960 4.300 -269.640 4.410 ;
        RECT -274.920 3.470 -272.980 3.620 ;
        RECT -269.300 3.620 -269.140 4.410 ;
        RECT -268.180 4.110 -268.020 4.900 ;
        RECT -264.340 4.900 -262.400 5.050 ;
        RECT -267.680 4.110 -267.360 4.220 ;
        RECT -268.180 3.970 -267.360 4.110 ;
        RECT -267.680 3.940 -267.360 3.970 ;
        RECT -265.000 4.110 -264.680 4.220 ;
        RECT -264.340 4.110 -264.180 4.900 ;
        RECT -262.740 4.750 -262.400 4.900 ;
        RECT -260.040 4.900 -258.100 5.050 ;
        RECT -260.040 4.750 -259.700 4.900 ;
        RECT -262.720 4.550 -262.400 4.580 ;
        RECT -265.000 3.970 -264.180 4.110 ;
        RECT -263.220 4.410 -262.400 4.550 ;
        RECT -265.000 3.940 -264.680 3.970 ;
        RECT -267.700 3.620 -267.360 3.770 ;
        RECT -269.300 3.470 -267.360 3.620 ;
        RECT -265.000 3.620 -264.660 3.770 ;
        RECT -263.220 3.620 -263.060 4.410 ;
        RECT -262.720 4.300 -262.400 4.410 ;
        RECT -260.040 4.550 -259.720 4.580 ;
        RECT -260.040 4.410 -259.220 4.550 ;
        RECT -260.040 4.300 -259.720 4.410 ;
        RECT -265.000 3.470 -263.060 3.620 ;
        RECT -259.380 3.620 -259.220 4.410 ;
        RECT -258.260 4.110 -258.100 4.900 ;
        RECT -254.420 4.900 -252.480 5.050 ;
        RECT -257.760 4.110 -257.440 4.220 ;
        RECT -258.260 3.970 -257.440 4.110 ;
        RECT -257.760 3.940 -257.440 3.970 ;
        RECT -255.080 4.110 -254.760 4.220 ;
        RECT -254.420 4.110 -254.260 4.900 ;
        RECT -252.820 4.750 -252.480 4.900 ;
        RECT -250.120 4.900 -248.180 5.050 ;
        RECT -250.120 4.750 -249.780 4.900 ;
        RECT -252.800 4.550 -252.480 4.580 ;
        RECT -255.080 3.970 -254.260 4.110 ;
        RECT -253.300 4.410 -252.480 4.550 ;
        RECT -255.080 3.940 -254.760 3.970 ;
        RECT -257.780 3.620 -257.440 3.770 ;
        RECT -259.380 3.470 -257.440 3.620 ;
        RECT -255.080 3.620 -254.740 3.770 ;
        RECT -253.300 3.620 -253.140 4.410 ;
        RECT -252.800 4.300 -252.480 4.410 ;
        RECT -250.120 4.550 -249.800 4.580 ;
        RECT -250.120 4.410 -249.300 4.550 ;
        RECT -250.120 4.300 -249.800 4.410 ;
        RECT -255.080 3.470 -253.140 3.620 ;
        RECT -249.460 3.620 -249.300 4.410 ;
        RECT -248.340 4.110 -248.180 4.900 ;
        RECT -244.500 4.900 -242.560 5.050 ;
        RECT -247.840 4.110 -247.520 4.220 ;
        RECT -248.340 3.970 -247.520 4.110 ;
        RECT -247.840 3.940 -247.520 3.970 ;
        RECT -245.160 4.110 -244.840 4.220 ;
        RECT -244.500 4.110 -244.340 4.900 ;
        RECT -242.900 4.750 -242.560 4.900 ;
        RECT -240.200 4.900 -238.260 5.050 ;
        RECT -240.200 4.750 -239.860 4.900 ;
        RECT -242.880 4.550 -242.560 4.580 ;
        RECT -245.160 3.970 -244.340 4.110 ;
        RECT -243.380 4.410 -242.560 4.550 ;
        RECT -245.160 3.940 -244.840 3.970 ;
        RECT -247.860 3.620 -247.520 3.770 ;
        RECT -249.460 3.470 -247.520 3.620 ;
        RECT -245.160 3.620 -244.820 3.770 ;
        RECT -243.380 3.620 -243.220 4.410 ;
        RECT -242.880 4.300 -242.560 4.410 ;
        RECT -240.200 4.550 -239.880 4.580 ;
        RECT -240.200 4.410 -239.380 4.550 ;
        RECT -240.200 4.300 -239.880 4.410 ;
        RECT -245.160 3.470 -243.220 3.620 ;
        RECT -239.540 3.620 -239.380 4.410 ;
        RECT -238.420 4.110 -238.260 4.900 ;
        RECT -234.580 4.900 -232.640 5.050 ;
        RECT -237.920 4.110 -237.600 4.220 ;
        RECT -238.420 3.970 -237.600 4.110 ;
        RECT -237.920 3.940 -237.600 3.970 ;
        RECT -235.240 4.110 -234.920 4.220 ;
        RECT -234.580 4.110 -234.420 4.900 ;
        RECT -232.980 4.750 -232.640 4.900 ;
        RECT -230.280 4.900 -228.340 5.050 ;
        RECT -230.280 4.750 -229.940 4.900 ;
        RECT -232.960 4.550 -232.640 4.580 ;
        RECT -235.240 3.970 -234.420 4.110 ;
        RECT -233.460 4.410 -232.640 4.550 ;
        RECT -235.240 3.940 -234.920 3.970 ;
        RECT -237.940 3.620 -237.600 3.770 ;
        RECT -239.540 3.470 -237.600 3.620 ;
        RECT -235.240 3.620 -234.900 3.770 ;
        RECT -233.460 3.620 -233.300 4.410 ;
        RECT -232.960 4.300 -232.640 4.410 ;
        RECT -230.280 4.550 -229.960 4.580 ;
        RECT -230.280 4.410 -229.460 4.550 ;
        RECT -230.280 4.300 -229.960 4.410 ;
        RECT -235.240 3.470 -233.300 3.620 ;
        RECT -229.620 3.620 -229.460 4.410 ;
        RECT -228.500 4.110 -228.340 4.900 ;
        RECT -224.660 4.900 -222.720 5.050 ;
        RECT -228.000 4.110 -227.680 4.220 ;
        RECT -228.500 3.970 -227.680 4.110 ;
        RECT -228.000 3.940 -227.680 3.970 ;
        RECT -225.320 4.110 -225.000 4.220 ;
        RECT -224.660 4.110 -224.500 4.900 ;
        RECT -223.060 4.750 -222.720 4.900 ;
        RECT -220.360 4.900 -218.420 5.050 ;
        RECT -220.360 4.750 -220.020 4.900 ;
        RECT -223.040 4.550 -222.720 4.580 ;
        RECT -225.320 3.970 -224.500 4.110 ;
        RECT -223.540 4.410 -222.720 4.550 ;
        RECT -225.320 3.940 -225.000 3.970 ;
        RECT -228.020 3.620 -227.680 3.770 ;
        RECT -229.620 3.470 -227.680 3.620 ;
        RECT -225.320 3.620 -224.980 3.770 ;
        RECT -223.540 3.620 -223.380 4.410 ;
        RECT -223.040 4.300 -222.720 4.410 ;
        RECT -220.360 4.550 -220.040 4.580 ;
        RECT -220.360 4.410 -219.540 4.550 ;
        RECT -220.360 4.300 -220.040 4.410 ;
        RECT -225.320 3.470 -223.380 3.620 ;
        RECT -219.700 3.620 -219.540 4.410 ;
        RECT -218.580 4.110 -218.420 4.900 ;
        RECT -214.740 4.900 -212.800 5.050 ;
        RECT -218.080 4.110 -217.760 4.220 ;
        RECT -218.580 3.970 -217.760 4.110 ;
        RECT -218.080 3.940 -217.760 3.970 ;
        RECT -215.400 4.110 -215.080 4.220 ;
        RECT -214.740 4.110 -214.580 4.900 ;
        RECT -213.140 4.750 -212.800 4.900 ;
        RECT -210.440 4.900 -208.500 5.050 ;
        RECT -210.440 4.750 -210.100 4.900 ;
        RECT -213.120 4.550 -212.800 4.580 ;
        RECT -215.400 3.970 -214.580 4.110 ;
        RECT -213.620 4.410 -212.800 4.550 ;
        RECT -215.400 3.940 -215.080 3.970 ;
        RECT -218.100 3.620 -217.760 3.770 ;
        RECT -219.700 3.470 -217.760 3.620 ;
        RECT -215.400 3.620 -215.060 3.770 ;
        RECT -213.620 3.620 -213.460 4.410 ;
        RECT -213.120 4.300 -212.800 4.410 ;
        RECT -210.440 4.550 -210.120 4.580 ;
        RECT -210.440 4.410 -209.620 4.550 ;
        RECT -210.440 4.300 -210.120 4.410 ;
        RECT -215.400 3.470 -213.460 3.620 ;
        RECT -209.780 3.620 -209.620 4.410 ;
        RECT -208.660 4.110 -208.500 4.900 ;
        RECT -204.820 4.900 -202.880 5.050 ;
        RECT -208.160 4.110 -207.840 4.220 ;
        RECT -208.660 3.970 -207.840 4.110 ;
        RECT -208.160 3.940 -207.840 3.970 ;
        RECT -205.480 4.110 -205.160 4.220 ;
        RECT -204.820 4.110 -204.660 4.900 ;
        RECT -203.220 4.750 -202.880 4.900 ;
        RECT -200.520 4.900 -198.580 5.050 ;
        RECT -200.520 4.750 -200.180 4.900 ;
        RECT -203.200 4.550 -202.880 4.580 ;
        RECT -205.480 3.970 -204.660 4.110 ;
        RECT -203.700 4.410 -202.880 4.550 ;
        RECT -205.480 3.940 -205.160 3.970 ;
        RECT -208.180 3.620 -207.840 3.770 ;
        RECT -209.780 3.470 -207.840 3.620 ;
        RECT -205.480 3.620 -205.140 3.770 ;
        RECT -203.700 3.620 -203.540 4.410 ;
        RECT -203.200 4.300 -202.880 4.410 ;
        RECT -200.520 4.550 -200.200 4.580 ;
        RECT -200.520 4.410 -199.700 4.550 ;
        RECT -200.520 4.300 -200.200 4.410 ;
        RECT -205.480 3.470 -203.540 3.620 ;
        RECT -199.860 3.620 -199.700 4.410 ;
        RECT -198.740 4.110 -198.580 4.900 ;
        RECT -194.900 4.900 -192.960 5.050 ;
        RECT -198.240 4.110 -197.920 4.220 ;
        RECT -198.740 3.970 -197.920 4.110 ;
        RECT -198.240 3.940 -197.920 3.970 ;
        RECT -195.560 4.110 -195.240 4.220 ;
        RECT -194.900 4.110 -194.740 4.900 ;
        RECT -193.300 4.750 -192.960 4.900 ;
        RECT -190.600 4.900 -188.660 5.050 ;
        RECT -190.600 4.750 -190.260 4.900 ;
        RECT -193.280 4.550 -192.960 4.580 ;
        RECT -195.560 3.970 -194.740 4.110 ;
        RECT -193.780 4.410 -192.960 4.550 ;
        RECT -195.560 3.940 -195.240 3.970 ;
        RECT -198.260 3.620 -197.920 3.770 ;
        RECT -199.860 3.470 -197.920 3.620 ;
        RECT -195.560 3.620 -195.220 3.770 ;
        RECT -193.780 3.620 -193.620 4.410 ;
        RECT -193.280 4.300 -192.960 4.410 ;
        RECT -190.600 4.550 -190.280 4.580 ;
        RECT -190.600 4.410 -189.780 4.550 ;
        RECT -190.600 4.300 -190.280 4.410 ;
        RECT -195.560 3.470 -193.620 3.620 ;
        RECT -189.940 3.620 -189.780 4.410 ;
        RECT -188.820 4.110 -188.660 4.900 ;
        RECT -184.980 4.900 -183.040 5.050 ;
        RECT -188.320 4.110 -188.000 4.220 ;
        RECT -188.820 3.970 -188.000 4.110 ;
        RECT -188.320 3.940 -188.000 3.970 ;
        RECT -185.640 4.110 -185.320 4.220 ;
        RECT -184.980 4.110 -184.820 4.900 ;
        RECT -183.380 4.750 -183.040 4.900 ;
        RECT -180.680 4.900 -178.740 5.050 ;
        RECT -180.680 4.750 -180.340 4.900 ;
        RECT -183.360 4.550 -183.040 4.580 ;
        RECT -185.640 3.970 -184.820 4.110 ;
        RECT -183.860 4.410 -183.040 4.550 ;
        RECT -185.640 3.940 -185.320 3.970 ;
        RECT -188.340 3.620 -188.000 3.770 ;
        RECT -189.940 3.470 -188.000 3.620 ;
        RECT -185.640 3.620 -185.300 3.770 ;
        RECT -183.860 3.620 -183.700 4.410 ;
        RECT -183.360 4.300 -183.040 4.410 ;
        RECT -180.680 4.550 -180.360 4.580 ;
        RECT -180.680 4.410 -179.860 4.550 ;
        RECT -180.680 4.300 -180.360 4.410 ;
        RECT -185.640 3.470 -183.700 3.620 ;
        RECT -180.020 3.620 -179.860 4.410 ;
        RECT -178.900 4.110 -178.740 4.900 ;
        RECT -175.060 4.900 -173.120 5.050 ;
        RECT -178.400 4.110 -178.080 4.220 ;
        RECT -178.900 3.970 -178.080 4.110 ;
        RECT -178.400 3.940 -178.080 3.970 ;
        RECT -175.720 4.110 -175.400 4.220 ;
        RECT -175.060 4.110 -174.900 4.900 ;
        RECT -173.460 4.750 -173.120 4.900 ;
        RECT -170.760 4.900 -168.820 5.050 ;
        RECT -170.760 4.750 -170.420 4.900 ;
        RECT -173.440 4.550 -173.120 4.580 ;
        RECT -175.720 3.970 -174.900 4.110 ;
        RECT -173.940 4.410 -173.120 4.550 ;
        RECT -175.720 3.940 -175.400 3.970 ;
        RECT -178.420 3.620 -178.080 3.770 ;
        RECT -180.020 3.470 -178.080 3.620 ;
        RECT -175.720 3.620 -175.380 3.770 ;
        RECT -173.940 3.620 -173.780 4.410 ;
        RECT -173.440 4.300 -173.120 4.410 ;
        RECT -170.760 4.550 -170.440 4.580 ;
        RECT -170.760 4.410 -169.940 4.550 ;
        RECT -170.760 4.300 -170.440 4.410 ;
        RECT -175.720 3.470 -173.780 3.620 ;
        RECT -170.100 3.620 -169.940 4.410 ;
        RECT -168.980 4.110 -168.820 4.900 ;
        RECT -165.140 4.900 -163.200 5.050 ;
        RECT -168.480 4.110 -168.160 4.220 ;
        RECT -168.980 3.970 -168.160 4.110 ;
        RECT -168.480 3.940 -168.160 3.970 ;
        RECT -165.800 4.110 -165.480 4.220 ;
        RECT -165.140 4.110 -164.980 4.900 ;
        RECT -163.540 4.750 -163.200 4.900 ;
        RECT -160.840 4.900 -158.900 5.050 ;
        RECT -160.840 4.750 -160.500 4.900 ;
        RECT -163.520 4.550 -163.200 4.580 ;
        RECT -165.800 3.970 -164.980 4.110 ;
        RECT -164.020 4.410 -163.200 4.550 ;
        RECT -165.800 3.940 -165.480 3.970 ;
        RECT -168.500 3.620 -168.160 3.770 ;
        RECT -170.100 3.470 -168.160 3.620 ;
        RECT -165.800 3.620 -165.460 3.770 ;
        RECT -164.020 3.620 -163.860 4.410 ;
        RECT -163.520 4.300 -163.200 4.410 ;
        RECT -160.840 4.550 -160.520 4.580 ;
        RECT -160.840 4.410 -160.020 4.550 ;
        RECT -160.840 4.300 -160.520 4.410 ;
        RECT -165.800 3.470 -163.860 3.620 ;
        RECT -160.180 3.620 -160.020 4.410 ;
        RECT -159.060 4.110 -158.900 4.900 ;
        RECT -155.220 4.900 -153.280 5.050 ;
        RECT -158.560 4.110 -158.240 4.220 ;
        RECT -159.060 3.970 -158.240 4.110 ;
        RECT -158.560 3.940 -158.240 3.970 ;
        RECT -155.880 4.110 -155.560 4.220 ;
        RECT -155.220 4.110 -155.060 4.900 ;
        RECT -153.620 4.750 -153.280 4.900 ;
        RECT -150.920 4.900 -148.980 5.050 ;
        RECT -150.920 4.750 -150.580 4.900 ;
        RECT -153.600 4.550 -153.280 4.580 ;
        RECT -155.880 3.970 -155.060 4.110 ;
        RECT -154.100 4.410 -153.280 4.550 ;
        RECT -155.880 3.940 -155.560 3.970 ;
        RECT -158.580 3.620 -158.240 3.770 ;
        RECT -160.180 3.470 -158.240 3.620 ;
        RECT -155.880 3.620 -155.540 3.770 ;
        RECT -154.100 3.620 -153.940 4.410 ;
        RECT -153.600 4.300 -153.280 4.410 ;
        RECT -150.920 4.550 -150.600 4.580 ;
        RECT -150.920 4.410 -150.100 4.550 ;
        RECT -150.920 4.300 -150.600 4.410 ;
        RECT -155.880 3.470 -153.940 3.620 ;
        RECT -150.260 3.620 -150.100 4.410 ;
        RECT -149.140 4.110 -148.980 4.900 ;
        RECT -145.300 4.900 -143.360 5.050 ;
        RECT -148.640 4.110 -148.320 4.220 ;
        RECT -149.140 3.970 -148.320 4.110 ;
        RECT -148.640 3.940 -148.320 3.970 ;
        RECT -145.960 4.110 -145.640 4.220 ;
        RECT -145.300 4.110 -145.140 4.900 ;
        RECT -143.700 4.750 -143.360 4.900 ;
        RECT -141.000 4.900 -139.060 5.050 ;
        RECT -141.000 4.750 -140.660 4.900 ;
        RECT -143.680 4.550 -143.360 4.580 ;
        RECT -145.960 3.970 -145.140 4.110 ;
        RECT -144.180 4.410 -143.360 4.550 ;
        RECT -145.960 3.940 -145.640 3.970 ;
        RECT -148.660 3.620 -148.320 3.770 ;
        RECT -150.260 3.470 -148.320 3.620 ;
        RECT -145.960 3.620 -145.620 3.770 ;
        RECT -144.180 3.620 -144.020 4.410 ;
        RECT -143.680 4.300 -143.360 4.410 ;
        RECT -141.000 4.550 -140.680 4.580 ;
        RECT -141.000 4.410 -140.180 4.550 ;
        RECT -141.000 4.300 -140.680 4.410 ;
        RECT -145.960 3.470 -144.020 3.620 ;
        RECT -140.340 3.620 -140.180 4.410 ;
        RECT -139.220 4.110 -139.060 4.900 ;
        RECT -135.380 4.900 -133.440 5.050 ;
        RECT -138.720 4.110 -138.400 4.220 ;
        RECT -139.220 3.970 -138.400 4.110 ;
        RECT -138.720 3.940 -138.400 3.970 ;
        RECT -136.040 4.110 -135.720 4.220 ;
        RECT -135.380 4.110 -135.220 4.900 ;
        RECT -133.780 4.750 -133.440 4.900 ;
        RECT -131.080 4.900 -129.140 5.050 ;
        RECT -131.080 4.750 -130.740 4.900 ;
        RECT -133.760 4.550 -133.440 4.580 ;
        RECT -136.040 3.970 -135.220 4.110 ;
        RECT -134.260 4.410 -133.440 4.550 ;
        RECT -136.040 3.940 -135.720 3.970 ;
        RECT -138.740 3.620 -138.400 3.770 ;
        RECT -140.340 3.470 -138.400 3.620 ;
        RECT -136.040 3.620 -135.700 3.770 ;
        RECT -134.260 3.620 -134.100 4.410 ;
        RECT -133.760 4.300 -133.440 4.410 ;
        RECT -131.080 4.550 -130.760 4.580 ;
        RECT -131.080 4.410 -130.260 4.550 ;
        RECT -131.080 4.300 -130.760 4.410 ;
        RECT -136.040 3.470 -134.100 3.620 ;
        RECT -130.420 3.620 -130.260 4.410 ;
        RECT -129.300 4.110 -129.140 4.900 ;
        RECT -125.460 4.900 -123.520 5.050 ;
        RECT -128.800 4.110 -128.480 4.220 ;
        RECT -129.300 3.970 -128.480 4.110 ;
        RECT -128.800 3.940 -128.480 3.970 ;
        RECT -126.120 4.110 -125.800 4.220 ;
        RECT -125.460 4.110 -125.300 4.900 ;
        RECT -123.860 4.750 -123.520 4.900 ;
        RECT -121.160 4.900 -119.220 5.050 ;
        RECT -121.160 4.750 -120.820 4.900 ;
        RECT -123.840 4.550 -123.520 4.580 ;
        RECT -126.120 3.970 -125.300 4.110 ;
        RECT -124.340 4.410 -123.520 4.550 ;
        RECT -126.120 3.940 -125.800 3.970 ;
        RECT -128.820 3.620 -128.480 3.770 ;
        RECT -130.420 3.470 -128.480 3.620 ;
        RECT -126.120 3.620 -125.780 3.770 ;
        RECT -124.340 3.620 -124.180 4.410 ;
        RECT -123.840 4.300 -123.520 4.410 ;
        RECT -121.160 4.550 -120.840 4.580 ;
        RECT -121.160 4.410 -120.340 4.550 ;
        RECT -121.160 4.300 -120.840 4.410 ;
        RECT -126.120 3.470 -124.180 3.620 ;
        RECT -120.500 3.620 -120.340 4.410 ;
        RECT -119.380 4.110 -119.220 4.900 ;
        RECT -115.540 4.900 -113.600 5.050 ;
        RECT -118.880 4.110 -118.560 4.220 ;
        RECT -119.380 3.970 -118.560 4.110 ;
        RECT -118.880 3.940 -118.560 3.970 ;
        RECT -116.200 4.110 -115.880 4.220 ;
        RECT -115.540 4.110 -115.380 4.900 ;
        RECT -113.940 4.750 -113.600 4.900 ;
        RECT -111.240 4.900 -109.300 5.050 ;
        RECT -111.240 4.750 -110.900 4.900 ;
        RECT -113.920 4.550 -113.600 4.580 ;
        RECT -116.200 3.970 -115.380 4.110 ;
        RECT -114.420 4.410 -113.600 4.550 ;
        RECT -116.200 3.940 -115.880 3.970 ;
        RECT -118.900 3.620 -118.560 3.770 ;
        RECT -120.500 3.470 -118.560 3.620 ;
        RECT -116.200 3.620 -115.860 3.770 ;
        RECT -114.420 3.620 -114.260 4.410 ;
        RECT -113.920 4.300 -113.600 4.410 ;
        RECT -111.240 4.550 -110.920 4.580 ;
        RECT -111.240 4.410 -110.420 4.550 ;
        RECT -111.240 4.300 -110.920 4.410 ;
        RECT -116.200 3.470 -114.260 3.620 ;
        RECT -110.580 3.620 -110.420 4.410 ;
        RECT -109.460 4.110 -109.300 4.900 ;
        RECT -105.620 4.900 -103.680 5.050 ;
        RECT -108.960 4.110 -108.640 4.220 ;
        RECT -109.460 3.970 -108.640 4.110 ;
        RECT -108.960 3.940 -108.640 3.970 ;
        RECT -106.280 4.110 -105.960 4.220 ;
        RECT -105.620 4.110 -105.460 4.900 ;
        RECT -104.020 4.750 -103.680 4.900 ;
        RECT -101.320 4.900 -99.380 5.050 ;
        RECT -101.320 4.750 -100.980 4.900 ;
        RECT -104.000 4.550 -103.680 4.580 ;
        RECT -106.280 3.970 -105.460 4.110 ;
        RECT -104.500 4.410 -103.680 4.550 ;
        RECT -106.280 3.940 -105.960 3.970 ;
        RECT -108.980 3.620 -108.640 3.770 ;
        RECT -110.580 3.470 -108.640 3.620 ;
        RECT -106.280 3.620 -105.940 3.770 ;
        RECT -104.500 3.620 -104.340 4.410 ;
        RECT -104.000 4.300 -103.680 4.410 ;
        RECT -101.320 4.550 -101.000 4.580 ;
        RECT -101.320 4.410 -100.500 4.550 ;
        RECT -101.320 4.300 -101.000 4.410 ;
        RECT -106.280 3.470 -104.340 3.620 ;
        RECT -100.660 3.620 -100.500 4.410 ;
        RECT -99.540 4.110 -99.380 4.900 ;
        RECT -95.700 4.900 -93.760 5.050 ;
        RECT -99.040 4.110 -98.720 4.220 ;
        RECT -99.540 3.970 -98.720 4.110 ;
        RECT -99.040 3.940 -98.720 3.970 ;
        RECT -96.360 4.110 -96.040 4.220 ;
        RECT -95.700 4.110 -95.540 4.900 ;
        RECT -94.100 4.750 -93.760 4.900 ;
        RECT -91.400 4.900 -89.460 5.050 ;
        RECT -91.400 4.750 -91.060 4.900 ;
        RECT -94.080 4.550 -93.760 4.580 ;
        RECT -96.360 3.970 -95.540 4.110 ;
        RECT -94.580 4.410 -93.760 4.550 ;
        RECT -96.360 3.940 -96.040 3.970 ;
        RECT -99.060 3.620 -98.720 3.770 ;
        RECT -100.660 3.470 -98.720 3.620 ;
        RECT -96.360 3.620 -96.020 3.770 ;
        RECT -94.580 3.620 -94.420 4.410 ;
        RECT -94.080 4.300 -93.760 4.410 ;
        RECT -91.400 4.550 -91.080 4.580 ;
        RECT -91.400 4.410 -90.580 4.550 ;
        RECT -91.400 4.300 -91.080 4.410 ;
        RECT -96.360 3.470 -94.420 3.620 ;
        RECT -90.740 3.620 -90.580 4.410 ;
        RECT -89.620 4.110 -89.460 4.900 ;
        RECT -85.780 4.900 -83.840 5.050 ;
        RECT -89.120 4.110 -88.800 4.220 ;
        RECT -89.620 3.970 -88.800 4.110 ;
        RECT -89.120 3.940 -88.800 3.970 ;
        RECT -86.440 4.110 -86.120 4.220 ;
        RECT -85.780 4.110 -85.620 4.900 ;
        RECT -84.180 4.750 -83.840 4.900 ;
        RECT -81.480 4.900 -79.540 5.050 ;
        RECT -81.480 4.750 -81.140 4.900 ;
        RECT -84.160 4.550 -83.840 4.580 ;
        RECT -86.440 3.970 -85.620 4.110 ;
        RECT -84.660 4.410 -83.840 4.550 ;
        RECT -86.440 3.940 -86.120 3.970 ;
        RECT -89.140 3.620 -88.800 3.770 ;
        RECT -90.740 3.470 -88.800 3.620 ;
        RECT -86.440 3.620 -86.100 3.770 ;
        RECT -84.660 3.620 -84.500 4.410 ;
        RECT -84.160 4.300 -83.840 4.410 ;
        RECT -81.480 4.550 -81.160 4.580 ;
        RECT -81.480 4.410 -80.660 4.550 ;
        RECT -81.480 4.300 -81.160 4.410 ;
        RECT -86.440 3.470 -84.500 3.620 ;
        RECT -80.820 3.620 -80.660 4.410 ;
        RECT -79.700 4.110 -79.540 4.900 ;
        RECT -75.860 4.900 -73.920 5.050 ;
        RECT -79.200 4.110 -78.880 4.220 ;
        RECT -79.700 3.970 -78.880 4.110 ;
        RECT -79.200 3.940 -78.880 3.970 ;
        RECT -76.520 4.110 -76.200 4.220 ;
        RECT -75.860 4.110 -75.700 4.900 ;
        RECT -74.260 4.750 -73.920 4.900 ;
        RECT -71.560 4.900 -69.620 5.050 ;
        RECT -71.560 4.750 -71.220 4.900 ;
        RECT -74.240 4.550 -73.920 4.580 ;
        RECT -76.520 3.970 -75.700 4.110 ;
        RECT -74.740 4.410 -73.920 4.550 ;
        RECT -76.520 3.940 -76.200 3.970 ;
        RECT -79.220 3.620 -78.880 3.770 ;
        RECT -80.820 3.470 -78.880 3.620 ;
        RECT -76.520 3.620 -76.180 3.770 ;
        RECT -74.740 3.620 -74.580 4.410 ;
        RECT -74.240 4.300 -73.920 4.410 ;
        RECT -71.560 4.550 -71.240 4.580 ;
        RECT -71.560 4.410 -70.740 4.550 ;
        RECT -71.560 4.300 -71.240 4.410 ;
        RECT -76.520 3.470 -74.580 3.620 ;
        RECT -70.900 3.620 -70.740 4.410 ;
        RECT -69.780 4.110 -69.620 4.900 ;
        RECT -65.940 4.900 -64.000 5.050 ;
        RECT -69.280 4.110 -68.960 4.220 ;
        RECT -69.780 3.970 -68.960 4.110 ;
        RECT -69.280 3.940 -68.960 3.970 ;
        RECT -66.600 4.110 -66.280 4.220 ;
        RECT -65.940 4.110 -65.780 4.900 ;
        RECT -64.340 4.750 -64.000 4.900 ;
        RECT -61.640 4.900 -59.700 5.050 ;
        RECT -61.640 4.750 -61.300 4.900 ;
        RECT -64.320 4.550 -64.000 4.580 ;
        RECT -66.600 3.970 -65.780 4.110 ;
        RECT -64.820 4.410 -64.000 4.550 ;
        RECT -66.600 3.940 -66.280 3.970 ;
        RECT -69.300 3.620 -68.960 3.770 ;
        RECT -70.900 3.470 -68.960 3.620 ;
        RECT -66.600 3.620 -66.260 3.770 ;
        RECT -64.820 3.620 -64.660 4.410 ;
        RECT -64.320 4.300 -64.000 4.410 ;
        RECT -61.640 4.550 -61.320 4.580 ;
        RECT -61.640 4.410 -60.820 4.550 ;
        RECT -61.640 4.300 -61.320 4.410 ;
        RECT -66.600 3.470 -64.660 3.620 ;
        RECT -60.980 3.620 -60.820 4.410 ;
        RECT -59.860 4.110 -59.700 4.900 ;
        RECT -56.020 4.900 -54.080 5.050 ;
        RECT -59.360 4.110 -59.040 4.220 ;
        RECT -59.860 3.970 -59.040 4.110 ;
        RECT -59.360 3.940 -59.040 3.970 ;
        RECT -56.680 4.110 -56.360 4.220 ;
        RECT -56.020 4.110 -55.860 4.900 ;
        RECT -54.420 4.750 -54.080 4.900 ;
        RECT -51.720 4.900 -49.780 5.050 ;
        RECT -51.720 4.750 -51.380 4.900 ;
        RECT -54.400 4.550 -54.080 4.580 ;
        RECT -56.680 3.970 -55.860 4.110 ;
        RECT -54.900 4.410 -54.080 4.550 ;
        RECT -56.680 3.940 -56.360 3.970 ;
        RECT -59.380 3.620 -59.040 3.770 ;
        RECT -60.980 3.470 -59.040 3.620 ;
        RECT -56.680 3.620 -56.340 3.770 ;
        RECT -54.900 3.620 -54.740 4.410 ;
        RECT -54.400 4.300 -54.080 4.410 ;
        RECT -51.720 4.550 -51.400 4.580 ;
        RECT -51.720 4.410 -50.900 4.550 ;
        RECT -51.720 4.300 -51.400 4.410 ;
        RECT -56.680 3.470 -54.740 3.620 ;
        RECT -51.060 3.620 -50.900 4.410 ;
        RECT -49.940 4.110 -49.780 4.900 ;
        RECT -46.100 4.900 -44.160 5.050 ;
        RECT -49.440 4.110 -49.120 4.220 ;
        RECT -49.940 3.970 -49.120 4.110 ;
        RECT -49.440 3.940 -49.120 3.970 ;
        RECT -46.760 4.110 -46.440 4.220 ;
        RECT -46.100 4.110 -45.940 4.900 ;
        RECT -44.500 4.750 -44.160 4.900 ;
        RECT -41.800 4.900 -39.860 5.050 ;
        RECT -41.800 4.750 -41.460 4.900 ;
        RECT -44.480 4.550 -44.160 4.580 ;
        RECT -46.760 3.970 -45.940 4.110 ;
        RECT -44.980 4.410 -44.160 4.550 ;
        RECT -46.760 3.940 -46.440 3.970 ;
        RECT -49.460 3.620 -49.120 3.770 ;
        RECT -51.060 3.470 -49.120 3.620 ;
        RECT -46.760 3.620 -46.420 3.770 ;
        RECT -44.980 3.620 -44.820 4.410 ;
        RECT -44.480 4.300 -44.160 4.410 ;
        RECT -41.800 4.550 -41.480 4.580 ;
        RECT -41.800 4.410 -40.980 4.550 ;
        RECT -41.800 4.300 -41.480 4.410 ;
        RECT -46.760 3.470 -44.820 3.620 ;
        RECT -41.140 3.620 -40.980 4.410 ;
        RECT -40.020 4.110 -39.860 4.900 ;
        RECT -36.180 4.900 -34.240 5.050 ;
        RECT -39.520 4.110 -39.200 4.220 ;
        RECT -40.020 3.970 -39.200 4.110 ;
        RECT -39.520 3.940 -39.200 3.970 ;
        RECT -36.840 4.110 -36.520 4.220 ;
        RECT -36.180 4.110 -36.020 4.900 ;
        RECT -34.580 4.750 -34.240 4.900 ;
        RECT -31.880 4.900 -29.940 5.050 ;
        RECT -31.880 4.750 -31.540 4.900 ;
        RECT -34.560 4.550 -34.240 4.580 ;
        RECT -36.840 3.970 -36.020 4.110 ;
        RECT -35.060 4.410 -34.240 4.550 ;
        RECT -36.840 3.940 -36.520 3.970 ;
        RECT -39.540 3.620 -39.200 3.770 ;
        RECT -41.140 3.470 -39.200 3.620 ;
        RECT -36.840 3.620 -36.500 3.770 ;
        RECT -35.060 3.620 -34.900 4.410 ;
        RECT -34.560 4.300 -34.240 4.410 ;
        RECT -31.880 4.550 -31.560 4.580 ;
        RECT -31.880 4.410 -31.060 4.550 ;
        RECT -31.880 4.300 -31.560 4.410 ;
        RECT -36.840 3.470 -34.900 3.620 ;
        RECT -31.220 3.620 -31.060 4.410 ;
        RECT -30.100 4.110 -29.940 4.900 ;
        RECT -26.260 4.900 -24.320 5.050 ;
        RECT -29.600 4.110 -29.280 4.220 ;
        RECT -30.100 3.970 -29.280 4.110 ;
        RECT -29.600 3.940 -29.280 3.970 ;
        RECT -26.920 4.110 -26.600 4.220 ;
        RECT -26.260 4.110 -26.100 4.900 ;
        RECT -24.660 4.750 -24.320 4.900 ;
        RECT -21.960 4.900 -20.020 5.050 ;
        RECT -21.960 4.750 -21.620 4.900 ;
        RECT -24.640 4.550 -24.320 4.580 ;
        RECT -26.920 3.970 -26.100 4.110 ;
        RECT -25.140 4.410 -24.320 4.550 ;
        RECT -26.920 3.940 -26.600 3.970 ;
        RECT -29.620 3.620 -29.280 3.770 ;
        RECT -31.220 3.470 -29.280 3.620 ;
        RECT -26.920 3.620 -26.580 3.770 ;
        RECT -25.140 3.620 -24.980 4.410 ;
        RECT -24.640 4.300 -24.320 4.410 ;
        RECT -21.960 4.550 -21.640 4.580 ;
        RECT -21.960 4.410 -21.140 4.550 ;
        RECT -21.960 4.300 -21.640 4.410 ;
        RECT -26.920 3.470 -24.980 3.620 ;
        RECT -21.300 3.620 -21.140 4.410 ;
        RECT -20.180 4.110 -20.020 4.900 ;
        RECT -16.340 4.900 -14.400 5.050 ;
        RECT -19.680 4.110 -19.360 4.220 ;
        RECT -20.180 3.970 -19.360 4.110 ;
        RECT -19.680 3.940 -19.360 3.970 ;
        RECT -17.000 4.110 -16.680 4.220 ;
        RECT -16.340 4.110 -16.180 4.900 ;
        RECT -14.740 4.750 -14.400 4.900 ;
        RECT -12.040 4.900 -10.100 5.050 ;
        RECT -12.040 4.750 -11.700 4.900 ;
        RECT -14.720 4.550 -14.400 4.580 ;
        RECT -17.000 3.970 -16.180 4.110 ;
        RECT -15.220 4.410 -14.400 4.550 ;
        RECT -17.000 3.940 -16.680 3.970 ;
        RECT -19.700 3.620 -19.360 3.770 ;
        RECT -21.300 3.470 -19.360 3.620 ;
        RECT -17.000 3.620 -16.660 3.770 ;
        RECT -15.220 3.620 -15.060 4.410 ;
        RECT -14.720 4.300 -14.400 4.410 ;
        RECT -12.040 4.550 -11.720 4.580 ;
        RECT -12.040 4.410 -11.220 4.550 ;
        RECT -12.040 4.300 -11.720 4.410 ;
        RECT -17.000 3.470 -15.060 3.620 ;
        RECT -11.380 3.620 -11.220 4.410 ;
        RECT -10.260 4.110 -10.100 4.900 ;
        RECT -6.420 4.900 -4.480 5.050 ;
        RECT -9.760 4.110 -9.440 4.220 ;
        RECT -10.260 3.970 -9.440 4.110 ;
        RECT -9.760 3.940 -9.440 3.970 ;
        RECT -7.080 4.110 -6.760 4.220 ;
        RECT -6.420 4.110 -6.260 4.900 ;
        RECT -4.820 4.750 -4.480 4.900 ;
        RECT -2.120 4.900 -0.180 5.050 ;
        RECT -2.120 4.750 -1.780 4.900 ;
        RECT -4.800 4.550 -4.480 4.580 ;
        RECT -7.080 3.970 -6.260 4.110 ;
        RECT -5.300 4.410 -4.480 4.550 ;
        RECT -7.080 3.940 -6.760 3.970 ;
        RECT -9.780 3.620 -9.440 3.770 ;
        RECT -11.380 3.470 -9.440 3.620 ;
        RECT -7.080 3.620 -6.740 3.770 ;
        RECT -5.300 3.620 -5.140 4.410 ;
        RECT -4.800 4.300 -4.480 4.410 ;
        RECT -2.120 4.550 -1.800 4.580 ;
        RECT -2.120 4.410 -1.300 4.550 ;
        RECT -2.120 4.300 -1.800 4.410 ;
        RECT -7.080 3.470 -5.140 3.620 ;
        RECT -1.460 3.620 -1.300 4.410 ;
        RECT -0.340 4.110 -0.180 4.900 ;
        RECT 3.500 4.900 5.440 5.050 ;
        RECT 0.160 4.110 0.480 4.220 ;
        RECT -0.340 3.970 0.480 4.110 ;
        RECT 0.160 3.940 0.480 3.970 ;
        RECT 2.840 4.110 3.160 4.220 ;
        RECT 3.500 4.110 3.660 4.900 ;
        RECT 5.100 4.750 5.440 4.900 ;
        RECT 7.800 4.900 9.740 5.050 ;
        RECT 7.800 4.750 8.140 4.900 ;
        RECT 5.120 4.550 5.440 4.580 ;
        RECT 2.840 3.970 3.660 4.110 ;
        RECT 4.620 4.410 5.440 4.550 ;
        RECT 2.840 3.940 3.160 3.970 ;
        RECT 0.140 3.620 0.480 3.770 ;
        RECT -1.460 3.470 0.480 3.620 ;
        RECT 2.840 3.620 3.180 3.770 ;
        RECT 4.620 3.620 4.780 4.410 ;
        RECT 5.120 4.300 5.440 4.410 ;
        RECT 7.800 4.550 8.120 4.580 ;
        RECT 7.800 4.410 8.620 4.550 ;
        RECT 7.800 4.300 8.120 4.410 ;
        RECT 2.840 3.470 4.780 3.620 ;
        RECT 8.460 3.620 8.620 4.410 ;
        RECT 9.580 4.110 9.740 4.900 ;
        RECT 13.420 4.900 15.360 5.050 ;
        RECT 10.080 4.110 10.400 4.220 ;
        RECT 9.580 3.970 10.400 4.110 ;
        RECT 10.080 3.940 10.400 3.970 ;
        RECT 12.760 4.110 13.080 4.220 ;
        RECT 13.420 4.110 13.580 4.900 ;
        RECT 15.020 4.750 15.360 4.900 ;
        RECT 17.720 4.900 19.660 5.050 ;
        RECT 17.720 4.750 18.060 4.900 ;
        RECT 15.040 4.550 15.360 4.580 ;
        RECT 12.760 3.970 13.580 4.110 ;
        RECT 14.540 4.410 15.360 4.550 ;
        RECT 12.760 3.940 13.080 3.970 ;
        RECT 10.060 3.620 10.400 3.770 ;
        RECT 8.460 3.470 10.400 3.620 ;
        RECT 12.760 3.620 13.100 3.770 ;
        RECT 14.540 3.620 14.700 4.410 ;
        RECT 15.040 4.300 15.360 4.410 ;
        RECT 17.720 4.550 18.040 4.580 ;
        RECT 17.720 4.410 18.540 4.550 ;
        RECT 17.720 4.300 18.040 4.410 ;
        RECT 12.760 3.470 14.700 3.620 ;
        RECT 18.380 3.620 18.540 4.410 ;
        RECT 19.500 4.110 19.660 4.900 ;
        RECT 23.340 4.900 25.280 5.050 ;
        RECT 20.000 4.110 20.320 4.220 ;
        RECT 19.500 3.970 20.320 4.110 ;
        RECT 20.000 3.940 20.320 3.970 ;
        RECT 22.680 4.110 23.000 4.220 ;
        RECT 23.340 4.110 23.500 4.900 ;
        RECT 24.940 4.750 25.280 4.900 ;
        RECT 24.960 4.550 25.280 4.580 ;
        RECT 22.680 3.970 23.500 4.110 ;
        RECT 24.460 4.410 25.280 4.550 ;
        RECT 22.680 3.940 23.000 3.970 ;
        RECT 19.980 3.620 20.320 3.770 ;
        RECT 18.380 3.470 20.320 3.620 ;
        RECT 22.680 3.620 23.020 3.770 ;
        RECT 24.460 3.620 24.620 4.410 ;
        RECT 24.960 4.300 25.280 4.410 ;
        RECT 22.680 3.470 24.620 3.620 ;
        RECT -291.210 2.660 -289.370 3.140 ;
        RECT -289.450 1.570 -288.970 2.470 ;
        RECT -288.150 2.340 -287.960 3.470 ;
        RECT -284.080 2.340 -283.890 3.470 ;
        RECT -278.230 2.340 -278.040 3.470 ;
        RECT -274.160 2.340 -273.970 3.470 ;
        RECT -268.310 2.340 -268.120 3.470 ;
        RECT -264.240 2.340 -264.050 3.470 ;
        RECT -258.390 2.340 -258.200 3.470 ;
        RECT -254.320 2.340 -254.130 3.470 ;
        RECT -248.470 2.340 -248.280 3.470 ;
        RECT -244.400 2.340 -244.210 3.470 ;
        RECT -238.550 2.340 -238.360 3.470 ;
        RECT -234.480 2.340 -234.290 3.470 ;
        RECT -228.630 2.340 -228.440 3.470 ;
        RECT -224.560 2.340 -224.370 3.470 ;
        RECT -218.710 2.340 -218.520 3.470 ;
        RECT -214.640 2.340 -214.450 3.470 ;
        RECT -208.790 2.340 -208.600 3.470 ;
        RECT -204.720 2.340 -204.530 3.470 ;
        RECT -198.870 2.340 -198.680 3.470 ;
        RECT -194.800 2.340 -194.610 3.470 ;
        RECT -188.950 2.340 -188.760 3.470 ;
        RECT -184.880 2.340 -184.690 3.470 ;
        RECT -179.030 2.340 -178.840 3.470 ;
        RECT -174.960 2.340 -174.770 3.470 ;
        RECT -169.110 2.340 -168.920 3.470 ;
        RECT -165.040 2.340 -164.850 3.470 ;
        RECT -159.190 2.340 -159.000 3.470 ;
        RECT -155.120 2.340 -154.930 3.470 ;
        RECT -149.270 2.340 -149.080 3.470 ;
        RECT -145.200 2.340 -145.010 3.470 ;
        RECT -139.350 2.340 -139.160 3.470 ;
        RECT -135.280 2.340 -135.090 3.470 ;
        RECT -129.430 2.340 -129.240 3.470 ;
        RECT -125.360 2.340 -125.170 3.470 ;
        RECT -119.510 2.340 -119.320 3.470 ;
        RECT -115.440 2.340 -115.250 3.470 ;
        RECT -109.590 2.340 -109.400 3.470 ;
        RECT -105.520 2.340 -105.330 3.470 ;
        RECT -99.670 2.340 -99.480 3.470 ;
        RECT -95.600 2.340 -95.410 3.470 ;
        RECT -89.750 2.340 -89.560 3.470 ;
        RECT -85.680 2.340 -85.490 3.470 ;
        RECT -79.830 2.340 -79.640 3.470 ;
        RECT -75.760 2.340 -75.570 3.470 ;
        RECT -69.910 2.340 -69.720 3.470 ;
        RECT -65.840 2.340 -65.650 3.470 ;
        RECT -59.990 2.340 -59.800 3.470 ;
        RECT -55.920 2.340 -55.730 3.470 ;
        RECT -50.070 2.340 -49.880 3.470 ;
        RECT -46.000 2.340 -45.810 3.470 ;
        RECT -40.150 2.340 -39.960 3.470 ;
        RECT -36.080 2.340 -35.890 3.470 ;
        RECT -30.230 2.340 -30.040 3.470 ;
        RECT -26.160 2.340 -25.970 3.470 ;
        RECT -20.310 2.340 -20.120 3.470 ;
        RECT -16.240 2.340 -16.050 3.470 ;
        RECT -10.390 2.340 -10.200 3.470 ;
        RECT -6.320 2.340 -6.130 3.470 ;
        RECT -0.470 2.340 -0.280 3.470 ;
        RECT 3.600 2.340 3.790 3.470 ;
        RECT 9.450 2.340 9.640 3.470 ;
        RECT 13.520 2.340 13.710 3.470 ;
        RECT 19.370 2.340 19.560 3.470 ;
        RECT 23.440 2.340 23.630 3.470 ;
        RECT -288.200 2.050 -287.880 2.340 ;
        RECT -284.160 2.050 -283.840 2.340 ;
        RECT -278.280 2.050 -277.960 2.340 ;
        RECT -274.240 2.050 -273.920 2.340 ;
        RECT -268.360 2.050 -268.040 2.340 ;
        RECT -264.320 2.050 -264.000 2.340 ;
        RECT -258.440 2.050 -258.120 2.340 ;
        RECT -254.400 2.050 -254.080 2.340 ;
        RECT -248.520 2.050 -248.200 2.340 ;
        RECT -244.480 2.050 -244.160 2.340 ;
        RECT -238.600 2.050 -238.280 2.340 ;
        RECT -234.560 2.050 -234.240 2.340 ;
        RECT -228.680 2.050 -228.360 2.340 ;
        RECT -224.640 2.050 -224.320 2.340 ;
        RECT -218.760 2.050 -218.440 2.340 ;
        RECT -214.720 2.050 -214.400 2.340 ;
        RECT -208.840 2.050 -208.520 2.340 ;
        RECT -204.800 2.050 -204.480 2.340 ;
        RECT -198.920 2.050 -198.600 2.340 ;
        RECT -194.880 2.050 -194.560 2.340 ;
        RECT -189.000 2.050 -188.680 2.340 ;
        RECT -184.960 2.050 -184.640 2.340 ;
        RECT -179.080 2.050 -178.760 2.340 ;
        RECT -175.040 2.050 -174.720 2.340 ;
        RECT -169.160 2.050 -168.840 2.340 ;
        RECT -165.120 2.050 -164.800 2.340 ;
        RECT -159.240 2.050 -158.920 2.340 ;
        RECT -155.200 2.050 -154.880 2.340 ;
        RECT -149.320 2.050 -149.000 2.340 ;
        RECT -145.280 2.050 -144.960 2.340 ;
        RECT -139.400 2.050 -139.080 2.340 ;
        RECT -135.360 2.050 -135.040 2.340 ;
        RECT -129.480 2.050 -129.160 2.340 ;
        RECT -125.440 2.050 -125.120 2.340 ;
        RECT -119.560 2.050 -119.240 2.340 ;
        RECT -115.520 2.050 -115.200 2.340 ;
        RECT -109.640 2.050 -109.320 2.340 ;
        RECT -105.600 2.050 -105.280 2.340 ;
        RECT -99.720 2.050 -99.400 2.340 ;
        RECT -95.680 2.050 -95.360 2.340 ;
        RECT -89.800 2.050 -89.480 2.340 ;
        RECT -85.760 2.050 -85.440 2.340 ;
        RECT -79.880 2.050 -79.560 2.340 ;
        RECT -75.840 2.050 -75.520 2.340 ;
        RECT -69.960 2.050 -69.640 2.340 ;
        RECT -65.920 2.050 -65.600 2.340 ;
        RECT -60.040 2.050 -59.720 2.340 ;
        RECT -56.000 2.050 -55.680 2.340 ;
        RECT -50.120 2.050 -49.800 2.340 ;
        RECT -46.080 2.050 -45.760 2.340 ;
        RECT -40.200 2.050 -39.880 2.340 ;
        RECT -36.160 2.050 -35.840 2.340 ;
        RECT -30.280 2.050 -29.960 2.340 ;
        RECT -26.240 2.050 -25.920 2.340 ;
        RECT -20.360 2.050 -20.040 2.340 ;
        RECT -16.320 2.050 -16.000 2.340 ;
        RECT -10.440 2.050 -10.120 2.340 ;
        RECT -6.400 2.050 -6.080 2.340 ;
        RECT -0.520 2.050 -0.200 2.340 ;
        RECT 3.520 2.050 3.840 2.340 ;
        RECT 9.400 2.050 9.720 2.340 ;
        RECT 13.440 2.050 13.760 2.340 ;
        RECT 19.320 2.050 19.640 2.340 ;
        RECT 23.360 2.050 23.680 2.340 ;
        RECT -289.910 1.090 -288.970 1.570 ;
        RECT 24.450 1.570 24.930 2.470 ;
        RECT -284.900 1.170 -283.210 1.470 ;
        RECT -274.980 1.170 -273.290 1.470 ;
        RECT -265.060 1.170 -263.370 1.470 ;
        RECT -255.140 1.170 -253.450 1.470 ;
        RECT -245.220 1.170 -243.530 1.470 ;
        RECT -235.300 1.170 -233.610 1.470 ;
        RECT -225.380 1.170 -223.690 1.470 ;
        RECT -215.460 1.170 -213.770 1.470 ;
        RECT -205.540 1.170 -203.850 1.470 ;
        RECT -195.620 1.170 -193.930 1.470 ;
        RECT -185.700 1.170 -184.010 1.470 ;
        RECT -175.780 1.170 -174.090 1.470 ;
        RECT -165.860 1.170 -164.170 1.470 ;
        RECT -155.940 1.170 -154.250 1.470 ;
        RECT -146.020 1.170 -144.330 1.470 ;
        RECT -136.100 1.170 -134.410 1.470 ;
        RECT -126.180 1.170 -124.490 1.470 ;
        RECT -116.260 1.170 -114.570 1.470 ;
        RECT -106.340 1.170 -104.650 1.470 ;
        RECT -96.420 1.170 -94.730 1.470 ;
        RECT -86.500 1.170 -84.810 1.470 ;
        RECT -76.580 1.170 -74.890 1.470 ;
        RECT -66.660 1.170 -64.970 1.470 ;
        RECT -56.740 1.170 -55.050 1.470 ;
        RECT -46.820 1.170 -45.130 1.470 ;
        RECT -36.900 1.170 -35.210 1.470 ;
        RECT -26.980 1.170 -25.290 1.470 ;
        RECT -17.060 1.170 -15.370 1.470 ;
        RECT -7.140 1.170 -5.450 1.470 ;
        RECT 2.780 1.170 4.470 1.470 ;
        RECT 12.700 1.170 14.390 1.470 ;
        RECT 22.620 1.170 24.310 1.470 ;
        RECT -284.390 0.470 -283.390 1.170 ;
        RECT -274.470 0.470 -273.470 1.170 ;
        RECT -264.550 0.470 -263.550 1.170 ;
        RECT -254.630 0.470 -253.630 1.170 ;
        RECT -244.710 0.470 -243.710 1.170 ;
        RECT -234.790 0.470 -233.790 1.170 ;
        RECT -224.870 0.470 -223.870 1.170 ;
        RECT -214.950 0.470 -213.950 1.170 ;
        RECT -205.030 0.470 -204.030 1.170 ;
        RECT -195.110 0.470 -194.110 1.170 ;
        RECT -185.190 0.470 -184.190 1.170 ;
        RECT -175.270 0.470 -174.270 1.170 ;
        RECT -165.350 0.470 -164.350 1.170 ;
        RECT -155.430 0.470 -154.430 1.170 ;
        RECT -145.510 0.470 -144.510 1.170 ;
        RECT -135.590 0.470 -134.590 1.170 ;
        RECT -125.670 0.470 -124.670 1.170 ;
        RECT -115.750 0.470 -114.750 1.170 ;
        RECT -105.830 0.470 -104.830 1.170 ;
        RECT -95.910 0.470 -94.910 1.170 ;
        RECT -85.990 0.470 -84.990 1.170 ;
        RECT -76.070 0.470 -75.070 1.170 ;
        RECT -66.150 0.470 -65.150 1.170 ;
        RECT -56.230 0.470 -55.230 1.170 ;
        RECT -46.310 0.470 -45.310 1.170 ;
        RECT -36.390 0.470 -35.390 1.170 ;
        RECT -26.470 0.470 -25.470 1.170 ;
        RECT -16.550 0.470 -15.550 1.170 ;
        RECT -6.630 0.470 -5.630 1.170 ;
        RECT 3.290 0.470 4.290 1.170 ;
        RECT 13.210 0.470 14.210 1.170 ;
        RECT 23.130 0.470 24.130 1.170 ;
        RECT 24.450 1.090 25.390 1.570 ;
        RECT -289.450 -85.920 -288.990 -85.915 ;
        RECT -289.450 -86.395 -288.510 -85.920 ;
        RECT -287.590 -86.000 -286.590 -85.300 ;
        RECT -277.670 -86.000 -276.670 -85.300 ;
        RECT -267.750 -86.000 -266.750 -85.300 ;
        RECT -257.830 -86.000 -256.830 -85.300 ;
        RECT -247.910 -86.000 -246.910 -85.300 ;
        RECT -237.990 -86.000 -236.990 -85.300 ;
        RECT -228.070 -86.000 -227.070 -85.300 ;
        RECT -218.150 -86.000 -217.150 -85.300 ;
        RECT -208.230 -86.000 -207.230 -85.300 ;
        RECT -198.310 -86.000 -197.310 -85.300 ;
        RECT -188.390 -86.000 -187.390 -85.300 ;
        RECT -178.470 -86.000 -177.470 -85.300 ;
        RECT -168.550 -86.000 -167.550 -85.300 ;
        RECT -158.630 -86.000 -157.630 -85.300 ;
        RECT -148.710 -86.000 -147.710 -85.300 ;
        RECT -138.790 -86.000 -137.790 -85.300 ;
        RECT -128.870 -86.000 -127.870 -85.300 ;
        RECT -118.950 -86.000 -117.950 -85.300 ;
        RECT -109.030 -86.000 -108.030 -85.300 ;
        RECT -99.110 -86.000 -98.110 -85.300 ;
        RECT -89.190 -86.000 -88.190 -85.300 ;
        RECT -79.270 -86.000 -78.270 -85.300 ;
        RECT -69.350 -86.000 -68.350 -85.300 ;
        RECT -59.430 -86.000 -58.430 -85.300 ;
        RECT -49.510 -86.000 -48.510 -85.300 ;
        RECT -39.590 -86.000 -38.590 -85.300 ;
        RECT -29.670 -86.000 -28.670 -85.300 ;
        RECT -19.750 -86.000 -18.750 -85.300 ;
        RECT -9.830 -86.000 -8.830 -85.300 ;
        RECT 0.090 -86.000 1.090 -85.300 ;
        RECT 10.010 -86.000 11.010 -85.300 ;
        RECT 19.930 -86.000 20.930 -85.300 ;
        RECT -288.100 -86.300 -286.410 -86.000 ;
        RECT -278.180 -86.300 -276.490 -86.000 ;
        RECT -268.260 -86.300 -266.570 -86.000 ;
        RECT -258.340 -86.300 -256.650 -86.000 ;
        RECT -248.420 -86.300 -246.730 -86.000 ;
        RECT -238.500 -86.300 -236.810 -86.000 ;
        RECT -228.580 -86.300 -226.890 -86.000 ;
        RECT -218.660 -86.300 -216.970 -86.000 ;
        RECT -208.740 -86.300 -207.050 -86.000 ;
        RECT -198.820 -86.300 -197.130 -86.000 ;
        RECT -188.900 -86.300 -187.210 -86.000 ;
        RECT -178.980 -86.300 -177.290 -86.000 ;
        RECT -169.060 -86.300 -167.370 -86.000 ;
        RECT -159.140 -86.300 -157.450 -86.000 ;
        RECT -149.220 -86.300 -147.530 -86.000 ;
        RECT -139.300 -86.300 -137.610 -86.000 ;
        RECT -129.380 -86.300 -127.690 -86.000 ;
        RECT -119.460 -86.300 -117.770 -86.000 ;
        RECT -109.540 -86.300 -107.850 -86.000 ;
        RECT -99.620 -86.300 -97.930 -86.000 ;
        RECT -89.700 -86.300 -88.010 -86.000 ;
        RECT -79.780 -86.300 -78.090 -86.000 ;
        RECT -69.860 -86.300 -68.170 -86.000 ;
        RECT -59.940 -86.300 -58.250 -86.000 ;
        RECT -50.020 -86.300 -48.330 -86.000 ;
        RECT -40.100 -86.300 -38.410 -86.000 ;
        RECT -30.180 -86.300 -28.490 -86.000 ;
        RECT -20.260 -86.300 -18.570 -86.000 ;
        RECT -10.340 -86.300 -8.650 -86.000 ;
        RECT -0.420 -86.300 1.270 -86.000 ;
        RECT 9.500 -86.300 11.190 -86.000 ;
        RECT 19.420 -86.300 21.110 -86.000 ;
        RECT -288.990 -87.300 -288.510 -86.395 ;
        RECT -287.360 -87.170 -287.040 -86.880 ;
        RECT -281.480 -87.170 -281.160 -86.880 ;
        RECT -277.440 -87.170 -277.120 -86.880 ;
        RECT -271.560 -87.170 -271.240 -86.880 ;
        RECT -267.520 -87.170 -267.200 -86.880 ;
        RECT -261.640 -87.170 -261.320 -86.880 ;
        RECT -257.600 -87.170 -257.280 -86.880 ;
        RECT -251.720 -87.170 -251.400 -86.880 ;
        RECT -247.680 -87.170 -247.360 -86.880 ;
        RECT -241.800 -87.170 -241.480 -86.880 ;
        RECT -237.760 -87.170 -237.440 -86.880 ;
        RECT -231.880 -87.170 -231.560 -86.880 ;
        RECT -227.840 -87.170 -227.520 -86.880 ;
        RECT -221.960 -87.170 -221.640 -86.880 ;
        RECT -217.920 -87.170 -217.600 -86.880 ;
        RECT -212.040 -87.170 -211.720 -86.880 ;
        RECT -208.000 -87.170 -207.680 -86.880 ;
        RECT -202.120 -87.170 -201.800 -86.880 ;
        RECT -198.080 -87.170 -197.760 -86.880 ;
        RECT -192.200 -87.170 -191.880 -86.880 ;
        RECT -188.160 -87.170 -187.840 -86.880 ;
        RECT -182.280 -87.170 -181.960 -86.880 ;
        RECT -178.240 -87.170 -177.920 -86.880 ;
        RECT -172.360 -87.170 -172.040 -86.880 ;
        RECT -168.320 -87.170 -168.000 -86.880 ;
        RECT -162.440 -87.170 -162.120 -86.880 ;
        RECT -158.400 -87.170 -158.080 -86.880 ;
        RECT -152.520 -87.170 -152.200 -86.880 ;
        RECT -148.480 -87.170 -148.160 -86.880 ;
        RECT -142.600 -87.170 -142.280 -86.880 ;
        RECT -138.560 -87.170 -138.240 -86.880 ;
        RECT -132.680 -87.170 -132.360 -86.880 ;
        RECT -128.640 -87.170 -128.320 -86.880 ;
        RECT -122.760 -87.170 -122.440 -86.880 ;
        RECT -118.720 -87.170 -118.400 -86.880 ;
        RECT -112.840 -87.170 -112.520 -86.880 ;
        RECT -108.800 -87.170 -108.480 -86.880 ;
        RECT -102.920 -87.170 -102.600 -86.880 ;
        RECT -98.880 -87.170 -98.560 -86.880 ;
        RECT -93.000 -87.170 -92.680 -86.880 ;
        RECT -88.960 -87.170 -88.640 -86.880 ;
        RECT -83.080 -87.170 -82.760 -86.880 ;
        RECT -79.040 -87.170 -78.720 -86.880 ;
        RECT -73.160 -87.170 -72.840 -86.880 ;
        RECT -69.120 -87.170 -68.800 -86.880 ;
        RECT -63.240 -87.170 -62.920 -86.880 ;
        RECT -59.200 -87.170 -58.880 -86.880 ;
        RECT -53.320 -87.170 -53.000 -86.880 ;
        RECT -49.280 -87.170 -48.960 -86.880 ;
        RECT -43.400 -87.170 -43.080 -86.880 ;
        RECT -39.360 -87.170 -39.040 -86.880 ;
        RECT -33.480 -87.170 -33.160 -86.880 ;
        RECT -29.440 -87.170 -29.120 -86.880 ;
        RECT -23.560 -87.170 -23.240 -86.880 ;
        RECT -19.520 -87.170 -19.200 -86.880 ;
        RECT -13.640 -87.170 -13.320 -86.880 ;
        RECT -9.600 -87.170 -9.280 -86.880 ;
        RECT -3.720 -87.170 -3.400 -86.880 ;
        RECT 0.320 -87.170 0.640 -86.880 ;
        RECT 6.200 -87.170 6.520 -86.880 ;
        RECT 10.240 -87.170 10.560 -86.880 ;
        RECT 16.120 -87.170 16.440 -86.880 ;
        RECT 20.160 -87.170 20.480 -86.880 ;
        RECT 26.040 -87.170 26.360 -86.880 ;
        RECT -289.450 -87.970 -287.610 -87.490 ;
        RECT -287.280 -88.300 -287.090 -87.170 ;
        RECT -281.430 -88.300 -281.240 -87.170 ;
        RECT -277.360 -88.300 -277.170 -87.170 ;
        RECT -271.510 -88.300 -271.320 -87.170 ;
        RECT -267.440 -88.300 -267.250 -87.170 ;
        RECT -261.590 -88.300 -261.400 -87.170 ;
        RECT -257.520 -88.300 -257.330 -87.170 ;
        RECT -251.670 -88.300 -251.480 -87.170 ;
        RECT -247.600 -88.300 -247.410 -87.170 ;
        RECT -241.750 -88.300 -241.560 -87.170 ;
        RECT -237.680 -88.300 -237.490 -87.170 ;
        RECT -231.830 -88.300 -231.640 -87.170 ;
        RECT -227.760 -88.300 -227.570 -87.170 ;
        RECT -221.910 -88.300 -221.720 -87.170 ;
        RECT -217.840 -88.300 -217.650 -87.170 ;
        RECT -211.990 -88.300 -211.800 -87.170 ;
        RECT -207.920 -88.300 -207.730 -87.170 ;
        RECT -202.070 -88.300 -201.880 -87.170 ;
        RECT -198.000 -88.300 -197.810 -87.170 ;
        RECT -192.150 -88.300 -191.960 -87.170 ;
        RECT -188.080 -88.300 -187.890 -87.170 ;
        RECT -182.230 -88.300 -182.040 -87.170 ;
        RECT -178.160 -88.300 -177.970 -87.170 ;
        RECT -172.310 -88.300 -172.120 -87.170 ;
        RECT -168.240 -88.300 -168.050 -87.170 ;
        RECT -162.390 -88.300 -162.200 -87.170 ;
        RECT -158.320 -88.300 -158.130 -87.170 ;
        RECT -152.470 -88.300 -152.280 -87.170 ;
        RECT -148.400 -88.300 -148.210 -87.170 ;
        RECT -142.550 -88.300 -142.360 -87.170 ;
        RECT -138.480 -88.300 -138.290 -87.170 ;
        RECT -132.630 -88.300 -132.440 -87.170 ;
        RECT -128.560 -88.300 -128.370 -87.170 ;
        RECT -122.710 -88.300 -122.520 -87.170 ;
        RECT -118.640 -88.300 -118.450 -87.170 ;
        RECT -112.790 -88.300 -112.600 -87.170 ;
        RECT -108.720 -88.300 -108.530 -87.170 ;
        RECT -102.870 -88.300 -102.680 -87.170 ;
        RECT -98.800 -88.300 -98.610 -87.170 ;
        RECT -92.950 -88.300 -92.760 -87.170 ;
        RECT -88.880 -88.300 -88.690 -87.170 ;
        RECT -83.030 -88.300 -82.840 -87.170 ;
        RECT -78.960 -88.300 -78.770 -87.170 ;
        RECT -73.110 -88.300 -72.920 -87.170 ;
        RECT -69.040 -88.300 -68.850 -87.170 ;
        RECT -63.190 -88.300 -63.000 -87.170 ;
        RECT -59.120 -88.300 -58.930 -87.170 ;
        RECT -53.270 -88.300 -53.080 -87.170 ;
        RECT -49.200 -88.300 -49.010 -87.170 ;
        RECT -43.350 -88.300 -43.160 -87.170 ;
        RECT -39.280 -88.300 -39.090 -87.170 ;
        RECT -33.430 -88.300 -33.240 -87.170 ;
        RECT -29.360 -88.300 -29.170 -87.170 ;
        RECT -23.510 -88.300 -23.320 -87.170 ;
        RECT -19.440 -88.300 -19.250 -87.170 ;
        RECT -13.590 -88.300 -13.400 -87.170 ;
        RECT -9.520 -88.300 -9.330 -87.170 ;
        RECT -3.670 -88.300 -3.480 -87.170 ;
        RECT 0.400 -88.300 0.590 -87.170 ;
        RECT 6.250 -88.300 6.440 -87.170 ;
        RECT 10.320 -88.300 10.510 -87.170 ;
        RECT 16.170 -88.300 16.360 -87.170 ;
        RECT 20.240 -88.300 20.430 -87.170 ;
        RECT 26.090 -88.300 26.280 -87.170 ;
        RECT 26.610 -87.970 28.450 -87.490 ;
        RECT -288.040 -88.450 -286.100 -88.300 ;
        RECT -288.040 -88.600 -287.700 -88.450 ;
        RECT -288.040 -88.800 -287.720 -88.770 ;
        RECT -288.040 -88.940 -287.220 -88.800 ;
        RECT -288.040 -89.050 -287.720 -88.940 ;
        RECT -287.380 -89.730 -287.220 -88.940 ;
        RECT -286.260 -89.240 -286.100 -88.450 ;
        RECT -282.420 -88.450 -280.480 -88.300 ;
        RECT -285.760 -89.240 -285.440 -89.130 ;
        RECT -286.260 -89.380 -285.440 -89.240 ;
        RECT -285.760 -89.410 -285.440 -89.380 ;
        RECT -283.080 -89.240 -282.760 -89.130 ;
        RECT -282.420 -89.240 -282.260 -88.450 ;
        RECT -280.820 -88.600 -280.480 -88.450 ;
        RECT -278.120 -88.450 -276.180 -88.300 ;
        RECT -278.120 -88.600 -277.780 -88.450 ;
        RECT -280.800 -88.800 -280.480 -88.770 ;
        RECT -283.080 -89.380 -282.260 -89.240 ;
        RECT -281.300 -88.940 -280.480 -88.800 ;
        RECT -283.080 -89.410 -282.760 -89.380 ;
        RECT -285.780 -89.730 -285.440 -89.580 ;
        RECT -287.380 -89.880 -285.440 -89.730 ;
        RECT -283.080 -89.730 -282.740 -89.580 ;
        RECT -281.300 -89.730 -281.140 -88.940 ;
        RECT -280.800 -89.050 -280.480 -88.940 ;
        RECT -278.120 -88.800 -277.800 -88.770 ;
        RECT -278.120 -88.940 -277.300 -88.800 ;
        RECT -278.120 -89.050 -277.800 -88.940 ;
        RECT -283.080 -89.880 -281.140 -89.730 ;
        RECT -277.460 -89.730 -277.300 -88.940 ;
        RECT -276.340 -89.240 -276.180 -88.450 ;
        RECT -272.500 -88.450 -270.560 -88.300 ;
        RECT -275.840 -89.240 -275.520 -89.130 ;
        RECT -276.340 -89.380 -275.520 -89.240 ;
        RECT -275.840 -89.410 -275.520 -89.380 ;
        RECT -273.160 -89.240 -272.840 -89.130 ;
        RECT -272.500 -89.240 -272.340 -88.450 ;
        RECT -270.900 -88.600 -270.560 -88.450 ;
        RECT -268.200 -88.450 -266.260 -88.300 ;
        RECT -268.200 -88.600 -267.860 -88.450 ;
        RECT -270.880 -88.800 -270.560 -88.770 ;
        RECT -273.160 -89.380 -272.340 -89.240 ;
        RECT -271.380 -88.940 -270.560 -88.800 ;
        RECT -273.160 -89.410 -272.840 -89.380 ;
        RECT -275.860 -89.730 -275.520 -89.580 ;
        RECT -277.460 -89.880 -275.520 -89.730 ;
        RECT -273.160 -89.730 -272.820 -89.580 ;
        RECT -271.380 -89.730 -271.220 -88.940 ;
        RECT -270.880 -89.050 -270.560 -88.940 ;
        RECT -268.200 -88.800 -267.880 -88.770 ;
        RECT -268.200 -88.940 -267.380 -88.800 ;
        RECT -268.200 -89.050 -267.880 -88.940 ;
        RECT -273.160 -89.880 -271.220 -89.730 ;
        RECT -267.540 -89.730 -267.380 -88.940 ;
        RECT -266.420 -89.240 -266.260 -88.450 ;
        RECT -262.580 -88.450 -260.640 -88.300 ;
        RECT -265.920 -89.240 -265.600 -89.130 ;
        RECT -266.420 -89.380 -265.600 -89.240 ;
        RECT -265.920 -89.410 -265.600 -89.380 ;
        RECT -263.240 -89.240 -262.920 -89.130 ;
        RECT -262.580 -89.240 -262.420 -88.450 ;
        RECT -260.980 -88.600 -260.640 -88.450 ;
        RECT -258.280 -88.450 -256.340 -88.300 ;
        RECT -258.280 -88.600 -257.940 -88.450 ;
        RECT -260.960 -88.800 -260.640 -88.770 ;
        RECT -263.240 -89.380 -262.420 -89.240 ;
        RECT -261.460 -88.940 -260.640 -88.800 ;
        RECT -263.240 -89.410 -262.920 -89.380 ;
        RECT -265.940 -89.730 -265.600 -89.580 ;
        RECT -267.540 -89.880 -265.600 -89.730 ;
        RECT -263.240 -89.730 -262.900 -89.580 ;
        RECT -261.460 -89.730 -261.300 -88.940 ;
        RECT -260.960 -89.050 -260.640 -88.940 ;
        RECT -258.280 -88.800 -257.960 -88.770 ;
        RECT -258.280 -88.940 -257.460 -88.800 ;
        RECT -258.280 -89.050 -257.960 -88.940 ;
        RECT -263.240 -89.880 -261.300 -89.730 ;
        RECT -257.620 -89.730 -257.460 -88.940 ;
        RECT -256.500 -89.240 -256.340 -88.450 ;
        RECT -252.660 -88.450 -250.720 -88.300 ;
        RECT -256.000 -89.240 -255.680 -89.130 ;
        RECT -256.500 -89.380 -255.680 -89.240 ;
        RECT -256.000 -89.410 -255.680 -89.380 ;
        RECT -253.320 -89.240 -253.000 -89.130 ;
        RECT -252.660 -89.240 -252.500 -88.450 ;
        RECT -251.060 -88.600 -250.720 -88.450 ;
        RECT -248.360 -88.450 -246.420 -88.300 ;
        RECT -248.360 -88.600 -248.020 -88.450 ;
        RECT -251.040 -88.800 -250.720 -88.770 ;
        RECT -253.320 -89.380 -252.500 -89.240 ;
        RECT -251.540 -88.940 -250.720 -88.800 ;
        RECT -253.320 -89.410 -253.000 -89.380 ;
        RECT -256.020 -89.730 -255.680 -89.580 ;
        RECT -257.620 -89.880 -255.680 -89.730 ;
        RECT -253.320 -89.730 -252.980 -89.580 ;
        RECT -251.540 -89.730 -251.380 -88.940 ;
        RECT -251.040 -89.050 -250.720 -88.940 ;
        RECT -248.360 -88.800 -248.040 -88.770 ;
        RECT -248.360 -88.940 -247.540 -88.800 ;
        RECT -248.360 -89.050 -248.040 -88.940 ;
        RECT -253.320 -89.880 -251.380 -89.730 ;
        RECT -247.700 -89.730 -247.540 -88.940 ;
        RECT -246.580 -89.240 -246.420 -88.450 ;
        RECT -242.740 -88.450 -240.800 -88.300 ;
        RECT -246.080 -89.240 -245.760 -89.130 ;
        RECT -246.580 -89.380 -245.760 -89.240 ;
        RECT -246.080 -89.410 -245.760 -89.380 ;
        RECT -243.400 -89.240 -243.080 -89.130 ;
        RECT -242.740 -89.240 -242.580 -88.450 ;
        RECT -241.140 -88.600 -240.800 -88.450 ;
        RECT -238.440 -88.450 -236.500 -88.300 ;
        RECT -238.440 -88.600 -238.100 -88.450 ;
        RECT -241.120 -88.800 -240.800 -88.770 ;
        RECT -243.400 -89.380 -242.580 -89.240 ;
        RECT -241.620 -88.940 -240.800 -88.800 ;
        RECT -243.400 -89.410 -243.080 -89.380 ;
        RECT -246.100 -89.730 -245.760 -89.580 ;
        RECT -247.700 -89.880 -245.760 -89.730 ;
        RECT -243.400 -89.730 -243.060 -89.580 ;
        RECT -241.620 -89.730 -241.460 -88.940 ;
        RECT -241.120 -89.050 -240.800 -88.940 ;
        RECT -238.440 -88.800 -238.120 -88.770 ;
        RECT -238.440 -88.940 -237.620 -88.800 ;
        RECT -238.440 -89.050 -238.120 -88.940 ;
        RECT -243.400 -89.880 -241.460 -89.730 ;
        RECT -237.780 -89.730 -237.620 -88.940 ;
        RECT -236.660 -89.240 -236.500 -88.450 ;
        RECT -232.820 -88.450 -230.880 -88.300 ;
        RECT -236.160 -89.240 -235.840 -89.130 ;
        RECT -236.660 -89.380 -235.840 -89.240 ;
        RECT -236.160 -89.410 -235.840 -89.380 ;
        RECT -233.480 -89.240 -233.160 -89.130 ;
        RECT -232.820 -89.240 -232.660 -88.450 ;
        RECT -231.220 -88.600 -230.880 -88.450 ;
        RECT -228.520 -88.450 -226.580 -88.300 ;
        RECT -228.520 -88.600 -228.180 -88.450 ;
        RECT -231.200 -88.800 -230.880 -88.770 ;
        RECT -233.480 -89.380 -232.660 -89.240 ;
        RECT -231.700 -88.940 -230.880 -88.800 ;
        RECT -233.480 -89.410 -233.160 -89.380 ;
        RECT -236.180 -89.730 -235.840 -89.580 ;
        RECT -237.780 -89.880 -235.840 -89.730 ;
        RECT -233.480 -89.730 -233.140 -89.580 ;
        RECT -231.700 -89.730 -231.540 -88.940 ;
        RECT -231.200 -89.050 -230.880 -88.940 ;
        RECT -228.520 -88.800 -228.200 -88.770 ;
        RECT -228.520 -88.940 -227.700 -88.800 ;
        RECT -228.520 -89.050 -228.200 -88.940 ;
        RECT -233.480 -89.880 -231.540 -89.730 ;
        RECT -227.860 -89.730 -227.700 -88.940 ;
        RECT -226.740 -89.240 -226.580 -88.450 ;
        RECT -222.900 -88.450 -220.960 -88.300 ;
        RECT -226.240 -89.240 -225.920 -89.130 ;
        RECT -226.740 -89.380 -225.920 -89.240 ;
        RECT -226.240 -89.410 -225.920 -89.380 ;
        RECT -223.560 -89.240 -223.240 -89.130 ;
        RECT -222.900 -89.240 -222.740 -88.450 ;
        RECT -221.300 -88.600 -220.960 -88.450 ;
        RECT -218.600 -88.450 -216.660 -88.300 ;
        RECT -218.600 -88.600 -218.260 -88.450 ;
        RECT -221.280 -88.800 -220.960 -88.770 ;
        RECT -223.560 -89.380 -222.740 -89.240 ;
        RECT -221.780 -88.940 -220.960 -88.800 ;
        RECT -223.560 -89.410 -223.240 -89.380 ;
        RECT -226.260 -89.730 -225.920 -89.580 ;
        RECT -227.860 -89.880 -225.920 -89.730 ;
        RECT -223.560 -89.730 -223.220 -89.580 ;
        RECT -221.780 -89.730 -221.620 -88.940 ;
        RECT -221.280 -89.050 -220.960 -88.940 ;
        RECT -218.600 -88.800 -218.280 -88.770 ;
        RECT -218.600 -88.940 -217.780 -88.800 ;
        RECT -218.600 -89.050 -218.280 -88.940 ;
        RECT -223.560 -89.880 -221.620 -89.730 ;
        RECT -217.940 -89.730 -217.780 -88.940 ;
        RECT -216.820 -89.240 -216.660 -88.450 ;
        RECT -212.980 -88.450 -211.040 -88.300 ;
        RECT -216.320 -89.240 -216.000 -89.130 ;
        RECT -216.820 -89.380 -216.000 -89.240 ;
        RECT -216.320 -89.410 -216.000 -89.380 ;
        RECT -213.640 -89.240 -213.320 -89.130 ;
        RECT -212.980 -89.240 -212.820 -88.450 ;
        RECT -211.380 -88.600 -211.040 -88.450 ;
        RECT -208.680 -88.450 -206.740 -88.300 ;
        RECT -208.680 -88.600 -208.340 -88.450 ;
        RECT -211.360 -88.800 -211.040 -88.770 ;
        RECT -213.640 -89.380 -212.820 -89.240 ;
        RECT -211.860 -88.940 -211.040 -88.800 ;
        RECT -213.640 -89.410 -213.320 -89.380 ;
        RECT -216.340 -89.730 -216.000 -89.580 ;
        RECT -217.940 -89.880 -216.000 -89.730 ;
        RECT -213.640 -89.730 -213.300 -89.580 ;
        RECT -211.860 -89.730 -211.700 -88.940 ;
        RECT -211.360 -89.050 -211.040 -88.940 ;
        RECT -208.680 -88.800 -208.360 -88.770 ;
        RECT -208.680 -88.940 -207.860 -88.800 ;
        RECT -208.680 -89.050 -208.360 -88.940 ;
        RECT -213.640 -89.880 -211.700 -89.730 ;
        RECT -208.020 -89.730 -207.860 -88.940 ;
        RECT -206.900 -89.240 -206.740 -88.450 ;
        RECT -203.060 -88.450 -201.120 -88.300 ;
        RECT -206.400 -89.240 -206.080 -89.130 ;
        RECT -206.900 -89.380 -206.080 -89.240 ;
        RECT -206.400 -89.410 -206.080 -89.380 ;
        RECT -203.720 -89.240 -203.400 -89.130 ;
        RECT -203.060 -89.240 -202.900 -88.450 ;
        RECT -201.460 -88.600 -201.120 -88.450 ;
        RECT -198.760 -88.450 -196.820 -88.300 ;
        RECT -198.760 -88.600 -198.420 -88.450 ;
        RECT -201.440 -88.800 -201.120 -88.770 ;
        RECT -203.720 -89.380 -202.900 -89.240 ;
        RECT -201.940 -88.940 -201.120 -88.800 ;
        RECT -203.720 -89.410 -203.400 -89.380 ;
        RECT -206.420 -89.730 -206.080 -89.580 ;
        RECT -208.020 -89.880 -206.080 -89.730 ;
        RECT -203.720 -89.730 -203.380 -89.580 ;
        RECT -201.940 -89.730 -201.780 -88.940 ;
        RECT -201.440 -89.050 -201.120 -88.940 ;
        RECT -198.760 -88.800 -198.440 -88.770 ;
        RECT -198.760 -88.940 -197.940 -88.800 ;
        RECT -198.760 -89.050 -198.440 -88.940 ;
        RECT -203.720 -89.880 -201.780 -89.730 ;
        RECT -198.100 -89.730 -197.940 -88.940 ;
        RECT -196.980 -89.240 -196.820 -88.450 ;
        RECT -193.140 -88.450 -191.200 -88.300 ;
        RECT -196.480 -89.240 -196.160 -89.130 ;
        RECT -196.980 -89.380 -196.160 -89.240 ;
        RECT -196.480 -89.410 -196.160 -89.380 ;
        RECT -193.800 -89.240 -193.480 -89.130 ;
        RECT -193.140 -89.240 -192.980 -88.450 ;
        RECT -191.540 -88.600 -191.200 -88.450 ;
        RECT -188.840 -88.450 -186.900 -88.300 ;
        RECT -188.840 -88.600 -188.500 -88.450 ;
        RECT -191.520 -88.800 -191.200 -88.770 ;
        RECT -193.800 -89.380 -192.980 -89.240 ;
        RECT -192.020 -88.940 -191.200 -88.800 ;
        RECT -193.800 -89.410 -193.480 -89.380 ;
        RECT -196.500 -89.730 -196.160 -89.580 ;
        RECT -198.100 -89.880 -196.160 -89.730 ;
        RECT -193.800 -89.730 -193.460 -89.580 ;
        RECT -192.020 -89.730 -191.860 -88.940 ;
        RECT -191.520 -89.050 -191.200 -88.940 ;
        RECT -188.840 -88.800 -188.520 -88.770 ;
        RECT -188.840 -88.940 -188.020 -88.800 ;
        RECT -188.840 -89.050 -188.520 -88.940 ;
        RECT -193.800 -89.880 -191.860 -89.730 ;
        RECT -188.180 -89.730 -188.020 -88.940 ;
        RECT -187.060 -89.240 -186.900 -88.450 ;
        RECT -183.220 -88.450 -181.280 -88.300 ;
        RECT -186.560 -89.240 -186.240 -89.130 ;
        RECT -187.060 -89.380 -186.240 -89.240 ;
        RECT -186.560 -89.410 -186.240 -89.380 ;
        RECT -183.880 -89.240 -183.560 -89.130 ;
        RECT -183.220 -89.240 -183.060 -88.450 ;
        RECT -181.620 -88.600 -181.280 -88.450 ;
        RECT -178.920 -88.450 -176.980 -88.300 ;
        RECT -178.920 -88.600 -178.580 -88.450 ;
        RECT -181.600 -88.800 -181.280 -88.770 ;
        RECT -183.880 -89.380 -183.060 -89.240 ;
        RECT -182.100 -88.940 -181.280 -88.800 ;
        RECT -183.880 -89.410 -183.560 -89.380 ;
        RECT -186.580 -89.730 -186.240 -89.580 ;
        RECT -188.180 -89.880 -186.240 -89.730 ;
        RECT -183.880 -89.730 -183.540 -89.580 ;
        RECT -182.100 -89.730 -181.940 -88.940 ;
        RECT -181.600 -89.050 -181.280 -88.940 ;
        RECT -178.920 -88.800 -178.600 -88.770 ;
        RECT -178.920 -88.940 -178.100 -88.800 ;
        RECT -178.920 -89.050 -178.600 -88.940 ;
        RECT -183.880 -89.880 -181.940 -89.730 ;
        RECT -178.260 -89.730 -178.100 -88.940 ;
        RECT -177.140 -89.240 -176.980 -88.450 ;
        RECT -173.300 -88.450 -171.360 -88.300 ;
        RECT -176.640 -89.240 -176.320 -89.130 ;
        RECT -177.140 -89.380 -176.320 -89.240 ;
        RECT -176.640 -89.410 -176.320 -89.380 ;
        RECT -173.960 -89.240 -173.640 -89.130 ;
        RECT -173.300 -89.240 -173.140 -88.450 ;
        RECT -171.700 -88.600 -171.360 -88.450 ;
        RECT -169.000 -88.450 -167.060 -88.300 ;
        RECT -169.000 -88.600 -168.660 -88.450 ;
        RECT -171.680 -88.800 -171.360 -88.770 ;
        RECT -173.960 -89.380 -173.140 -89.240 ;
        RECT -172.180 -88.940 -171.360 -88.800 ;
        RECT -173.960 -89.410 -173.640 -89.380 ;
        RECT -176.660 -89.730 -176.320 -89.580 ;
        RECT -178.260 -89.880 -176.320 -89.730 ;
        RECT -173.960 -89.730 -173.620 -89.580 ;
        RECT -172.180 -89.730 -172.020 -88.940 ;
        RECT -171.680 -89.050 -171.360 -88.940 ;
        RECT -169.000 -88.800 -168.680 -88.770 ;
        RECT -169.000 -88.940 -168.180 -88.800 ;
        RECT -169.000 -89.050 -168.680 -88.940 ;
        RECT -173.960 -89.880 -172.020 -89.730 ;
        RECT -168.340 -89.730 -168.180 -88.940 ;
        RECT -167.220 -89.240 -167.060 -88.450 ;
        RECT -163.380 -88.450 -161.440 -88.300 ;
        RECT -166.720 -89.240 -166.400 -89.130 ;
        RECT -167.220 -89.380 -166.400 -89.240 ;
        RECT -166.720 -89.410 -166.400 -89.380 ;
        RECT -164.040 -89.240 -163.720 -89.130 ;
        RECT -163.380 -89.240 -163.220 -88.450 ;
        RECT -161.780 -88.600 -161.440 -88.450 ;
        RECT -159.080 -88.450 -157.140 -88.300 ;
        RECT -159.080 -88.600 -158.740 -88.450 ;
        RECT -161.760 -88.800 -161.440 -88.770 ;
        RECT -164.040 -89.380 -163.220 -89.240 ;
        RECT -162.260 -88.940 -161.440 -88.800 ;
        RECT -164.040 -89.410 -163.720 -89.380 ;
        RECT -166.740 -89.730 -166.400 -89.580 ;
        RECT -168.340 -89.880 -166.400 -89.730 ;
        RECT -164.040 -89.730 -163.700 -89.580 ;
        RECT -162.260 -89.730 -162.100 -88.940 ;
        RECT -161.760 -89.050 -161.440 -88.940 ;
        RECT -159.080 -88.800 -158.760 -88.770 ;
        RECT -159.080 -88.940 -158.260 -88.800 ;
        RECT -159.080 -89.050 -158.760 -88.940 ;
        RECT -164.040 -89.880 -162.100 -89.730 ;
        RECT -158.420 -89.730 -158.260 -88.940 ;
        RECT -157.300 -89.240 -157.140 -88.450 ;
        RECT -153.460 -88.450 -151.520 -88.300 ;
        RECT -156.800 -89.240 -156.480 -89.130 ;
        RECT -157.300 -89.380 -156.480 -89.240 ;
        RECT -156.800 -89.410 -156.480 -89.380 ;
        RECT -154.120 -89.240 -153.800 -89.130 ;
        RECT -153.460 -89.240 -153.300 -88.450 ;
        RECT -151.860 -88.600 -151.520 -88.450 ;
        RECT -149.160 -88.450 -147.220 -88.300 ;
        RECT -149.160 -88.600 -148.820 -88.450 ;
        RECT -151.840 -88.800 -151.520 -88.770 ;
        RECT -154.120 -89.380 -153.300 -89.240 ;
        RECT -152.340 -88.940 -151.520 -88.800 ;
        RECT -154.120 -89.410 -153.800 -89.380 ;
        RECT -156.820 -89.730 -156.480 -89.580 ;
        RECT -158.420 -89.880 -156.480 -89.730 ;
        RECT -154.120 -89.730 -153.780 -89.580 ;
        RECT -152.340 -89.730 -152.180 -88.940 ;
        RECT -151.840 -89.050 -151.520 -88.940 ;
        RECT -149.160 -88.800 -148.840 -88.770 ;
        RECT -149.160 -88.940 -148.340 -88.800 ;
        RECT -149.160 -89.050 -148.840 -88.940 ;
        RECT -154.120 -89.880 -152.180 -89.730 ;
        RECT -148.500 -89.730 -148.340 -88.940 ;
        RECT -147.380 -89.240 -147.220 -88.450 ;
        RECT -143.540 -88.450 -141.600 -88.300 ;
        RECT -146.880 -89.240 -146.560 -89.130 ;
        RECT -147.380 -89.380 -146.560 -89.240 ;
        RECT -146.880 -89.410 -146.560 -89.380 ;
        RECT -144.200 -89.240 -143.880 -89.130 ;
        RECT -143.540 -89.240 -143.380 -88.450 ;
        RECT -141.940 -88.600 -141.600 -88.450 ;
        RECT -139.240 -88.450 -137.300 -88.300 ;
        RECT -139.240 -88.600 -138.900 -88.450 ;
        RECT -141.920 -88.800 -141.600 -88.770 ;
        RECT -144.200 -89.380 -143.380 -89.240 ;
        RECT -142.420 -88.940 -141.600 -88.800 ;
        RECT -144.200 -89.410 -143.880 -89.380 ;
        RECT -146.900 -89.730 -146.560 -89.580 ;
        RECT -148.500 -89.880 -146.560 -89.730 ;
        RECT -144.200 -89.730 -143.860 -89.580 ;
        RECT -142.420 -89.730 -142.260 -88.940 ;
        RECT -141.920 -89.050 -141.600 -88.940 ;
        RECT -139.240 -88.800 -138.920 -88.770 ;
        RECT -139.240 -88.940 -138.420 -88.800 ;
        RECT -139.240 -89.050 -138.920 -88.940 ;
        RECT -144.200 -89.880 -142.260 -89.730 ;
        RECT -138.580 -89.730 -138.420 -88.940 ;
        RECT -137.460 -89.240 -137.300 -88.450 ;
        RECT -133.620 -88.450 -131.680 -88.300 ;
        RECT -136.960 -89.240 -136.640 -89.130 ;
        RECT -137.460 -89.380 -136.640 -89.240 ;
        RECT -136.960 -89.410 -136.640 -89.380 ;
        RECT -134.280 -89.240 -133.960 -89.130 ;
        RECT -133.620 -89.240 -133.460 -88.450 ;
        RECT -132.020 -88.600 -131.680 -88.450 ;
        RECT -129.320 -88.450 -127.380 -88.300 ;
        RECT -129.320 -88.600 -128.980 -88.450 ;
        RECT -132.000 -88.800 -131.680 -88.770 ;
        RECT -134.280 -89.380 -133.460 -89.240 ;
        RECT -132.500 -88.940 -131.680 -88.800 ;
        RECT -134.280 -89.410 -133.960 -89.380 ;
        RECT -136.980 -89.730 -136.640 -89.580 ;
        RECT -138.580 -89.880 -136.640 -89.730 ;
        RECT -134.280 -89.730 -133.940 -89.580 ;
        RECT -132.500 -89.730 -132.340 -88.940 ;
        RECT -132.000 -89.050 -131.680 -88.940 ;
        RECT -129.320 -88.800 -129.000 -88.770 ;
        RECT -129.320 -88.940 -128.500 -88.800 ;
        RECT -129.320 -89.050 -129.000 -88.940 ;
        RECT -134.280 -89.880 -132.340 -89.730 ;
        RECT -128.660 -89.730 -128.500 -88.940 ;
        RECT -127.540 -89.240 -127.380 -88.450 ;
        RECT -123.700 -88.450 -121.760 -88.300 ;
        RECT -127.040 -89.240 -126.720 -89.130 ;
        RECT -127.540 -89.380 -126.720 -89.240 ;
        RECT -127.040 -89.410 -126.720 -89.380 ;
        RECT -124.360 -89.240 -124.040 -89.130 ;
        RECT -123.700 -89.240 -123.540 -88.450 ;
        RECT -122.100 -88.600 -121.760 -88.450 ;
        RECT -119.400 -88.450 -117.460 -88.300 ;
        RECT -119.400 -88.600 -119.060 -88.450 ;
        RECT -122.080 -88.800 -121.760 -88.770 ;
        RECT -124.360 -89.380 -123.540 -89.240 ;
        RECT -122.580 -88.940 -121.760 -88.800 ;
        RECT -124.360 -89.410 -124.040 -89.380 ;
        RECT -127.060 -89.730 -126.720 -89.580 ;
        RECT -128.660 -89.880 -126.720 -89.730 ;
        RECT -124.360 -89.730 -124.020 -89.580 ;
        RECT -122.580 -89.730 -122.420 -88.940 ;
        RECT -122.080 -89.050 -121.760 -88.940 ;
        RECT -119.400 -88.800 -119.080 -88.770 ;
        RECT -119.400 -88.940 -118.580 -88.800 ;
        RECT -119.400 -89.050 -119.080 -88.940 ;
        RECT -124.360 -89.880 -122.420 -89.730 ;
        RECT -118.740 -89.730 -118.580 -88.940 ;
        RECT -117.620 -89.240 -117.460 -88.450 ;
        RECT -113.780 -88.450 -111.840 -88.300 ;
        RECT -117.120 -89.240 -116.800 -89.130 ;
        RECT -117.620 -89.380 -116.800 -89.240 ;
        RECT -117.120 -89.410 -116.800 -89.380 ;
        RECT -114.440 -89.240 -114.120 -89.130 ;
        RECT -113.780 -89.240 -113.620 -88.450 ;
        RECT -112.180 -88.600 -111.840 -88.450 ;
        RECT -109.480 -88.450 -107.540 -88.300 ;
        RECT -109.480 -88.600 -109.140 -88.450 ;
        RECT -112.160 -88.800 -111.840 -88.770 ;
        RECT -114.440 -89.380 -113.620 -89.240 ;
        RECT -112.660 -88.940 -111.840 -88.800 ;
        RECT -114.440 -89.410 -114.120 -89.380 ;
        RECT -117.140 -89.730 -116.800 -89.580 ;
        RECT -118.740 -89.880 -116.800 -89.730 ;
        RECT -114.440 -89.730 -114.100 -89.580 ;
        RECT -112.660 -89.730 -112.500 -88.940 ;
        RECT -112.160 -89.050 -111.840 -88.940 ;
        RECT -109.480 -88.800 -109.160 -88.770 ;
        RECT -109.480 -88.940 -108.660 -88.800 ;
        RECT -109.480 -89.050 -109.160 -88.940 ;
        RECT -114.440 -89.880 -112.500 -89.730 ;
        RECT -108.820 -89.730 -108.660 -88.940 ;
        RECT -107.700 -89.240 -107.540 -88.450 ;
        RECT -103.860 -88.450 -101.920 -88.300 ;
        RECT -107.200 -89.240 -106.880 -89.130 ;
        RECT -107.700 -89.380 -106.880 -89.240 ;
        RECT -107.200 -89.410 -106.880 -89.380 ;
        RECT -104.520 -89.240 -104.200 -89.130 ;
        RECT -103.860 -89.240 -103.700 -88.450 ;
        RECT -102.260 -88.600 -101.920 -88.450 ;
        RECT -99.560 -88.450 -97.620 -88.300 ;
        RECT -99.560 -88.600 -99.220 -88.450 ;
        RECT -102.240 -88.800 -101.920 -88.770 ;
        RECT -104.520 -89.380 -103.700 -89.240 ;
        RECT -102.740 -88.940 -101.920 -88.800 ;
        RECT -104.520 -89.410 -104.200 -89.380 ;
        RECT -107.220 -89.730 -106.880 -89.580 ;
        RECT -108.820 -89.880 -106.880 -89.730 ;
        RECT -104.520 -89.730 -104.180 -89.580 ;
        RECT -102.740 -89.730 -102.580 -88.940 ;
        RECT -102.240 -89.050 -101.920 -88.940 ;
        RECT -99.560 -88.800 -99.240 -88.770 ;
        RECT -99.560 -88.940 -98.740 -88.800 ;
        RECT -99.560 -89.050 -99.240 -88.940 ;
        RECT -104.520 -89.880 -102.580 -89.730 ;
        RECT -98.900 -89.730 -98.740 -88.940 ;
        RECT -97.780 -89.240 -97.620 -88.450 ;
        RECT -93.940 -88.450 -92.000 -88.300 ;
        RECT -97.280 -89.240 -96.960 -89.130 ;
        RECT -97.780 -89.380 -96.960 -89.240 ;
        RECT -97.280 -89.410 -96.960 -89.380 ;
        RECT -94.600 -89.240 -94.280 -89.130 ;
        RECT -93.940 -89.240 -93.780 -88.450 ;
        RECT -92.340 -88.600 -92.000 -88.450 ;
        RECT -89.640 -88.450 -87.700 -88.300 ;
        RECT -89.640 -88.600 -89.300 -88.450 ;
        RECT -92.320 -88.800 -92.000 -88.770 ;
        RECT -94.600 -89.380 -93.780 -89.240 ;
        RECT -92.820 -88.940 -92.000 -88.800 ;
        RECT -94.600 -89.410 -94.280 -89.380 ;
        RECT -97.300 -89.730 -96.960 -89.580 ;
        RECT -98.900 -89.880 -96.960 -89.730 ;
        RECT -94.600 -89.730 -94.260 -89.580 ;
        RECT -92.820 -89.730 -92.660 -88.940 ;
        RECT -92.320 -89.050 -92.000 -88.940 ;
        RECT -89.640 -88.800 -89.320 -88.770 ;
        RECT -89.640 -88.940 -88.820 -88.800 ;
        RECT -89.640 -89.050 -89.320 -88.940 ;
        RECT -94.600 -89.880 -92.660 -89.730 ;
        RECT -88.980 -89.730 -88.820 -88.940 ;
        RECT -87.860 -89.240 -87.700 -88.450 ;
        RECT -84.020 -88.450 -82.080 -88.300 ;
        RECT -87.360 -89.240 -87.040 -89.130 ;
        RECT -87.860 -89.380 -87.040 -89.240 ;
        RECT -87.360 -89.410 -87.040 -89.380 ;
        RECT -84.680 -89.240 -84.360 -89.130 ;
        RECT -84.020 -89.240 -83.860 -88.450 ;
        RECT -82.420 -88.600 -82.080 -88.450 ;
        RECT -79.720 -88.450 -77.780 -88.300 ;
        RECT -79.720 -88.600 -79.380 -88.450 ;
        RECT -82.400 -88.800 -82.080 -88.770 ;
        RECT -84.680 -89.380 -83.860 -89.240 ;
        RECT -82.900 -88.940 -82.080 -88.800 ;
        RECT -84.680 -89.410 -84.360 -89.380 ;
        RECT -87.380 -89.730 -87.040 -89.580 ;
        RECT -88.980 -89.880 -87.040 -89.730 ;
        RECT -84.680 -89.730 -84.340 -89.580 ;
        RECT -82.900 -89.730 -82.740 -88.940 ;
        RECT -82.400 -89.050 -82.080 -88.940 ;
        RECT -79.720 -88.800 -79.400 -88.770 ;
        RECT -79.720 -88.940 -78.900 -88.800 ;
        RECT -79.720 -89.050 -79.400 -88.940 ;
        RECT -84.680 -89.880 -82.740 -89.730 ;
        RECT -79.060 -89.730 -78.900 -88.940 ;
        RECT -77.940 -89.240 -77.780 -88.450 ;
        RECT -74.100 -88.450 -72.160 -88.300 ;
        RECT -77.440 -89.240 -77.120 -89.130 ;
        RECT -77.940 -89.380 -77.120 -89.240 ;
        RECT -77.440 -89.410 -77.120 -89.380 ;
        RECT -74.760 -89.240 -74.440 -89.130 ;
        RECT -74.100 -89.240 -73.940 -88.450 ;
        RECT -72.500 -88.600 -72.160 -88.450 ;
        RECT -69.800 -88.450 -67.860 -88.300 ;
        RECT -69.800 -88.600 -69.460 -88.450 ;
        RECT -72.480 -88.800 -72.160 -88.770 ;
        RECT -74.760 -89.380 -73.940 -89.240 ;
        RECT -72.980 -88.940 -72.160 -88.800 ;
        RECT -74.760 -89.410 -74.440 -89.380 ;
        RECT -77.460 -89.730 -77.120 -89.580 ;
        RECT -79.060 -89.880 -77.120 -89.730 ;
        RECT -74.760 -89.730 -74.420 -89.580 ;
        RECT -72.980 -89.730 -72.820 -88.940 ;
        RECT -72.480 -89.050 -72.160 -88.940 ;
        RECT -69.800 -88.800 -69.480 -88.770 ;
        RECT -69.800 -88.940 -68.980 -88.800 ;
        RECT -69.800 -89.050 -69.480 -88.940 ;
        RECT -74.760 -89.880 -72.820 -89.730 ;
        RECT -69.140 -89.730 -68.980 -88.940 ;
        RECT -68.020 -89.240 -67.860 -88.450 ;
        RECT -64.180 -88.450 -62.240 -88.300 ;
        RECT -67.520 -89.240 -67.200 -89.130 ;
        RECT -68.020 -89.380 -67.200 -89.240 ;
        RECT -67.520 -89.410 -67.200 -89.380 ;
        RECT -64.840 -89.240 -64.520 -89.130 ;
        RECT -64.180 -89.240 -64.020 -88.450 ;
        RECT -62.580 -88.600 -62.240 -88.450 ;
        RECT -59.880 -88.450 -57.940 -88.300 ;
        RECT -59.880 -88.600 -59.540 -88.450 ;
        RECT -62.560 -88.800 -62.240 -88.770 ;
        RECT -64.840 -89.380 -64.020 -89.240 ;
        RECT -63.060 -88.940 -62.240 -88.800 ;
        RECT -64.840 -89.410 -64.520 -89.380 ;
        RECT -67.540 -89.730 -67.200 -89.580 ;
        RECT -69.140 -89.880 -67.200 -89.730 ;
        RECT -64.840 -89.730 -64.500 -89.580 ;
        RECT -63.060 -89.730 -62.900 -88.940 ;
        RECT -62.560 -89.050 -62.240 -88.940 ;
        RECT -59.880 -88.800 -59.560 -88.770 ;
        RECT -59.880 -88.940 -59.060 -88.800 ;
        RECT -59.880 -89.050 -59.560 -88.940 ;
        RECT -64.840 -89.880 -62.900 -89.730 ;
        RECT -59.220 -89.730 -59.060 -88.940 ;
        RECT -58.100 -89.240 -57.940 -88.450 ;
        RECT -54.260 -88.450 -52.320 -88.300 ;
        RECT -57.600 -89.240 -57.280 -89.130 ;
        RECT -58.100 -89.380 -57.280 -89.240 ;
        RECT -57.600 -89.410 -57.280 -89.380 ;
        RECT -54.920 -89.240 -54.600 -89.130 ;
        RECT -54.260 -89.240 -54.100 -88.450 ;
        RECT -52.660 -88.600 -52.320 -88.450 ;
        RECT -49.960 -88.450 -48.020 -88.300 ;
        RECT -49.960 -88.600 -49.620 -88.450 ;
        RECT -52.640 -88.800 -52.320 -88.770 ;
        RECT -54.920 -89.380 -54.100 -89.240 ;
        RECT -53.140 -88.940 -52.320 -88.800 ;
        RECT -54.920 -89.410 -54.600 -89.380 ;
        RECT -57.620 -89.730 -57.280 -89.580 ;
        RECT -59.220 -89.880 -57.280 -89.730 ;
        RECT -54.920 -89.730 -54.580 -89.580 ;
        RECT -53.140 -89.730 -52.980 -88.940 ;
        RECT -52.640 -89.050 -52.320 -88.940 ;
        RECT -49.960 -88.800 -49.640 -88.770 ;
        RECT -49.960 -88.940 -49.140 -88.800 ;
        RECT -49.960 -89.050 -49.640 -88.940 ;
        RECT -54.920 -89.880 -52.980 -89.730 ;
        RECT -49.300 -89.730 -49.140 -88.940 ;
        RECT -48.180 -89.240 -48.020 -88.450 ;
        RECT -44.340 -88.450 -42.400 -88.300 ;
        RECT -47.680 -89.240 -47.360 -89.130 ;
        RECT -48.180 -89.380 -47.360 -89.240 ;
        RECT -47.680 -89.410 -47.360 -89.380 ;
        RECT -45.000 -89.240 -44.680 -89.130 ;
        RECT -44.340 -89.240 -44.180 -88.450 ;
        RECT -42.740 -88.600 -42.400 -88.450 ;
        RECT -40.040 -88.450 -38.100 -88.300 ;
        RECT -40.040 -88.600 -39.700 -88.450 ;
        RECT -42.720 -88.800 -42.400 -88.770 ;
        RECT -45.000 -89.380 -44.180 -89.240 ;
        RECT -43.220 -88.940 -42.400 -88.800 ;
        RECT -45.000 -89.410 -44.680 -89.380 ;
        RECT -47.700 -89.730 -47.360 -89.580 ;
        RECT -49.300 -89.880 -47.360 -89.730 ;
        RECT -45.000 -89.730 -44.660 -89.580 ;
        RECT -43.220 -89.730 -43.060 -88.940 ;
        RECT -42.720 -89.050 -42.400 -88.940 ;
        RECT -40.040 -88.800 -39.720 -88.770 ;
        RECT -40.040 -88.940 -39.220 -88.800 ;
        RECT -40.040 -89.050 -39.720 -88.940 ;
        RECT -45.000 -89.880 -43.060 -89.730 ;
        RECT -39.380 -89.730 -39.220 -88.940 ;
        RECT -38.260 -89.240 -38.100 -88.450 ;
        RECT -34.420 -88.450 -32.480 -88.300 ;
        RECT -37.760 -89.240 -37.440 -89.130 ;
        RECT -38.260 -89.380 -37.440 -89.240 ;
        RECT -37.760 -89.410 -37.440 -89.380 ;
        RECT -35.080 -89.240 -34.760 -89.130 ;
        RECT -34.420 -89.240 -34.260 -88.450 ;
        RECT -32.820 -88.600 -32.480 -88.450 ;
        RECT -30.120 -88.450 -28.180 -88.300 ;
        RECT -30.120 -88.600 -29.780 -88.450 ;
        RECT -32.800 -88.800 -32.480 -88.770 ;
        RECT -35.080 -89.380 -34.260 -89.240 ;
        RECT -33.300 -88.940 -32.480 -88.800 ;
        RECT -35.080 -89.410 -34.760 -89.380 ;
        RECT -37.780 -89.730 -37.440 -89.580 ;
        RECT -39.380 -89.880 -37.440 -89.730 ;
        RECT -35.080 -89.730 -34.740 -89.580 ;
        RECT -33.300 -89.730 -33.140 -88.940 ;
        RECT -32.800 -89.050 -32.480 -88.940 ;
        RECT -30.120 -88.800 -29.800 -88.770 ;
        RECT -30.120 -88.940 -29.300 -88.800 ;
        RECT -30.120 -89.050 -29.800 -88.940 ;
        RECT -35.080 -89.880 -33.140 -89.730 ;
        RECT -29.460 -89.730 -29.300 -88.940 ;
        RECT -28.340 -89.240 -28.180 -88.450 ;
        RECT -24.500 -88.450 -22.560 -88.300 ;
        RECT -27.840 -89.240 -27.520 -89.130 ;
        RECT -28.340 -89.380 -27.520 -89.240 ;
        RECT -27.840 -89.410 -27.520 -89.380 ;
        RECT -25.160 -89.240 -24.840 -89.130 ;
        RECT -24.500 -89.240 -24.340 -88.450 ;
        RECT -22.900 -88.600 -22.560 -88.450 ;
        RECT -20.200 -88.450 -18.260 -88.300 ;
        RECT -20.200 -88.600 -19.860 -88.450 ;
        RECT -22.880 -88.800 -22.560 -88.770 ;
        RECT -25.160 -89.380 -24.340 -89.240 ;
        RECT -23.380 -88.940 -22.560 -88.800 ;
        RECT -25.160 -89.410 -24.840 -89.380 ;
        RECT -27.860 -89.730 -27.520 -89.580 ;
        RECT -29.460 -89.880 -27.520 -89.730 ;
        RECT -25.160 -89.730 -24.820 -89.580 ;
        RECT -23.380 -89.730 -23.220 -88.940 ;
        RECT -22.880 -89.050 -22.560 -88.940 ;
        RECT -20.200 -88.800 -19.880 -88.770 ;
        RECT -20.200 -88.940 -19.380 -88.800 ;
        RECT -20.200 -89.050 -19.880 -88.940 ;
        RECT -25.160 -89.880 -23.220 -89.730 ;
        RECT -19.540 -89.730 -19.380 -88.940 ;
        RECT -18.420 -89.240 -18.260 -88.450 ;
        RECT -14.580 -88.450 -12.640 -88.300 ;
        RECT -17.920 -89.240 -17.600 -89.130 ;
        RECT -18.420 -89.380 -17.600 -89.240 ;
        RECT -17.920 -89.410 -17.600 -89.380 ;
        RECT -15.240 -89.240 -14.920 -89.130 ;
        RECT -14.580 -89.240 -14.420 -88.450 ;
        RECT -12.980 -88.600 -12.640 -88.450 ;
        RECT -10.280 -88.450 -8.340 -88.300 ;
        RECT -10.280 -88.600 -9.940 -88.450 ;
        RECT -12.960 -88.800 -12.640 -88.770 ;
        RECT -15.240 -89.380 -14.420 -89.240 ;
        RECT -13.460 -88.940 -12.640 -88.800 ;
        RECT -15.240 -89.410 -14.920 -89.380 ;
        RECT -17.940 -89.730 -17.600 -89.580 ;
        RECT -19.540 -89.880 -17.600 -89.730 ;
        RECT -15.240 -89.730 -14.900 -89.580 ;
        RECT -13.460 -89.730 -13.300 -88.940 ;
        RECT -12.960 -89.050 -12.640 -88.940 ;
        RECT -10.280 -88.800 -9.960 -88.770 ;
        RECT -10.280 -88.940 -9.460 -88.800 ;
        RECT -10.280 -89.050 -9.960 -88.940 ;
        RECT -15.240 -89.880 -13.300 -89.730 ;
        RECT -9.620 -89.730 -9.460 -88.940 ;
        RECT -8.500 -89.240 -8.340 -88.450 ;
        RECT -4.660 -88.450 -2.720 -88.300 ;
        RECT -8.000 -89.240 -7.680 -89.130 ;
        RECT -8.500 -89.380 -7.680 -89.240 ;
        RECT -8.000 -89.410 -7.680 -89.380 ;
        RECT -5.320 -89.240 -5.000 -89.130 ;
        RECT -4.660 -89.240 -4.500 -88.450 ;
        RECT -3.060 -88.600 -2.720 -88.450 ;
        RECT -0.360 -88.450 1.580 -88.300 ;
        RECT -0.360 -88.600 -0.020 -88.450 ;
        RECT -3.040 -88.800 -2.720 -88.770 ;
        RECT -5.320 -89.380 -4.500 -89.240 ;
        RECT -3.540 -88.940 -2.720 -88.800 ;
        RECT -5.320 -89.410 -5.000 -89.380 ;
        RECT -8.020 -89.730 -7.680 -89.580 ;
        RECT -9.620 -89.880 -7.680 -89.730 ;
        RECT -5.320 -89.730 -4.980 -89.580 ;
        RECT -3.540 -89.730 -3.380 -88.940 ;
        RECT -3.040 -89.050 -2.720 -88.940 ;
        RECT -0.360 -88.800 -0.040 -88.770 ;
        RECT -0.360 -88.940 0.460 -88.800 ;
        RECT -0.360 -89.050 -0.040 -88.940 ;
        RECT -5.320 -89.880 -3.380 -89.730 ;
        RECT 0.300 -89.730 0.460 -88.940 ;
        RECT 1.420 -89.240 1.580 -88.450 ;
        RECT 5.260 -88.450 7.200 -88.300 ;
        RECT 1.920 -89.240 2.240 -89.130 ;
        RECT 1.420 -89.380 2.240 -89.240 ;
        RECT 1.920 -89.410 2.240 -89.380 ;
        RECT 4.600 -89.240 4.920 -89.130 ;
        RECT 5.260 -89.240 5.420 -88.450 ;
        RECT 6.860 -88.600 7.200 -88.450 ;
        RECT 9.560 -88.450 11.500 -88.300 ;
        RECT 9.560 -88.600 9.900 -88.450 ;
        RECT 6.880 -88.800 7.200 -88.770 ;
        RECT 4.600 -89.380 5.420 -89.240 ;
        RECT 6.380 -88.940 7.200 -88.800 ;
        RECT 4.600 -89.410 4.920 -89.380 ;
        RECT 1.900 -89.730 2.240 -89.580 ;
        RECT 0.300 -89.880 2.240 -89.730 ;
        RECT 4.600 -89.730 4.940 -89.580 ;
        RECT 6.380 -89.730 6.540 -88.940 ;
        RECT 6.880 -89.050 7.200 -88.940 ;
        RECT 9.560 -88.800 9.880 -88.770 ;
        RECT 9.560 -88.940 10.380 -88.800 ;
        RECT 9.560 -89.050 9.880 -88.940 ;
        RECT 4.600 -89.880 6.540 -89.730 ;
        RECT 10.220 -89.730 10.380 -88.940 ;
        RECT 11.340 -89.240 11.500 -88.450 ;
        RECT 15.180 -88.450 17.120 -88.300 ;
        RECT 11.840 -89.240 12.160 -89.130 ;
        RECT 11.340 -89.380 12.160 -89.240 ;
        RECT 11.840 -89.410 12.160 -89.380 ;
        RECT 14.520 -89.240 14.840 -89.130 ;
        RECT 15.180 -89.240 15.340 -88.450 ;
        RECT 16.780 -88.600 17.120 -88.450 ;
        RECT 19.480 -88.450 21.420 -88.300 ;
        RECT 19.480 -88.600 19.820 -88.450 ;
        RECT 16.800 -88.800 17.120 -88.770 ;
        RECT 14.520 -89.380 15.340 -89.240 ;
        RECT 16.300 -88.940 17.120 -88.800 ;
        RECT 14.520 -89.410 14.840 -89.380 ;
        RECT 11.820 -89.730 12.160 -89.580 ;
        RECT 10.220 -89.880 12.160 -89.730 ;
        RECT 14.520 -89.730 14.860 -89.580 ;
        RECT 16.300 -89.730 16.460 -88.940 ;
        RECT 16.800 -89.050 17.120 -88.940 ;
        RECT 19.480 -88.800 19.800 -88.770 ;
        RECT 19.480 -88.940 20.300 -88.800 ;
        RECT 19.480 -89.050 19.800 -88.940 ;
        RECT 14.520 -89.880 16.460 -89.730 ;
        RECT 20.140 -89.730 20.300 -88.940 ;
        RECT 21.260 -89.240 21.420 -88.450 ;
        RECT 25.100 -88.450 27.040 -88.300 ;
        RECT 21.760 -89.240 22.080 -89.130 ;
        RECT 21.260 -89.380 22.080 -89.240 ;
        RECT 21.760 -89.410 22.080 -89.380 ;
        RECT 24.440 -89.240 24.760 -89.130 ;
        RECT 25.100 -89.240 25.260 -88.450 ;
        RECT 26.700 -88.600 27.040 -88.450 ;
        RECT 26.720 -88.800 27.040 -88.770 ;
        RECT 24.440 -89.380 25.260 -89.240 ;
        RECT 26.220 -88.940 27.040 -88.800 ;
        RECT 24.440 -89.410 24.760 -89.380 ;
        RECT 21.740 -89.730 22.080 -89.580 ;
        RECT 20.140 -89.880 22.080 -89.730 ;
        RECT 24.440 -89.730 24.780 -89.580 ;
        RECT 26.220 -89.730 26.380 -88.940 ;
        RECT 26.720 -89.050 27.040 -88.940 ;
        RECT 24.440 -89.880 26.380 -89.730 ;
        RECT -289.450 -90.690 -287.610 -90.210 ;
        RECT -287.690 -91.780 -287.210 -90.880 ;
        RECT -286.390 -91.010 -286.200 -89.880 ;
        RECT -282.320 -91.010 -282.130 -89.880 ;
        RECT -276.470 -91.010 -276.280 -89.880 ;
        RECT -272.400 -91.010 -272.210 -89.880 ;
        RECT -266.550 -91.010 -266.360 -89.880 ;
        RECT -262.480 -91.010 -262.290 -89.880 ;
        RECT -256.630 -91.010 -256.440 -89.880 ;
        RECT -252.560 -91.010 -252.370 -89.880 ;
        RECT -246.710 -91.010 -246.520 -89.880 ;
        RECT -242.640 -91.010 -242.450 -89.880 ;
        RECT -236.790 -91.010 -236.600 -89.880 ;
        RECT -232.720 -91.010 -232.530 -89.880 ;
        RECT -226.870 -91.010 -226.680 -89.880 ;
        RECT -222.800 -91.010 -222.610 -89.880 ;
        RECT -216.950 -91.010 -216.760 -89.880 ;
        RECT -212.880 -91.010 -212.690 -89.880 ;
        RECT -207.030 -91.010 -206.840 -89.880 ;
        RECT -202.960 -91.010 -202.770 -89.880 ;
        RECT -197.110 -91.010 -196.920 -89.880 ;
        RECT -193.040 -91.010 -192.850 -89.880 ;
        RECT -187.190 -91.010 -187.000 -89.880 ;
        RECT -183.120 -91.010 -182.930 -89.880 ;
        RECT -177.270 -91.010 -177.080 -89.880 ;
        RECT -173.200 -91.010 -173.010 -89.880 ;
        RECT -167.350 -91.010 -167.160 -89.880 ;
        RECT -163.280 -91.010 -163.090 -89.880 ;
        RECT -157.430 -91.010 -157.240 -89.880 ;
        RECT -153.360 -91.010 -153.170 -89.880 ;
        RECT -147.510 -91.010 -147.320 -89.880 ;
        RECT -143.440 -91.010 -143.250 -89.880 ;
        RECT -137.590 -91.010 -137.400 -89.880 ;
        RECT -133.520 -91.010 -133.330 -89.880 ;
        RECT -127.670 -91.010 -127.480 -89.880 ;
        RECT -123.600 -91.010 -123.410 -89.880 ;
        RECT -117.750 -91.010 -117.560 -89.880 ;
        RECT -113.680 -91.010 -113.490 -89.880 ;
        RECT -107.830 -91.010 -107.640 -89.880 ;
        RECT -103.760 -91.010 -103.570 -89.880 ;
        RECT -97.910 -91.010 -97.720 -89.880 ;
        RECT -93.840 -91.010 -93.650 -89.880 ;
        RECT -87.990 -91.010 -87.800 -89.880 ;
        RECT -83.920 -91.010 -83.730 -89.880 ;
        RECT -78.070 -91.010 -77.880 -89.880 ;
        RECT -74.000 -91.010 -73.810 -89.880 ;
        RECT -68.150 -91.010 -67.960 -89.880 ;
        RECT -64.080 -91.010 -63.890 -89.880 ;
        RECT -58.230 -91.010 -58.040 -89.880 ;
        RECT -54.160 -91.010 -53.970 -89.880 ;
        RECT -48.310 -91.010 -48.120 -89.880 ;
        RECT -44.240 -91.010 -44.050 -89.880 ;
        RECT -38.390 -91.010 -38.200 -89.880 ;
        RECT -34.320 -91.010 -34.130 -89.880 ;
        RECT -28.470 -91.010 -28.280 -89.880 ;
        RECT -24.400 -91.010 -24.210 -89.880 ;
        RECT -18.550 -91.010 -18.360 -89.880 ;
        RECT -14.480 -91.010 -14.290 -89.880 ;
        RECT -8.630 -91.010 -8.440 -89.880 ;
        RECT -4.560 -91.010 -4.370 -89.880 ;
        RECT 1.290 -91.010 1.480 -89.880 ;
        RECT 5.360 -91.010 5.550 -89.880 ;
        RECT 11.210 -91.010 11.400 -89.880 ;
        RECT 15.280 -91.010 15.470 -89.880 ;
        RECT 21.130 -91.010 21.320 -89.880 ;
        RECT 25.200 -91.010 25.390 -89.880 ;
        RECT -286.440 -91.300 -286.120 -91.010 ;
        RECT -282.400 -91.300 -282.080 -91.010 ;
        RECT -276.520 -91.300 -276.200 -91.010 ;
        RECT -272.480 -91.300 -272.160 -91.010 ;
        RECT -266.600 -91.300 -266.280 -91.010 ;
        RECT -262.560 -91.300 -262.240 -91.010 ;
        RECT -256.680 -91.300 -256.360 -91.010 ;
        RECT -252.640 -91.300 -252.320 -91.010 ;
        RECT -246.760 -91.300 -246.440 -91.010 ;
        RECT -242.720 -91.300 -242.400 -91.010 ;
        RECT -236.840 -91.300 -236.520 -91.010 ;
        RECT -232.800 -91.300 -232.480 -91.010 ;
        RECT -226.920 -91.300 -226.600 -91.010 ;
        RECT -222.880 -91.300 -222.560 -91.010 ;
        RECT -217.000 -91.300 -216.680 -91.010 ;
        RECT -212.960 -91.300 -212.640 -91.010 ;
        RECT -207.080 -91.300 -206.760 -91.010 ;
        RECT -203.040 -91.300 -202.720 -91.010 ;
        RECT -197.160 -91.300 -196.840 -91.010 ;
        RECT -193.120 -91.300 -192.800 -91.010 ;
        RECT -187.240 -91.300 -186.920 -91.010 ;
        RECT -183.200 -91.300 -182.880 -91.010 ;
        RECT -177.320 -91.300 -177.000 -91.010 ;
        RECT -173.280 -91.300 -172.960 -91.010 ;
        RECT -167.400 -91.300 -167.080 -91.010 ;
        RECT -163.360 -91.300 -163.040 -91.010 ;
        RECT -157.480 -91.300 -157.160 -91.010 ;
        RECT -153.440 -91.300 -153.120 -91.010 ;
        RECT -147.560 -91.300 -147.240 -91.010 ;
        RECT -143.520 -91.300 -143.200 -91.010 ;
        RECT -137.640 -91.300 -137.320 -91.010 ;
        RECT -133.600 -91.300 -133.280 -91.010 ;
        RECT -127.720 -91.300 -127.400 -91.010 ;
        RECT -123.680 -91.300 -123.360 -91.010 ;
        RECT -117.800 -91.300 -117.480 -91.010 ;
        RECT -113.760 -91.300 -113.440 -91.010 ;
        RECT -107.880 -91.300 -107.560 -91.010 ;
        RECT -103.840 -91.300 -103.520 -91.010 ;
        RECT -97.960 -91.300 -97.640 -91.010 ;
        RECT -93.920 -91.300 -93.600 -91.010 ;
        RECT -88.040 -91.300 -87.720 -91.010 ;
        RECT -84.000 -91.300 -83.680 -91.010 ;
        RECT -78.120 -91.300 -77.800 -91.010 ;
        RECT -74.080 -91.300 -73.760 -91.010 ;
        RECT -68.200 -91.300 -67.880 -91.010 ;
        RECT -64.160 -91.300 -63.840 -91.010 ;
        RECT -58.280 -91.300 -57.960 -91.010 ;
        RECT -54.240 -91.300 -53.920 -91.010 ;
        RECT -48.360 -91.300 -48.040 -91.010 ;
        RECT -44.320 -91.300 -44.000 -91.010 ;
        RECT -38.440 -91.300 -38.120 -91.010 ;
        RECT -34.400 -91.300 -34.080 -91.010 ;
        RECT -28.520 -91.300 -28.200 -91.010 ;
        RECT -24.480 -91.300 -24.160 -91.010 ;
        RECT -18.600 -91.300 -18.280 -91.010 ;
        RECT -14.560 -91.300 -14.240 -91.010 ;
        RECT -8.680 -91.300 -8.360 -91.010 ;
        RECT -4.640 -91.300 -4.320 -91.010 ;
        RECT 1.240 -91.300 1.560 -91.010 ;
        RECT 5.280 -91.300 5.600 -91.010 ;
        RECT 11.160 -91.300 11.480 -91.010 ;
        RECT 15.200 -91.300 15.520 -91.010 ;
        RECT 21.080 -91.300 21.400 -91.010 ;
        RECT 25.120 -91.300 25.440 -91.010 ;
        RECT -288.150 -92.260 -287.210 -91.780 ;
        RECT 26.210 -91.780 26.690 -90.880 ;
        RECT -283.140 -92.180 -281.450 -91.880 ;
        RECT -273.220 -92.180 -271.530 -91.880 ;
        RECT -263.300 -92.180 -261.610 -91.880 ;
        RECT -253.380 -92.180 -251.690 -91.880 ;
        RECT -243.460 -92.180 -241.770 -91.880 ;
        RECT -233.540 -92.180 -231.850 -91.880 ;
        RECT -223.620 -92.180 -221.930 -91.880 ;
        RECT -213.700 -92.180 -212.010 -91.880 ;
        RECT -203.780 -92.180 -202.090 -91.880 ;
        RECT -193.860 -92.180 -192.170 -91.880 ;
        RECT -183.940 -92.180 -182.250 -91.880 ;
        RECT -174.020 -92.180 -172.330 -91.880 ;
        RECT -164.100 -92.180 -162.410 -91.880 ;
        RECT -154.180 -92.180 -152.490 -91.880 ;
        RECT -144.260 -92.180 -142.570 -91.880 ;
        RECT -134.340 -92.180 -132.650 -91.880 ;
        RECT -124.420 -92.180 -122.730 -91.880 ;
        RECT -114.500 -92.180 -112.810 -91.880 ;
        RECT -104.580 -92.180 -102.890 -91.880 ;
        RECT -94.660 -92.180 -92.970 -91.880 ;
        RECT -84.740 -92.180 -83.050 -91.880 ;
        RECT -74.820 -92.180 -73.130 -91.880 ;
        RECT -64.900 -92.180 -63.210 -91.880 ;
        RECT -54.980 -92.180 -53.290 -91.880 ;
        RECT -45.060 -92.180 -43.370 -91.880 ;
        RECT -35.140 -92.180 -33.450 -91.880 ;
        RECT -25.220 -92.180 -23.530 -91.880 ;
        RECT -15.300 -92.180 -13.610 -91.880 ;
        RECT -5.380 -92.180 -3.690 -91.880 ;
        RECT 4.540 -92.180 6.230 -91.880 ;
        RECT 14.460 -92.180 16.150 -91.880 ;
        RECT 24.380 -92.180 26.070 -91.880 ;
        RECT -282.630 -92.880 -281.630 -92.180 ;
        RECT -272.710 -92.880 -271.710 -92.180 ;
        RECT -262.790 -92.880 -261.790 -92.180 ;
        RECT -252.870 -92.880 -251.870 -92.180 ;
        RECT -242.950 -92.880 -241.950 -92.180 ;
        RECT -233.030 -92.880 -232.030 -92.180 ;
        RECT -223.110 -92.880 -222.110 -92.180 ;
        RECT -213.190 -92.880 -212.190 -92.180 ;
        RECT -203.270 -92.880 -202.270 -92.180 ;
        RECT -193.350 -92.880 -192.350 -92.180 ;
        RECT -183.430 -92.880 -182.430 -92.180 ;
        RECT -173.510 -92.880 -172.510 -92.180 ;
        RECT -163.590 -92.880 -162.590 -92.180 ;
        RECT -153.670 -92.880 -152.670 -92.180 ;
        RECT -143.750 -92.880 -142.750 -92.180 ;
        RECT -133.830 -92.880 -132.830 -92.180 ;
        RECT -123.910 -92.880 -122.910 -92.180 ;
        RECT -113.990 -92.880 -112.990 -92.180 ;
        RECT -104.070 -92.880 -103.070 -92.180 ;
        RECT -94.150 -92.880 -93.150 -92.180 ;
        RECT -84.230 -92.880 -83.230 -92.180 ;
        RECT -74.310 -92.880 -73.310 -92.180 ;
        RECT -64.390 -92.880 -63.390 -92.180 ;
        RECT -54.470 -92.880 -53.470 -92.180 ;
        RECT -44.550 -92.880 -43.550 -92.180 ;
        RECT -34.630 -92.880 -33.630 -92.180 ;
        RECT -24.710 -92.880 -23.710 -92.180 ;
        RECT -14.790 -92.880 -13.790 -92.180 ;
        RECT -4.870 -92.880 -3.870 -92.180 ;
        RECT 5.050 -92.880 6.050 -92.180 ;
        RECT 14.970 -92.880 15.970 -92.180 ;
        RECT 24.890 -92.880 25.890 -92.180 ;
        RECT 26.210 -92.260 27.150 -91.780 ;
        RECT -289.200 -173.630 -288.740 -173.625 ;
        RECT -289.200 -174.105 -288.260 -173.630 ;
        RECT -287.340 -173.710 -286.340 -173.010 ;
        RECT -277.420 -173.710 -276.420 -173.010 ;
        RECT -267.500 -173.710 -266.500 -173.010 ;
        RECT -257.580 -173.710 -256.580 -173.010 ;
        RECT -247.660 -173.710 -246.660 -173.010 ;
        RECT -237.740 -173.710 -236.740 -173.010 ;
        RECT -227.820 -173.710 -226.820 -173.010 ;
        RECT -217.900 -173.710 -216.900 -173.010 ;
        RECT -207.980 -173.710 -206.980 -173.010 ;
        RECT -198.060 -173.710 -197.060 -173.010 ;
        RECT -188.140 -173.710 -187.140 -173.010 ;
        RECT -178.220 -173.710 -177.220 -173.010 ;
        RECT -168.300 -173.710 -167.300 -173.010 ;
        RECT -158.380 -173.710 -157.380 -173.010 ;
        RECT -148.460 -173.710 -147.460 -173.010 ;
        RECT -138.540 -173.710 -137.540 -173.010 ;
        RECT -128.620 -173.710 -127.620 -173.010 ;
        RECT -118.700 -173.710 -117.700 -173.010 ;
        RECT -108.780 -173.710 -107.780 -173.010 ;
        RECT -98.860 -173.710 -97.860 -173.010 ;
        RECT -88.940 -173.710 -87.940 -173.010 ;
        RECT -79.020 -173.710 -78.020 -173.010 ;
        RECT -69.100 -173.710 -68.100 -173.010 ;
        RECT -59.180 -173.710 -58.180 -173.010 ;
        RECT -49.260 -173.710 -48.260 -173.010 ;
        RECT -39.340 -173.710 -38.340 -173.010 ;
        RECT -29.420 -173.710 -28.420 -173.010 ;
        RECT -19.500 -173.710 -18.500 -173.010 ;
        RECT -9.580 -173.710 -8.580 -173.010 ;
        RECT 0.340 -173.710 1.340 -173.010 ;
        RECT 10.260 -173.710 11.260 -173.010 ;
        RECT 20.180 -173.710 21.180 -173.010 ;
        RECT -287.850 -174.010 -286.160 -173.710 ;
        RECT -277.930 -174.010 -276.240 -173.710 ;
        RECT -268.010 -174.010 -266.320 -173.710 ;
        RECT -258.090 -174.010 -256.400 -173.710 ;
        RECT -248.170 -174.010 -246.480 -173.710 ;
        RECT -238.250 -174.010 -236.560 -173.710 ;
        RECT -228.330 -174.010 -226.640 -173.710 ;
        RECT -218.410 -174.010 -216.720 -173.710 ;
        RECT -208.490 -174.010 -206.800 -173.710 ;
        RECT -198.570 -174.010 -196.880 -173.710 ;
        RECT -188.650 -174.010 -186.960 -173.710 ;
        RECT -178.730 -174.010 -177.040 -173.710 ;
        RECT -168.810 -174.010 -167.120 -173.710 ;
        RECT -158.890 -174.010 -157.200 -173.710 ;
        RECT -148.970 -174.010 -147.280 -173.710 ;
        RECT -139.050 -174.010 -137.360 -173.710 ;
        RECT -129.130 -174.010 -127.440 -173.710 ;
        RECT -119.210 -174.010 -117.520 -173.710 ;
        RECT -109.290 -174.010 -107.600 -173.710 ;
        RECT -99.370 -174.010 -97.680 -173.710 ;
        RECT -89.450 -174.010 -87.760 -173.710 ;
        RECT -79.530 -174.010 -77.840 -173.710 ;
        RECT -69.610 -174.010 -67.920 -173.710 ;
        RECT -59.690 -174.010 -58.000 -173.710 ;
        RECT -49.770 -174.010 -48.080 -173.710 ;
        RECT -39.850 -174.010 -38.160 -173.710 ;
        RECT -29.930 -174.010 -28.240 -173.710 ;
        RECT -20.010 -174.010 -18.320 -173.710 ;
        RECT -10.090 -174.010 -8.400 -173.710 ;
        RECT -0.170 -174.010 1.520 -173.710 ;
        RECT 9.750 -174.010 11.440 -173.710 ;
        RECT 19.670 -174.010 21.360 -173.710 ;
        RECT -288.740 -175.010 -288.260 -174.105 ;
        RECT -287.110 -174.880 -286.790 -174.590 ;
        RECT -281.230 -174.880 -280.910 -174.590 ;
        RECT -277.190 -174.880 -276.870 -174.590 ;
        RECT -271.310 -174.880 -270.990 -174.590 ;
        RECT -267.270 -174.880 -266.950 -174.590 ;
        RECT -261.390 -174.880 -261.070 -174.590 ;
        RECT -257.350 -174.880 -257.030 -174.590 ;
        RECT -251.470 -174.880 -251.150 -174.590 ;
        RECT -247.430 -174.880 -247.110 -174.590 ;
        RECT -241.550 -174.880 -241.230 -174.590 ;
        RECT -237.510 -174.880 -237.190 -174.590 ;
        RECT -231.630 -174.880 -231.310 -174.590 ;
        RECT -227.590 -174.880 -227.270 -174.590 ;
        RECT -221.710 -174.880 -221.390 -174.590 ;
        RECT -217.670 -174.880 -217.350 -174.590 ;
        RECT -211.790 -174.880 -211.470 -174.590 ;
        RECT -207.750 -174.880 -207.430 -174.590 ;
        RECT -201.870 -174.880 -201.550 -174.590 ;
        RECT -197.830 -174.880 -197.510 -174.590 ;
        RECT -191.950 -174.880 -191.630 -174.590 ;
        RECT -187.910 -174.880 -187.590 -174.590 ;
        RECT -182.030 -174.880 -181.710 -174.590 ;
        RECT -177.990 -174.880 -177.670 -174.590 ;
        RECT -172.110 -174.880 -171.790 -174.590 ;
        RECT -168.070 -174.880 -167.750 -174.590 ;
        RECT -162.190 -174.880 -161.870 -174.590 ;
        RECT -158.150 -174.880 -157.830 -174.590 ;
        RECT -152.270 -174.880 -151.950 -174.590 ;
        RECT -148.230 -174.880 -147.910 -174.590 ;
        RECT -142.350 -174.880 -142.030 -174.590 ;
        RECT -138.310 -174.880 -137.990 -174.590 ;
        RECT -132.430 -174.880 -132.110 -174.590 ;
        RECT -128.390 -174.880 -128.070 -174.590 ;
        RECT -122.510 -174.880 -122.190 -174.590 ;
        RECT -118.470 -174.880 -118.150 -174.590 ;
        RECT -112.590 -174.880 -112.270 -174.590 ;
        RECT -108.550 -174.880 -108.230 -174.590 ;
        RECT -102.670 -174.880 -102.350 -174.590 ;
        RECT -98.630 -174.880 -98.310 -174.590 ;
        RECT -92.750 -174.880 -92.430 -174.590 ;
        RECT -88.710 -174.880 -88.390 -174.590 ;
        RECT -82.830 -174.880 -82.510 -174.590 ;
        RECT -78.790 -174.880 -78.470 -174.590 ;
        RECT -72.910 -174.880 -72.590 -174.590 ;
        RECT -68.870 -174.880 -68.550 -174.590 ;
        RECT -62.990 -174.880 -62.670 -174.590 ;
        RECT -58.950 -174.880 -58.630 -174.590 ;
        RECT -53.070 -174.880 -52.750 -174.590 ;
        RECT -49.030 -174.880 -48.710 -174.590 ;
        RECT -43.150 -174.880 -42.830 -174.590 ;
        RECT -39.110 -174.880 -38.790 -174.590 ;
        RECT -33.230 -174.880 -32.910 -174.590 ;
        RECT -29.190 -174.880 -28.870 -174.590 ;
        RECT -23.310 -174.880 -22.990 -174.590 ;
        RECT -19.270 -174.880 -18.950 -174.590 ;
        RECT -13.390 -174.880 -13.070 -174.590 ;
        RECT -9.350 -174.880 -9.030 -174.590 ;
        RECT -3.470 -174.880 -3.150 -174.590 ;
        RECT 0.570 -174.880 0.890 -174.590 ;
        RECT 6.450 -174.880 6.770 -174.590 ;
        RECT 10.490 -174.880 10.810 -174.590 ;
        RECT 16.370 -174.880 16.690 -174.590 ;
        RECT 20.410 -174.880 20.730 -174.590 ;
        RECT 26.290 -174.880 26.610 -174.590 ;
        RECT -289.200 -175.680 -287.360 -175.200 ;
        RECT -287.030 -176.010 -286.840 -174.880 ;
        RECT -281.180 -176.010 -280.990 -174.880 ;
        RECT -277.110 -176.010 -276.920 -174.880 ;
        RECT -271.260 -176.010 -271.070 -174.880 ;
        RECT -267.190 -176.010 -267.000 -174.880 ;
        RECT -261.340 -176.010 -261.150 -174.880 ;
        RECT -257.270 -176.010 -257.080 -174.880 ;
        RECT -251.420 -176.010 -251.230 -174.880 ;
        RECT -247.350 -176.010 -247.160 -174.880 ;
        RECT -241.500 -176.010 -241.310 -174.880 ;
        RECT -237.430 -176.010 -237.240 -174.880 ;
        RECT -231.580 -176.010 -231.390 -174.880 ;
        RECT -227.510 -176.010 -227.320 -174.880 ;
        RECT -221.660 -176.010 -221.470 -174.880 ;
        RECT -217.590 -176.010 -217.400 -174.880 ;
        RECT -211.740 -176.010 -211.550 -174.880 ;
        RECT -207.670 -176.010 -207.480 -174.880 ;
        RECT -201.820 -176.010 -201.630 -174.880 ;
        RECT -197.750 -176.010 -197.560 -174.880 ;
        RECT -191.900 -176.010 -191.710 -174.880 ;
        RECT -187.830 -176.010 -187.640 -174.880 ;
        RECT -181.980 -176.010 -181.790 -174.880 ;
        RECT -177.910 -176.010 -177.720 -174.880 ;
        RECT -172.060 -176.010 -171.870 -174.880 ;
        RECT -167.990 -176.010 -167.800 -174.880 ;
        RECT -162.140 -176.010 -161.950 -174.880 ;
        RECT -158.070 -176.010 -157.880 -174.880 ;
        RECT -152.220 -176.010 -152.030 -174.880 ;
        RECT -148.150 -176.010 -147.960 -174.880 ;
        RECT -142.300 -176.010 -142.110 -174.880 ;
        RECT -138.230 -176.010 -138.040 -174.880 ;
        RECT -132.380 -176.010 -132.190 -174.880 ;
        RECT -128.310 -176.010 -128.120 -174.880 ;
        RECT -122.460 -176.010 -122.270 -174.880 ;
        RECT -118.390 -176.010 -118.200 -174.880 ;
        RECT -112.540 -176.010 -112.350 -174.880 ;
        RECT -108.470 -176.010 -108.280 -174.880 ;
        RECT -102.620 -176.010 -102.430 -174.880 ;
        RECT -98.550 -176.010 -98.360 -174.880 ;
        RECT -92.700 -176.010 -92.510 -174.880 ;
        RECT -88.630 -176.010 -88.440 -174.880 ;
        RECT -82.780 -176.010 -82.590 -174.880 ;
        RECT -78.710 -176.010 -78.520 -174.880 ;
        RECT -72.860 -176.010 -72.670 -174.880 ;
        RECT -68.790 -176.010 -68.600 -174.880 ;
        RECT -62.940 -176.010 -62.750 -174.880 ;
        RECT -58.870 -176.010 -58.680 -174.880 ;
        RECT -53.020 -176.010 -52.830 -174.880 ;
        RECT -48.950 -176.010 -48.760 -174.880 ;
        RECT -43.100 -176.010 -42.910 -174.880 ;
        RECT -39.030 -176.010 -38.840 -174.880 ;
        RECT -33.180 -176.010 -32.990 -174.880 ;
        RECT -29.110 -176.010 -28.920 -174.880 ;
        RECT -23.260 -176.010 -23.070 -174.880 ;
        RECT -19.190 -176.010 -19.000 -174.880 ;
        RECT -13.340 -176.010 -13.150 -174.880 ;
        RECT -9.270 -176.010 -9.080 -174.880 ;
        RECT -3.420 -176.010 -3.230 -174.880 ;
        RECT 0.650 -176.010 0.840 -174.880 ;
        RECT 6.500 -176.010 6.690 -174.880 ;
        RECT 10.570 -176.010 10.760 -174.880 ;
        RECT 16.420 -176.010 16.610 -174.880 ;
        RECT 20.490 -176.010 20.680 -174.880 ;
        RECT 26.340 -176.010 26.530 -174.880 ;
        RECT 26.860 -175.680 28.700 -175.200 ;
        RECT -287.790 -176.160 -285.850 -176.010 ;
        RECT -287.790 -176.310 -287.450 -176.160 ;
        RECT -287.790 -176.510 -287.470 -176.480 ;
        RECT -287.790 -176.650 -286.970 -176.510 ;
        RECT -287.790 -176.760 -287.470 -176.650 ;
        RECT -287.130 -177.440 -286.970 -176.650 ;
        RECT -286.010 -176.950 -285.850 -176.160 ;
        RECT -282.170 -176.160 -280.230 -176.010 ;
        RECT -285.510 -176.950 -285.190 -176.840 ;
        RECT -286.010 -177.090 -285.190 -176.950 ;
        RECT -285.510 -177.120 -285.190 -177.090 ;
        RECT -282.830 -176.950 -282.510 -176.840 ;
        RECT -282.170 -176.950 -282.010 -176.160 ;
        RECT -280.570 -176.310 -280.230 -176.160 ;
        RECT -277.870 -176.160 -275.930 -176.010 ;
        RECT -277.870 -176.310 -277.530 -176.160 ;
        RECT -280.550 -176.510 -280.230 -176.480 ;
        RECT -282.830 -177.090 -282.010 -176.950 ;
        RECT -281.050 -176.650 -280.230 -176.510 ;
        RECT -282.830 -177.120 -282.510 -177.090 ;
        RECT -285.530 -177.440 -285.190 -177.290 ;
        RECT -287.130 -177.590 -285.190 -177.440 ;
        RECT -282.830 -177.440 -282.490 -177.290 ;
        RECT -281.050 -177.440 -280.890 -176.650 ;
        RECT -280.550 -176.760 -280.230 -176.650 ;
        RECT -277.870 -176.510 -277.550 -176.480 ;
        RECT -277.870 -176.650 -277.050 -176.510 ;
        RECT -277.870 -176.760 -277.550 -176.650 ;
        RECT -282.830 -177.590 -280.890 -177.440 ;
        RECT -277.210 -177.440 -277.050 -176.650 ;
        RECT -276.090 -176.950 -275.930 -176.160 ;
        RECT -272.250 -176.160 -270.310 -176.010 ;
        RECT -275.590 -176.950 -275.270 -176.840 ;
        RECT -276.090 -177.090 -275.270 -176.950 ;
        RECT -275.590 -177.120 -275.270 -177.090 ;
        RECT -272.910 -176.950 -272.590 -176.840 ;
        RECT -272.250 -176.950 -272.090 -176.160 ;
        RECT -270.650 -176.310 -270.310 -176.160 ;
        RECT -267.950 -176.160 -266.010 -176.010 ;
        RECT -267.950 -176.310 -267.610 -176.160 ;
        RECT -270.630 -176.510 -270.310 -176.480 ;
        RECT -272.910 -177.090 -272.090 -176.950 ;
        RECT -271.130 -176.650 -270.310 -176.510 ;
        RECT -272.910 -177.120 -272.590 -177.090 ;
        RECT -275.610 -177.440 -275.270 -177.290 ;
        RECT -277.210 -177.590 -275.270 -177.440 ;
        RECT -272.910 -177.440 -272.570 -177.290 ;
        RECT -271.130 -177.440 -270.970 -176.650 ;
        RECT -270.630 -176.760 -270.310 -176.650 ;
        RECT -267.950 -176.510 -267.630 -176.480 ;
        RECT -267.950 -176.650 -267.130 -176.510 ;
        RECT -267.950 -176.760 -267.630 -176.650 ;
        RECT -272.910 -177.590 -270.970 -177.440 ;
        RECT -267.290 -177.440 -267.130 -176.650 ;
        RECT -266.170 -176.950 -266.010 -176.160 ;
        RECT -262.330 -176.160 -260.390 -176.010 ;
        RECT -265.670 -176.950 -265.350 -176.840 ;
        RECT -266.170 -177.090 -265.350 -176.950 ;
        RECT -265.670 -177.120 -265.350 -177.090 ;
        RECT -262.990 -176.950 -262.670 -176.840 ;
        RECT -262.330 -176.950 -262.170 -176.160 ;
        RECT -260.730 -176.310 -260.390 -176.160 ;
        RECT -258.030 -176.160 -256.090 -176.010 ;
        RECT -258.030 -176.310 -257.690 -176.160 ;
        RECT -260.710 -176.510 -260.390 -176.480 ;
        RECT -262.990 -177.090 -262.170 -176.950 ;
        RECT -261.210 -176.650 -260.390 -176.510 ;
        RECT -262.990 -177.120 -262.670 -177.090 ;
        RECT -265.690 -177.440 -265.350 -177.290 ;
        RECT -267.290 -177.590 -265.350 -177.440 ;
        RECT -262.990 -177.440 -262.650 -177.290 ;
        RECT -261.210 -177.440 -261.050 -176.650 ;
        RECT -260.710 -176.760 -260.390 -176.650 ;
        RECT -258.030 -176.510 -257.710 -176.480 ;
        RECT -258.030 -176.650 -257.210 -176.510 ;
        RECT -258.030 -176.760 -257.710 -176.650 ;
        RECT -262.990 -177.590 -261.050 -177.440 ;
        RECT -257.370 -177.440 -257.210 -176.650 ;
        RECT -256.250 -176.950 -256.090 -176.160 ;
        RECT -252.410 -176.160 -250.470 -176.010 ;
        RECT -255.750 -176.950 -255.430 -176.840 ;
        RECT -256.250 -177.090 -255.430 -176.950 ;
        RECT -255.750 -177.120 -255.430 -177.090 ;
        RECT -253.070 -176.950 -252.750 -176.840 ;
        RECT -252.410 -176.950 -252.250 -176.160 ;
        RECT -250.810 -176.310 -250.470 -176.160 ;
        RECT -248.110 -176.160 -246.170 -176.010 ;
        RECT -248.110 -176.310 -247.770 -176.160 ;
        RECT -250.790 -176.510 -250.470 -176.480 ;
        RECT -253.070 -177.090 -252.250 -176.950 ;
        RECT -251.290 -176.650 -250.470 -176.510 ;
        RECT -253.070 -177.120 -252.750 -177.090 ;
        RECT -255.770 -177.440 -255.430 -177.290 ;
        RECT -257.370 -177.590 -255.430 -177.440 ;
        RECT -253.070 -177.440 -252.730 -177.290 ;
        RECT -251.290 -177.440 -251.130 -176.650 ;
        RECT -250.790 -176.760 -250.470 -176.650 ;
        RECT -248.110 -176.510 -247.790 -176.480 ;
        RECT -248.110 -176.650 -247.290 -176.510 ;
        RECT -248.110 -176.760 -247.790 -176.650 ;
        RECT -253.070 -177.590 -251.130 -177.440 ;
        RECT -247.450 -177.440 -247.290 -176.650 ;
        RECT -246.330 -176.950 -246.170 -176.160 ;
        RECT -242.490 -176.160 -240.550 -176.010 ;
        RECT -245.830 -176.950 -245.510 -176.840 ;
        RECT -246.330 -177.090 -245.510 -176.950 ;
        RECT -245.830 -177.120 -245.510 -177.090 ;
        RECT -243.150 -176.950 -242.830 -176.840 ;
        RECT -242.490 -176.950 -242.330 -176.160 ;
        RECT -240.890 -176.310 -240.550 -176.160 ;
        RECT -238.190 -176.160 -236.250 -176.010 ;
        RECT -238.190 -176.310 -237.850 -176.160 ;
        RECT -240.870 -176.510 -240.550 -176.480 ;
        RECT -243.150 -177.090 -242.330 -176.950 ;
        RECT -241.370 -176.650 -240.550 -176.510 ;
        RECT -243.150 -177.120 -242.830 -177.090 ;
        RECT -245.850 -177.440 -245.510 -177.290 ;
        RECT -247.450 -177.590 -245.510 -177.440 ;
        RECT -243.150 -177.440 -242.810 -177.290 ;
        RECT -241.370 -177.440 -241.210 -176.650 ;
        RECT -240.870 -176.760 -240.550 -176.650 ;
        RECT -238.190 -176.510 -237.870 -176.480 ;
        RECT -238.190 -176.650 -237.370 -176.510 ;
        RECT -238.190 -176.760 -237.870 -176.650 ;
        RECT -243.150 -177.590 -241.210 -177.440 ;
        RECT -237.530 -177.440 -237.370 -176.650 ;
        RECT -236.410 -176.950 -236.250 -176.160 ;
        RECT -232.570 -176.160 -230.630 -176.010 ;
        RECT -235.910 -176.950 -235.590 -176.840 ;
        RECT -236.410 -177.090 -235.590 -176.950 ;
        RECT -235.910 -177.120 -235.590 -177.090 ;
        RECT -233.230 -176.950 -232.910 -176.840 ;
        RECT -232.570 -176.950 -232.410 -176.160 ;
        RECT -230.970 -176.310 -230.630 -176.160 ;
        RECT -228.270 -176.160 -226.330 -176.010 ;
        RECT -228.270 -176.310 -227.930 -176.160 ;
        RECT -230.950 -176.510 -230.630 -176.480 ;
        RECT -233.230 -177.090 -232.410 -176.950 ;
        RECT -231.450 -176.650 -230.630 -176.510 ;
        RECT -233.230 -177.120 -232.910 -177.090 ;
        RECT -235.930 -177.440 -235.590 -177.290 ;
        RECT -237.530 -177.590 -235.590 -177.440 ;
        RECT -233.230 -177.440 -232.890 -177.290 ;
        RECT -231.450 -177.440 -231.290 -176.650 ;
        RECT -230.950 -176.760 -230.630 -176.650 ;
        RECT -228.270 -176.510 -227.950 -176.480 ;
        RECT -228.270 -176.650 -227.450 -176.510 ;
        RECT -228.270 -176.760 -227.950 -176.650 ;
        RECT -233.230 -177.590 -231.290 -177.440 ;
        RECT -227.610 -177.440 -227.450 -176.650 ;
        RECT -226.490 -176.950 -226.330 -176.160 ;
        RECT -222.650 -176.160 -220.710 -176.010 ;
        RECT -225.990 -176.950 -225.670 -176.840 ;
        RECT -226.490 -177.090 -225.670 -176.950 ;
        RECT -225.990 -177.120 -225.670 -177.090 ;
        RECT -223.310 -176.950 -222.990 -176.840 ;
        RECT -222.650 -176.950 -222.490 -176.160 ;
        RECT -221.050 -176.310 -220.710 -176.160 ;
        RECT -218.350 -176.160 -216.410 -176.010 ;
        RECT -218.350 -176.310 -218.010 -176.160 ;
        RECT -221.030 -176.510 -220.710 -176.480 ;
        RECT -223.310 -177.090 -222.490 -176.950 ;
        RECT -221.530 -176.650 -220.710 -176.510 ;
        RECT -223.310 -177.120 -222.990 -177.090 ;
        RECT -226.010 -177.440 -225.670 -177.290 ;
        RECT -227.610 -177.590 -225.670 -177.440 ;
        RECT -223.310 -177.440 -222.970 -177.290 ;
        RECT -221.530 -177.440 -221.370 -176.650 ;
        RECT -221.030 -176.760 -220.710 -176.650 ;
        RECT -218.350 -176.510 -218.030 -176.480 ;
        RECT -218.350 -176.650 -217.530 -176.510 ;
        RECT -218.350 -176.760 -218.030 -176.650 ;
        RECT -223.310 -177.590 -221.370 -177.440 ;
        RECT -217.690 -177.440 -217.530 -176.650 ;
        RECT -216.570 -176.950 -216.410 -176.160 ;
        RECT -212.730 -176.160 -210.790 -176.010 ;
        RECT -216.070 -176.950 -215.750 -176.840 ;
        RECT -216.570 -177.090 -215.750 -176.950 ;
        RECT -216.070 -177.120 -215.750 -177.090 ;
        RECT -213.390 -176.950 -213.070 -176.840 ;
        RECT -212.730 -176.950 -212.570 -176.160 ;
        RECT -211.130 -176.310 -210.790 -176.160 ;
        RECT -208.430 -176.160 -206.490 -176.010 ;
        RECT -208.430 -176.310 -208.090 -176.160 ;
        RECT -211.110 -176.510 -210.790 -176.480 ;
        RECT -213.390 -177.090 -212.570 -176.950 ;
        RECT -211.610 -176.650 -210.790 -176.510 ;
        RECT -213.390 -177.120 -213.070 -177.090 ;
        RECT -216.090 -177.440 -215.750 -177.290 ;
        RECT -217.690 -177.590 -215.750 -177.440 ;
        RECT -213.390 -177.440 -213.050 -177.290 ;
        RECT -211.610 -177.440 -211.450 -176.650 ;
        RECT -211.110 -176.760 -210.790 -176.650 ;
        RECT -208.430 -176.510 -208.110 -176.480 ;
        RECT -208.430 -176.650 -207.610 -176.510 ;
        RECT -208.430 -176.760 -208.110 -176.650 ;
        RECT -213.390 -177.590 -211.450 -177.440 ;
        RECT -207.770 -177.440 -207.610 -176.650 ;
        RECT -206.650 -176.950 -206.490 -176.160 ;
        RECT -202.810 -176.160 -200.870 -176.010 ;
        RECT -206.150 -176.950 -205.830 -176.840 ;
        RECT -206.650 -177.090 -205.830 -176.950 ;
        RECT -206.150 -177.120 -205.830 -177.090 ;
        RECT -203.470 -176.950 -203.150 -176.840 ;
        RECT -202.810 -176.950 -202.650 -176.160 ;
        RECT -201.210 -176.310 -200.870 -176.160 ;
        RECT -198.510 -176.160 -196.570 -176.010 ;
        RECT -198.510 -176.310 -198.170 -176.160 ;
        RECT -201.190 -176.510 -200.870 -176.480 ;
        RECT -203.470 -177.090 -202.650 -176.950 ;
        RECT -201.690 -176.650 -200.870 -176.510 ;
        RECT -203.470 -177.120 -203.150 -177.090 ;
        RECT -206.170 -177.440 -205.830 -177.290 ;
        RECT -207.770 -177.590 -205.830 -177.440 ;
        RECT -203.470 -177.440 -203.130 -177.290 ;
        RECT -201.690 -177.440 -201.530 -176.650 ;
        RECT -201.190 -176.760 -200.870 -176.650 ;
        RECT -198.510 -176.510 -198.190 -176.480 ;
        RECT -198.510 -176.650 -197.690 -176.510 ;
        RECT -198.510 -176.760 -198.190 -176.650 ;
        RECT -203.470 -177.590 -201.530 -177.440 ;
        RECT -197.850 -177.440 -197.690 -176.650 ;
        RECT -196.730 -176.950 -196.570 -176.160 ;
        RECT -192.890 -176.160 -190.950 -176.010 ;
        RECT -196.230 -176.950 -195.910 -176.840 ;
        RECT -196.730 -177.090 -195.910 -176.950 ;
        RECT -196.230 -177.120 -195.910 -177.090 ;
        RECT -193.550 -176.950 -193.230 -176.840 ;
        RECT -192.890 -176.950 -192.730 -176.160 ;
        RECT -191.290 -176.310 -190.950 -176.160 ;
        RECT -188.590 -176.160 -186.650 -176.010 ;
        RECT -188.590 -176.310 -188.250 -176.160 ;
        RECT -191.270 -176.510 -190.950 -176.480 ;
        RECT -193.550 -177.090 -192.730 -176.950 ;
        RECT -191.770 -176.650 -190.950 -176.510 ;
        RECT -193.550 -177.120 -193.230 -177.090 ;
        RECT -196.250 -177.440 -195.910 -177.290 ;
        RECT -197.850 -177.590 -195.910 -177.440 ;
        RECT -193.550 -177.440 -193.210 -177.290 ;
        RECT -191.770 -177.440 -191.610 -176.650 ;
        RECT -191.270 -176.760 -190.950 -176.650 ;
        RECT -188.590 -176.510 -188.270 -176.480 ;
        RECT -188.590 -176.650 -187.770 -176.510 ;
        RECT -188.590 -176.760 -188.270 -176.650 ;
        RECT -193.550 -177.590 -191.610 -177.440 ;
        RECT -187.930 -177.440 -187.770 -176.650 ;
        RECT -186.810 -176.950 -186.650 -176.160 ;
        RECT -182.970 -176.160 -181.030 -176.010 ;
        RECT -186.310 -176.950 -185.990 -176.840 ;
        RECT -186.810 -177.090 -185.990 -176.950 ;
        RECT -186.310 -177.120 -185.990 -177.090 ;
        RECT -183.630 -176.950 -183.310 -176.840 ;
        RECT -182.970 -176.950 -182.810 -176.160 ;
        RECT -181.370 -176.310 -181.030 -176.160 ;
        RECT -178.670 -176.160 -176.730 -176.010 ;
        RECT -178.670 -176.310 -178.330 -176.160 ;
        RECT -181.350 -176.510 -181.030 -176.480 ;
        RECT -183.630 -177.090 -182.810 -176.950 ;
        RECT -181.850 -176.650 -181.030 -176.510 ;
        RECT -183.630 -177.120 -183.310 -177.090 ;
        RECT -186.330 -177.440 -185.990 -177.290 ;
        RECT -187.930 -177.590 -185.990 -177.440 ;
        RECT -183.630 -177.440 -183.290 -177.290 ;
        RECT -181.850 -177.440 -181.690 -176.650 ;
        RECT -181.350 -176.760 -181.030 -176.650 ;
        RECT -178.670 -176.510 -178.350 -176.480 ;
        RECT -178.670 -176.650 -177.850 -176.510 ;
        RECT -178.670 -176.760 -178.350 -176.650 ;
        RECT -183.630 -177.590 -181.690 -177.440 ;
        RECT -178.010 -177.440 -177.850 -176.650 ;
        RECT -176.890 -176.950 -176.730 -176.160 ;
        RECT -173.050 -176.160 -171.110 -176.010 ;
        RECT -176.390 -176.950 -176.070 -176.840 ;
        RECT -176.890 -177.090 -176.070 -176.950 ;
        RECT -176.390 -177.120 -176.070 -177.090 ;
        RECT -173.710 -176.950 -173.390 -176.840 ;
        RECT -173.050 -176.950 -172.890 -176.160 ;
        RECT -171.450 -176.310 -171.110 -176.160 ;
        RECT -168.750 -176.160 -166.810 -176.010 ;
        RECT -168.750 -176.310 -168.410 -176.160 ;
        RECT -171.430 -176.510 -171.110 -176.480 ;
        RECT -173.710 -177.090 -172.890 -176.950 ;
        RECT -171.930 -176.650 -171.110 -176.510 ;
        RECT -173.710 -177.120 -173.390 -177.090 ;
        RECT -176.410 -177.440 -176.070 -177.290 ;
        RECT -178.010 -177.590 -176.070 -177.440 ;
        RECT -173.710 -177.440 -173.370 -177.290 ;
        RECT -171.930 -177.440 -171.770 -176.650 ;
        RECT -171.430 -176.760 -171.110 -176.650 ;
        RECT -168.750 -176.510 -168.430 -176.480 ;
        RECT -168.750 -176.650 -167.930 -176.510 ;
        RECT -168.750 -176.760 -168.430 -176.650 ;
        RECT -173.710 -177.590 -171.770 -177.440 ;
        RECT -168.090 -177.440 -167.930 -176.650 ;
        RECT -166.970 -176.950 -166.810 -176.160 ;
        RECT -163.130 -176.160 -161.190 -176.010 ;
        RECT -166.470 -176.950 -166.150 -176.840 ;
        RECT -166.970 -177.090 -166.150 -176.950 ;
        RECT -166.470 -177.120 -166.150 -177.090 ;
        RECT -163.790 -176.950 -163.470 -176.840 ;
        RECT -163.130 -176.950 -162.970 -176.160 ;
        RECT -161.530 -176.310 -161.190 -176.160 ;
        RECT -158.830 -176.160 -156.890 -176.010 ;
        RECT -158.830 -176.310 -158.490 -176.160 ;
        RECT -161.510 -176.510 -161.190 -176.480 ;
        RECT -163.790 -177.090 -162.970 -176.950 ;
        RECT -162.010 -176.650 -161.190 -176.510 ;
        RECT -163.790 -177.120 -163.470 -177.090 ;
        RECT -166.490 -177.440 -166.150 -177.290 ;
        RECT -168.090 -177.590 -166.150 -177.440 ;
        RECT -163.790 -177.440 -163.450 -177.290 ;
        RECT -162.010 -177.440 -161.850 -176.650 ;
        RECT -161.510 -176.760 -161.190 -176.650 ;
        RECT -158.830 -176.510 -158.510 -176.480 ;
        RECT -158.830 -176.650 -158.010 -176.510 ;
        RECT -158.830 -176.760 -158.510 -176.650 ;
        RECT -163.790 -177.590 -161.850 -177.440 ;
        RECT -158.170 -177.440 -158.010 -176.650 ;
        RECT -157.050 -176.950 -156.890 -176.160 ;
        RECT -153.210 -176.160 -151.270 -176.010 ;
        RECT -156.550 -176.950 -156.230 -176.840 ;
        RECT -157.050 -177.090 -156.230 -176.950 ;
        RECT -156.550 -177.120 -156.230 -177.090 ;
        RECT -153.870 -176.950 -153.550 -176.840 ;
        RECT -153.210 -176.950 -153.050 -176.160 ;
        RECT -151.610 -176.310 -151.270 -176.160 ;
        RECT -148.910 -176.160 -146.970 -176.010 ;
        RECT -148.910 -176.310 -148.570 -176.160 ;
        RECT -151.590 -176.510 -151.270 -176.480 ;
        RECT -153.870 -177.090 -153.050 -176.950 ;
        RECT -152.090 -176.650 -151.270 -176.510 ;
        RECT -153.870 -177.120 -153.550 -177.090 ;
        RECT -156.570 -177.440 -156.230 -177.290 ;
        RECT -158.170 -177.590 -156.230 -177.440 ;
        RECT -153.870 -177.440 -153.530 -177.290 ;
        RECT -152.090 -177.440 -151.930 -176.650 ;
        RECT -151.590 -176.760 -151.270 -176.650 ;
        RECT -148.910 -176.510 -148.590 -176.480 ;
        RECT -148.910 -176.650 -148.090 -176.510 ;
        RECT -148.910 -176.760 -148.590 -176.650 ;
        RECT -153.870 -177.590 -151.930 -177.440 ;
        RECT -148.250 -177.440 -148.090 -176.650 ;
        RECT -147.130 -176.950 -146.970 -176.160 ;
        RECT -143.290 -176.160 -141.350 -176.010 ;
        RECT -146.630 -176.950 -146.310 -176.840 ;
        RECT -147.130 -177.090 -146.310 -176.950 ;
        RECT -146.630 -177.120 -146.310 -177.090 ;
        RECT -143.950 -176.950 -143.630 -176.840 ;
        RECT -143.290 -176.950 -143.130 -176.160 ;
        RECT -141.690 -176.310 -141.350 -176.160 ;
        RECT -138.990 -176.160 -137.050 -176.010 ;
        RECT -138.990 -176.310 -138.650 -176.160 ;
        RECT -141.670 -176.510 -141.350 -176.480 ;
        RECT -143.950 -177.090 -143.130 -176.950 ;
        RECT -142.170 -176.650 -141.350 -176.510 ;
        RECT -143.950 -177.120 -143.630 -177.090 ;
        RECT -146.650 -177.440 -146.310 -177.290 ;
        RECT -148.250 -177.590 -146.310 -177.440 ;
        RECT -143.950 -177.440 -143.610 -177.290 ;
        RECT -142.170 -177.440 -142.010 -176.650 ;
        RECT -141.670 -176.760 -141.350 -176.650 ;
        RECT -138.990 -176.510 -138.670 -176.480 ;
        RECT -138.990 -176.650 -138.170 -176.510 ;
        RECT -138.990 -176.760 -138.670 -176.650 ;
        RECT -143.950 -177.590 -142.010 -177.440 ;
        RECT -138.330 -177.440 -138.170 -176.650 ;
        RECT -137.210 -176.950 -137.050 -176.160 ;
        RECT -133.370 -176.160 -131.430 -176.010 ;
        RECT -136.710 -176.950 -136.390 -176.840 ;
        RECT -137.210 -177.090 -136.390 -176.950 ;
        RECT -136.710 -177.120 -136.390 -177.090 ;
        RECT -134.030 -176.950 -133.710 -176.840 ;
        RECT -133.370 -176.950 -133.210 -176.160 ;
        RECT -131.770 -176.310 -131.430 -176.160 ;
        RECT -129.070 -176.160 -127.130 -176.010 ;
        RECT -129.070 -176.310 -128.730 -176.160 ;
        RECT -131.750 -176.510 -131.430 -176.480 ;
        RECT -134.030 -177.090 -133.210 -176.950 ;
        RECT -132.250 -176.650 -131.430 -176.510 ;
        RECT -134.030 -177.120 -133.710 -177.090 ;
        RECT -136.730 -177.440 -136.390 -177.290 ;
        RECT -138.330 -177.590 -136.390 -177.440 ;
        RECT -134.030 -177.440 -133.690 -177.290 ;
        RECT -132.250 -177.440 -132.090 -176.650 ;
        RECT -131.750 -176.760 -131.430 -176.650 ;
        RECT -129.070 -176.510 -128.750 -176.480 ;
        RECT -129.070 -176.650 -128.250 -176.510 ;
        RECT -129.070 -176.760 -128.750 -176.650 ;
        RECT -134.030 -177.590 -132.090 -177.440 ;
        RECT -128.410 -177.440 -128.250 -176.650 ;
        RECT -127.290 -176.950 -127.130 -176.160 ;
        RECT -123.450 -176.160 -121.510 -176.010 ;
        RECT -126.790 -176.950 -126.470 -176.840 ;
        RECT -127.290 -177.090 -126.470 -176.950 ;
        RECT -126.790 -177.120 -126.470 -177.090 ;
        RECT -124.110 -176.950 -123.790 -176.840 ;
        RECT -123.450 -176.950 -123.290 -176.160 ;
        RECT -121.850 -176.310 -121.510 -176.160 ;
        RECT -119.150 -176.160 -117.210 -176.010 ;
        RECT -119.150 -176.310 -118.810 -176.160 ;
        RECT -121.830 -176.510 -121.510 -176.480 ;
        RECT -124.110 -177.090 -123.290 -176.950 ;
        RECT -122.330 -176.650 -121.510 -176.510 ;
        RECT -124.110 -177.120 -123.790 -177.090 ;
        RECT -126.810 -177.440 -126.470 -177.290 ;
        RECT -128.410 -177.590 -126.470 -177.440 ;
        RECT -124.110 -177.440 -123.770 -177.290 ;
        RECT -122.330 -177.440 -122.170 -176.650 ;
        RECT -121.830 -176.760 -121.510 -176.650 ;
        RECT -119.150 -176.510 -118.830 -176.480 ;
        RECT -119.150 -176.650 -118.330 -176.510 ;
        RECT -119.150 -176.760 -118.830 -176.650 ;
        RECT -124.110 -177.590 -122.170 -177.440 ;
        RECT -118.490 -177.440 -118.330 -176.650 ;
        RECT -117.370 -176.950 -117.210 -176.160 ;
        RECT -113.530 -176.160 -111.590 -176.010 ;
        RECT -116.870 -176.950 -116.550 -176.840 ;
        RECT -117.370 -177.090 -116.550 -176.950 ;
        RECT -116.870 -177.120 -116.550 -177.090 ;
        RECT -114.190 -176.950 -113.870 -176.840 ;
        RECT -113.530 -176.950 -113.370 -176.160 ;
        RECT -111.930 -176.310 -111.590 -176.160 ;
        RECT -109.230 -176.160 -107.290 -176.010 ;
        RECT -109.230 -176.310 -108.890 -176.160 ;
        RECT -111.910 -176.510 -111.590 -176.480 ;
        RECT -114.190 -177.090 -113.370 -176.950 ;
        RECT -112.410 -176.650 -111.590 -176.510 ;
        RECT -114.190 -177.120 -113.870 -177.090 ;
        RECT -116.890 -177.440 -116.550 -177.290 ;
        RECT -118.490 -177.590 -116.550 -177.440 ;
        RECT -114.190 -177.440 -113.850 -177.290 ;
        RECT -112.410 -177.440 -112.250 -176.650 ;
        RECT -111.910 -176.760 -111.590 -176.650 ;
        RECT -109.230 -176.510 -108.910 -176.480 ;
        RECT -109.230 -176.650 -108.410 -176.510 ;
        RECT -109.230 -176.760 -108.910 -176.650 ;
        RECT -114.190 -177.590 -112.250 -177.440 ;
        RECT -108.570 -177.440 -108.410 -176.650 ;
        RECT -107.450 -176.950 -107.290 -176.160 ;
        RECT -103.610 -176.160 -101.670 -176.010 ;
        RECT -106.950 -176.950 -106.630 -176.840 ;
        RECT -107.450 -177.090 -106.630 -176.950 ;
        RECT -106.950 -177.120 -106.630 -177.090 ;
        RECT -104.270 -176.950 -103.950 -176.840 ;
        RECT -103.610 -176.950 -103.450 -176.160 ;
        RECT -102.010 -176.310 -101.670 -176.160 ;
        RECT -99.310 -176.160 -97.370 -176.010 ;
        RECT -99.310 -176.310 -98.970 -176.160 ;
        RECT -101.990 -176.510 -101.670 -176.480 ;
        RECT -104.270 -177.090 -103.450 -176.950 ;
        RECT -102.490 -176.650 -101.670 -176.510 ;
        RECT -104.270 -177.120 -103.950 -177.090 ;
        RECT -106.970 -177.440 -106.630 -177.290 ;
        RECT -108.570 -177.590 -106.630 -177.440 ;
        RECT -104.270 -177.440 -103.930 -177.290 ;
        RECT -102.490 -177.440 -102.330 -176.650 ;
        RECT -101.990 -176.760 -101.670 -176.650 ;
        RECT -99.310 -176.510 -98.990 -176.480 ;
        RECT -99.310 -176.650 -98.490 -176.510 ;
        RECT -99.310 -176.760 -98.990 -176.650 ;
        RECT -104.270 -177.590 -102.330 -177.440 ;
        RECT -98.650 -177.440 -98.490 -176.650 ;
        RECT -97.530 -176.950 -97.370 -176.160 ;
        RECT -93.690 -176.160 -91.750 -176.010 ;
        RECT -97.030 -176.950 -96.710 -176.840 ;
        RECT -97.530 -177.090 -96.710 -176.950 ;
        RECT -97.030 -177.120 -96.710 -177.090 ;
        RECT -94.350 -176.950 -94.030 -176.840 ;
        RECT -93.690 -176.950 -93.530 -176.160 ;
        RECT -92.090 -176.310 -91.750 -176.160 ;
        RECT -89.390 -176.160 -87.450 -176.010 ;
        RECT -89.390 -176.310 -89.050 -176.160 ;
        RECT -92.070 -176.510 -91.750 -176.480 ;
        RECT -94.350 -177.090 -93.530 -176.950 ;
        RECT -92.570 -176.650 -91.750 -176.510 ;
        RECT -94.350 -177.120 -94.030 -177.090 ;
        RECT -97.050 -177.440 -96.710 -177.290 ;
        RECT -98.650 -177.590 -96.710 -177.440 ;
        RECT -94.350 -177.440 -94.010 -177.290 ;
        RECT -92.570 -177.440 -92.410 -176.650 ;
        RECT -92.070 -176.760 -91.750 -176.650 ;
        RECT -89.390 -176.510 -89.070 -176.480 ;
        RECT -89.390 -176.650 -88.570 -176.510 ;
        RECT -89.390 -176.760 -89.070 -176.650 ;
        RECT -94.350 -177.590 -92.410 -177.440 ;
        RECT -88.730 -177.440 -88.570 -176.650 ;
        RECT -87.610 -176.950 -87.450 -176.160 ;
        RECT -83.770 -176.160 -81.830 -176.010 ;
        RECT -87.110 -176.950 -86.790 -176.840 ;
        RECT -87.610 -177.090 -86.790 -176.950 ;
        RECT -87.110 -177.120 -86.790 -177.090 ;
        RECT -84.430 -176.950 -84.110 -176.840 ;
        RECT -83.770 -176.950 -83.610 -176.160 ;
        RECT -82.170 -176.310 -81.830 -176.160 ;
        RECT -79.470 -176.160 -77.530 -176.010 ;
        RECT -79.470 -176.310 -79.130 -176.160 ;
        RECT -82.150 -176.510 -81.830 -176.480 ;
        RECT -84.430 -177.090 -83.610 -176.950 ;
        RECT -82.650 -176.650 -81.830 -176.510 ;
        RECT -84.430 -177.120 -84.110 -177.090 ;
        RECT -87.130 -177.440 -86.790 -177.290 ;
        RECT -88.730 -177.590 -86.790 -177.440 ;
        RECT -84.430 -177.440 -84.090 -177.290 ;
        RECT -82.650 -177.440 -82.490 -176.650 ;
        RECT -82.150 -176.760 -81.830 -176.650 ;
        RECT -79.470 -176.510 -79.150 -176.480 ;
        RECT -79.470 -176.650 -78.650 -176.510 ;
        RECT -79.470 -176.760 -79.150 -176.650 ;
        RECT -84.430 -177.590 -82.490 -177.440 ;
        RECT -78.810 -177.440 -78.650 -176.650 ;
        RECT -77.690 -176.950 -77.530 -176.160 ;
        RECT -73.850 -176.160 -71.910 -176.010 ;
        RECT -77.190 -176.950 -76.870 -176.840 ;
        RECT -77.690 -177.090 -76.870 -176.950 ;
        RECT -77.190 -177.120 -76.870 -177.090 ;
        RECT -74.510 -176.950 -74.190 -176.840 ;
        RECT -73.850 -176.950 -73.690 -176.160 ;
        RECT -72.250 -176.310 -71.910 -176.160 ;
        RECT -69.550 -176.160 -67.610 -176.010 ;
        RECT -69.550 -176.310 -69.210 -176.160 ;
        RECT -72.230 -176.510 -71.910 -176.480 ;
        RECT -74.510 -177.090 -73.690 -176.950 ;
        RECT -72.730 -176.650 -71.910 -176.510 ;
        RECT -74.510 -177.120 -74.190 -177.090 ;
        RECT -77.210 -177.440 -76.870 -177.290 ;
        RECT -78.810 -177.590 -76.870 -177.440 ;
        RECT -74.510 -177.440 -74.170 -177.290 ;
        RECT -72.730 -177.440 -72.570 -176.650 ;
        RECT -72.230 -176.760 -71.910 -176.650 ;
        RECT -69.550 -176.510 -69.230 -176.480 ;
        RECT -69.550 -176.650 -68.730 -176.510 ;
        RECT -69.550 -176.760 -69.230 -176.650 ;
        RECT -74.510 -177.590 -72.570 -177.440 ;
        RECT -68.890 -177.440 -68.730 -176.650 ;
        RECT -67.770 -176.950 -67.610 -176.160 ;
        RECT -63.930 -176.160 -61.990 -176.010 ;
        RECT -67.270 -176.950 -66.950 -176.840 ;
        RECT -67.770 -177.090 -66.950 -176.950 ;
        RECT -67.270 -177.120 -66.950 -177.090 ;
        RECT -64.590 -176.950 -64.270 -176.840 ;
        RECT -63.930 -176.950 -63.770 -176.160 ;
        RECT -62.330 -176.310 -61.990 -176.160 ;
        RECT -59.630 -176.160 -57.690 -176.010 ;
        RECT -59.630 -176.310 -59.290 -176.160 ;
        RECT -62.310 -176.510 -61.990 -176.480 ;
        RECT -64.590 -177.090 -63.770 -176.950 ;
        RECT -62.810 -176.650 -61.990 -176.510 ;
        RECT -64.590 -177.120 -64.270 -177.090 ;
        RECT -67.290 -177.440 -66.950 -177.290 ;
        RECT -68.890 -177.590 -66.950 -177.440 ;
        RECT -64.590 -177.440 -64.250 -177.290 ;
        RECT -62.810 -177.440 -62.650 -176.650 ;
        RECT -62.310 -176.760 -61.990 -176.650 ;
        RECT -59.630 -176.510 -59.310 -176.480 ;
        RECT -59.630 -176.650 -58.810 -176.510 ;
        RECT -59.630 -176.760 -59.310 -176.650 ;
        RECT -64.590 -177.590 -62.650 -177.440 ;
        RECT -58.970 -177.440 -58.810 -176.650 ;
        RECT -57.850 -176.950 -57.690 -176.160 ;
        RECT -54.010 -176.160 -52.070 -176.010 ;
        RECT -57.350 -176.950 -57.030 -176.840 ;
        RECT -57.850 -177.090 -57.030 -176.950 ;
        RECT -57.350 -177.120 -57.030 -177.090 ;
        RECT -54.670 -176.950 -54.350 -176.840 ;
        RECT -54.010 -176.950 -53.850 -176.160 ;
        RECT -52.410 -176.310 -52.070 -176.160 ;
        RECT -49.710 -176.160 -47.770 -176.010 ;
        RECT -49.710 -176.310 -49.370 -176.160 ;
        RECT -52.390 -176.510 -52.070 -176.480 ;
        RECT -54.670 -177.090 -53.850 -176.950 ;
        RECT -52.890 -176.650 -52.070 -176.510 ;
        RECT -54.670 -177.120 -54.350 -177.090 ;
        RECT -57.370 -177.440 -57.030 -177.290 ;
        RECT -58.970 -177.590 -57.030 -177.440 ;
        RECT -54.670 -177.440 -54.330 -177.290 ;
        RECT -52.890 -177.440 -52.730 -176.650 ;
        RECT -52.390 -176.760 -52.070 -176.650 ;
        RECT -49.710 -176.510 -49.390 -176.480 ;
        RECT -49.710 -176.650 -48.890 -176.510 ;
        RECT -49.710 -176.760 -49.390 -176.650 ;
        RECT -54.670 -177.590 -52.730 -177.440 ;
        RECT -49.050 -177.440 -48.890 -176.650 ;
        RECT -47.930 -176.950 -47.770 -176.160 ;
        RECT -44.090 -176.160 -42.150 -176.010 ;
        RECT -47.430 -176.950 -47.110 -176.840 ;
        RECT -47.930 -177.090 -47.110 -176.950 ;
        RECT -47.430 -177.120 -47.110 -177.090 ;
        RECT -44.750 -176.950 -44.430 -176.840 ;
        RECT -44.090 -176.950 -43.930 -176.160 ;
        RECT -42.490 -176.310 -42.150 -176.160 ;
        RECT -39.790 -176.160 -37.850 -176.010 ;
        RECT -39.790 -176.310 -39.450 -176.160 ;
        RECT -42.470 -176.510 -42.150 -176.480 ;
        RECT -44.750 -177.090 -43.930 -176.950 ;
        RECT -42.970 -176.650 -42.150 -176.510 ;
        RECT -44.750 -177.120 -44.430 -177.090 ;
        RECT -47.450 -177.440 -47.110 -177.290 ;
        RECT -49.050 -177.590 -47.110 -177.440 ;
        RECT -44.750 -177.440 -44.410 -177.290 ;
        RECT -42.970 -177.440 -42.810 -176.650 ;
        RECT -42.470 -176.760 -42.150 -176.650 ;
        RECT -39.790 -176.510 -39.470 -176.480 ;
        RECT -39.790 -176.650 -38.970 -176.510 ;
        RECT -39.790 -176.760 -39.470 -176.650 ;
        RECT -44.750 -177.590 -42.810 -177.440 ;
        RECT -39.130 -177.440 -38.970 -176.650 ;
        RECT -38.010 -176.950 -37.850 -176.160 ;
        RECT -34.170 -176.160 -32.230 -176.010 ;
        RECT -37.510 -176.950 -37.190 -176.840 ;
        RECT -38.010 -177.090 -37.190 -176.950 ;
        RECT -37.510 -177.120 -37.190 -177.090 ;
        RECT -34.830 -176.950 -34.510 -176.840 ;
        RECT -34.170 -176.950 -34.010 -176.160 ;
        RECT -32.570 -176.310 -32.230 -176.160 ;
        RECT -29.870 -176.160 -27.930 -176.010 ;
        RECT -29.870 -176.310 -29.530 -176.160 ;
        RECT -32.550 -176.510 -32.230 -176.480 ;
        RECT -34.830 -177.090 -34.010 -176.950 ;
        RECT -33.050 -176.650 -32.230 -176.510 ;
        RECT -34.830 -177.120 -34.510 -177.090 ;
        RECT -37.530 -177.440 -37.190 -177.290 ;
        RECT -39.130 -177.590 -37.190 -177.440 ;
        RECT -34.830 -177.440 -34.490 -177.290 ;
        RECT -33.050 -177.440 -32.890 -176.650 ;
        RECT -32.550 -176.760 -32.230 -176.650 ;
        RECT -29.870 -176.510 -29.550 -176.480 ;
        RECT -29.870 -176.650 -29.050 -176.510 ;
        RECT -29.870 -176.760 -29.550 -176.650 ;
        RECT -34.830 -177.590 -32.890 -177.440 ;
        RECT -29.210 -177.440 -29.050 -176.650 ;
        RECT -28.090 -176.950 -27.930 -176.160 ;
        RECT -24.250 -176.160 -22.310 -176.010 ;
        RECT -27.590 -176.950 -27.270 -176.840 ;
        RECT -28.090 -177.090 -27.270 -176.950 ;
        RECT -27.590 -177.120 -27.270 -177.090 ;
        RECT -24.910 -176.950 -24.590 -176.840 ;
        RECT -24.250 -176.950 -24.090 -176.160 ;
        RECT -22.650 -176.310 -22.310 -176.160 ;
        RECT -19.950 -176.160 -18.010 -176.010 ;
        RECT -19.950 -176.310 -19.610 -176.160 ;
        RECT -22.630 -176.510 -22.310 -176.480 ;
        RECT -24.910 -177.090 -24.090 -176.950 ;
        RECT -23.130 -176.650 -22.310 -176.510 ;
        RECT -24.910 -177.120 -24.590 -177.090 ;
        RECT -27.610 -177.440 -27.270 -177.290 ;
        RECT -29.210 -177.590 -27.270 -177.440 ;
        RECT -24.910 -177.440 -24.570 -177.290 ;
        RECT -23.130 -177.440 -22.970 -176.650 ;
        RECT -22.630 -176.760 -22.310 -176.650 ;
        RECT -19.950 -176.510 -19.630 -176.480 ;
        RECT -19.950 -176.650 -19.130 -176.510 ;
        RECT -19.950 -176.760 -19.630 -176.650 ;
        RECT -24.910 -177.590 -22.970 -177.440 ;
        RECT -19.290 -177.440 -19.130 -176.650 ;
        RECT -18.170 -176.950 -18.010 -176.160 ;
        RECT -14.330 -176.160 -12.390 -176.010 ;
        RECT -17.670 -176.950 -17.350 -176.840 ;
        RECT -18.170 -177.090 -17.350 -176.950 ;
        RECT -17.670 -177.120 -17.350 -177.090 ;
        RECT -14.990 -176.950 -14.670 -176.840 ;
        RECT -14.330 -176.950 -14.170 -176.160 ;
        RECT -12.730 -176.310 -12.390 -176.160 ;
        RECT -10.030 -176.160 -8.090 -176.010 ;
        RECT -10.030 -176.310 -9.690 -176.160 ;
        RECT -12.710 -176.510 -12.390 -176.480 ;
        RECT -14.990 -177.090 -14.170 -176.950 ;
        RECT -13.210 -176.650 -12.390 -176.510 ;
        RECT -14.990 -177.120 -14.670 -177.090 ;
        RECT -17.690 -177.440 -17.350 -177.290 ;
        RECT -19.290 -177.590 -17.350 -177.440 ;
        RECT -14.990 -177.440 -14.650 -177.290 ;
        RECT -13.210 -177.440 -13.050 -176.650 ;
        RECT -12.710 -176.760 -12.390 -176.650 ;
        RECT -10.030 -176.510 -9.710 -176.480 ;
        RECT -10.030 -176.650 -9.210 -176.510 ;
        RECT -10.030 -176.760 -9.710 -176.650 ;
        RECT -14.990 -177.590 -13.050 -177.440 ;
        RECT -9.370 -177.440 -9.210 -176.650 ;
        RECT -8.250 -176.950 -8.090 -176.160 ;
        RECT -4.410 -176.160 -2.470 -176.010 ;
        RECT -7.750 -176.950 -7.430 -176.840 ;
        RECT -8.250 -177.090 -7.430 -176.950 ;
        RECT -7.750 -177.120 -7.430 -177.090 ;
        RECT -5.070 -176.950 -4.750 -176.840 ;
        RECT -4.410 -176.950 -4.250 -176.160 ;
        RECT -2.810 -176.310 -2.470 -176.160 ;
        RECT -0.110 -176.160 1.830 -176.010 ;
        RECT -0.110 -176.310 0.230 -176.160 ;
        RECT -2.790 -176.510 -2.470 -176.480 ;
        RECT -5.070 -177.090 -4.250 -176.950 ;
        RECT -3.290 -176.650 -2.470 -176.510 ;
        RECT -5.070 -177.120 -4.750 -177.090 ;
        RECT -7.770 -177.440 -7.430 -177.290 ;
        RECT -9.370 -177.590 -7.430 -177.440 ;
        RECT -5.070 -177.440 -4.730 -177.290 ;
        RECT -3.290 -177.440 -3.130 -176.650 ;
        RECT -2.790 -176.760 -2.470 -176.650 ;
        RECT -0.110 -176.510 0.210 -176.480 ;
        RECT -0.110 -176.650 0.710 -176.510 ;
        RECT -0.110 -176.760 0.210 -176.650 ;
        RECT -5.070 -177.590 -3.130 -177.440 ;
        RECT 0.550 -177.440 0.710 -176.650 ;
        RECT 1.670 -176.950 1.830 -176.160 ;
        RECT 5.510 -176.160 7.450 -176.010 ;
        RECT 2.170 -176.950 2.490 -176.840 ;
        RECT 1.670 -177.090 2.490 -176.950 ;
        RECT 2.170 -177.120 2.490 -177.090 ;
        RECT 4.850 -176.950 5.170 -176.840 ;
        RECT 5.510 -176.950 5.670 -176.160 ;
        RECT 7.110 -176.310 7.450 -176.160 ;
        RECT 9.810 -176.160 11.750 -176.010 ;
        RECT 9.810 -176.310 10.150 -176.160 ;
        RECT 7.130 -176.510 7.450 -176.480 ;
        RECT 4.850 -177.090 5.670 -176.950 ;
        RECT 6.630 -176.650 7.450 -176.510 ;
        RECT 4.850 -177.120 5.170 -177.090 ;
        RECT 2.150 -177.440 2.490 -177.290 ;
        RECT 0.550 -177.590 2.490 -177.440 ;
        RECT 4.850 -177.440 5.190 -177.290 ;
        RECT 6.630 -177.440 6.790 -176.650 ;
        RECT 7.130 -176.760 7.450 -176.650 ;
        RECT 9.810 -176.510 10.130 -176.480 ;
        RECT 9.810 -176.650 10.630 -176.510 ;
        RECT 9.810 -176.760 10.130 -176.650 ;
        RECT 4.850 -177.590 6.790 -177.440 ;
        RECT 10.470 -177.440 10.630 -176.650 ;
        RECT 11.590 -176.950 11.750 -176.160 ;
        RECT 15.430 -176.160 17.370 -176.010 ;
        RECT 12.090 -176.950 12.410 -176.840 ;
        RECT 11.590 -177.090 12.410 -176.950 ;
        RECT 12.090 -177.120 12.410 -177.090 ;
        RECT 14.770 -176.950 15.090 -176.840 ;
        RECT 15.430 -176.950 15.590 -176.160 ;
        RECT 17.030 -176.310 17.370 -176.160 ;
        RECT 19.730 -176.160 21.670 -176.010 ;
        RECT 19.730 -176.310 20.070 -176.160 ;
        RECT 17.050 -176.510 17.370 -176.480 ;
        RECT 14.770 -177.090 15.590 -176.950 ;
        RECT 16.550 -176.650 17.370 -176.510 ;
        RECT 14.770 -177.120 15.090 -177.090 ;
        RECT 12.070 -177.440 12.410 -177.290 ;
        RECT 10.470 -177.590 12.410 -177.440 ;
        RECT 14.770 -177.440 15.110 -177.290 ;
        RECT 16.550 -177.440 16.710 -176.650 ;
        RECT 17.050 -176.760 17.370 -176.650 ;
        RECT 19.730 -176.510 20.050 -176.480 ;
        RECT 19.730 -176.650 20.550 -176.510 ;
        RECT 19.730 -176.760 20.050 -176.650 ;
        RECT 14.770 -177.590 16.710 -177.440 ;
        RECT 20.390 -177.440 20.550 -176.650 ;
        RECT 21.510 -176.950 21.670 -176.160 ;
        RECT 25.350 -176.160 27.290 -176.010 ;
        RECT 22.010 -176.950 22.330 -176.840 ;
        RECT 21.510 -177.090 22.330 -176.950 ;
        RECT 22.010 -177.120 22.330 -177.090 ;
        RECT 24.690 -176.950 25.010 -176.840 ;
        RECT 25.350 -176.950 25.510 -176.160 ;
        RECT 26.950 -176.310 27.290 -176.160 ;
        RECT 26.970 -176.510 27.290 -176.480 ;
        RECT 24.690 -177.090 25.510 -176.950 ;
        RECT 26.470 -176.650 27.290 -176.510 ;
        RECT 24.690 -177.120 25.010 -177.090 ;
        RECT 21.990 -177.440 22.330 -177.290 ;
        RECT 20.390 -177.590 22.330 -177.440 ;
        RECT 24.690 -177.440 25.030 -177.290 ;
        RECT 26.470 -177.440 26.630 -176.650 ;
        RECT 26.970 -176.760 27.290 -176.650 ;
        RECT 24.690 -177.590 26.630 -177.440 ;
        RECT -289.200 -178.400 -287.360 -177.920 ;
        RECT -287.440 -179.490 -286.960 -178.590 ;
        RECT -286.140 -178.720 -285.950 -177.590 ;
        RECT -282.070 -178.720 -281.880 -177.590 ;
        RECT -276.220 -178.720 -276.030 -177.590 ;
        RECT -272.150 -178.720 -271.960 -177.590 ;
        RECT -266.300 -178.720 -266.110 -177.590 ;
        RECT -262.230 -178.720 -262.040 -177.590 ;
        RECT -256.380 -178.720 -256.190 -177.590 ;
        RECT -252.310 -178.720 -252.120 -177.590 ;
        RECT -246.460 -178.720 -246.270 -177.590 ;
        RECT -242.390 -178.720 -242.200 -177.590 ;
        RECT -236.540 -178.720 -236.350 -177.590 ;
        RECT -232.470 -178.720 -232.280 -177.590 ;
        RECT -226.620 -178.720 -226.430 -177.590 ;
        RECT -222.550 -178.720 -222.360 -177.590 ;
        RECT -216.700 -178.720 -216.510 -177.590 ;
        RECT -212.630 -178.720 -212.440 -177.590 ;
        RECT -206.780 -178.720 -206.590 -177.590 ;
        RECT -202.710 -178.720 -202.520 -177.590 ;
        RECT -196.860 -178.720 -196.670 -177.590 ;
        RECT -192.790 -178.720 -192.600 -177.590 ;
        RECT -186.940 -178.720 -186.750 -177.590 ;
        RECT -182.870 -178.720 -182.680 -177.590 ;
        RECT -177.020 -178.720 -176.830 -177.590 ;
        RECT -172.950 -178.720 -172.760 -177.590 ;
        RECT -167.100 -178.720 -166.910 -177.590 ;
        RECT -163.030 -178.720 -162.840 -177.590 ;
        RECT -157.180 -178.720 -156.990 -177.590 ;
        RECT -153.110 -178.720 -152.920 -177.590 ;
        RECT -147.260 -178.720 -147.070 -177.590 ;
        RECT -143.190 -178.720 -143.000 -177.590 ;
        RECT -137.340 -178.720 -137.150 -177.590 ;
        RECT -133.270 -178.720 -133.080 -177.590 ;
        RECT -127.420 -178.720 -127.230 -177.590 ;
        RECT -123.350 -178.720 -123.160 -177.590 ;
        RECT -117.500 -178.720 -117.310 -177.590 ;
        RECT -113.430 -178.720 -113.240 -177.590 ;
        RECT -107.580 -178.720 -107.390 -177.590 ;
        RECT -103.510 -178.720 -103.320 -177.590 ;
        RECT -97.660 -178.720 -97.470 -177.590 ;
        RECT -93.590 -178.720 -93.400 -177.590 ;
        RECT -87.740 -178.720 -87.550 -177.590 ;
        RECT -83.670 -178.720 -83.480 -177.590 ;
        RECT -77.820 -178.720 -77.630 -177.590 ;
        RECT -73.750 -178.720 -73.560 -177.590 ;
        RECT -67.900 -178.720 -67.710 -177.590 ;
        RECT -63.830 -178.720 -63.640 -177.590 ;
        RECT -57.980 -178.720 -57.790 -177.590 ;
        RECT -53.910 -178.720 -53.720 -177.590 ;
        RECT -48.060 -178.720 -47.870 -177.590 ;
        RECT -43.990 -178.720 -43.800 -177.590 ;
        RECT -38.140 -178.720 -37.950 -177.590 ;
        RECT -34.070 -178.720 -33.880 -177.590 ;
        RECT -28.220 -178.720 -28.030 -177.590 ;
        RECT -24.150 -178.720 -23.960 -177.590 ;
        RECT -18.300 -178.720 -18.110 -177.590 ;
        RECT -14.230 -178.720 -14.040 -177.590 ;
        RECT -8.380 -178.720 -8.190 -177.590 ;
        RECT -4.310 -178.720 -4.120 -177.590 ;
        RECT 1.540 -178.720 1.730 -177.590 ;
        RECT 5.610 -178.720 5.800 -177.590 ;
        RECT 11.460 -178.720 11.650 -177.590 ;
        RECT 15.530 -178.720 15.720 -177.590 ;
        RECT 21.380 -178.720 21.570 -177.590 ;
        RECT 25.450 -178.720 25.640 -177.590 ;
        RECT -286.190 -179.010 -285.870 -178.720 ;
        RECT -282.150 -179.010 -281.830 -178.720 ;
        RECT -276.270 -179.010 -275.950 -178.720 ;
        RECT -272.230 -179.010 -271.910 -178.720 ;
        RECT -266.350 -179.010 -266.030 -178.720 ;
        RECT -262.310 -179.010 -261.990 -178.720 ;
        RECT -256.430 -179.010 -256.110 -178.720 ;
        RECT -252.390 -179.010 -252.070 -178.720 ;
        RECT -246.510 -179.010 -246.190 -178.720 ;
        RECT -242.470 -179.010 -242.150 -178.720 ;
        RECT -236.590 -179.010 -236.270 -178.720 ;
        RECT -232.550 -179.010 -232.230 -178.720 ;
        RECT -226.670 -179.010 -226.350 -178.720 ;
        RECT -222.630 -179.010 -222.310 -178.720 ;
        RECT -216.750 -179.010 -216.430 -178.720 ;
        RECT -212.710 -179.010 -212.390 -178.720 ;
        RECT -206.830 -179.010 -206.510 -178.720 ;
        RECT -202.790 -179.010 -202.470 -178.720 ;
        RECT -196.910 -179.010 -196.590 -178.720 ;
        RECT -192.870 -179.010 -192.550 -178.720 ;
        RECT -186.990 -179.010 -186.670 -178.720 ;
        RECT -182.950 -179.010 -182.630 -178.720 ;
        RECT -177.070 -179.010 -176.750 -178.720 ;
        RECT -173.030 -179.010 -172.710 -178.720 ;
        RECT -167.150 -179.010 -166.830 -178.720 ;
        RECT -163.110 -179.010 -162.790 -178.720 ;
        RECT -157.230 -179.010 -156.910 -178.720 ;
        RECT -153.190 -179.010 -152.870 -178.720 ;
        RECT -147.310 -179.010 -146.990 -178.720 ;
        RECT -143.270 -179.010 -142.950 -178.720 ;
        RECT -137.390 -179.010 -137.070 -178.720 ;
        RECT -133.350 -179.010 -133.030 -178.720 ;
        RECT -127.470 -179.010 -127.150 -178.720 ;
        RECT -123.430 -179.010 -123.110 -178.720 ;
        RECT -117.550 -179.010 -117.230 -178.720 ;
        RECT -113.510 -179.010 -113.190 -178.720 ;
        RECT -107.630 -179.010 -107.310 -178.720 ;
        RECT -103.590 -179.010 -103.270 -178.720 ;
        RECT -97.710 -179.010 -97.390 -178.720 ;
        RECT -93.670 -179.010 -93.350 -178.720 ;
        RECT -87.790 -179.010 -87.470 -178.720 ;
        RECT -83.750 -179.010 -83.430 -178.720 ;
        RECT -77.870 -179.010 -77.550 -178.720 ;
        RECT -73.830 -179.010 -73.510 -178.720 ;
        RECT -67.950 -179.010 -67.630 -178.720 ;
        RECT -63.910 -179.010 -63.590 -178.720 ;
        RECT -58.030 -179.010 -57.710 -178.720 ;
        RECT -53.990 -179.010 -53.670 -178.720 ;
        RECT -48.110 -179.010 -47.790 -178.720 ;
        RECT -44.070 -179.010 -43.750 -178.720 ;
        RECT -38.190 -179.010 -37.870 -178.720 ;
        RECT -34.150 -179.010 -33.830 -178.720 ;
        RECT -28.270 -179.010 -27.950 -178.720 ;
        RECT -24.230 -179.010 -23.910 -178.720 ;
        RECT -18.350 -179.010 -18.030 -178.720 ;
        RECT -14.310 -179.010 -13.990 -178.720 ;
        RECT -8.430 -179.010 -8.110 -178.720 ;
        RECT -4.390 -179.010 -4.070 -178.720 ;
        RECT 1.490 -179.010 1.810 -178.720 ;
        RECT 5.530 -179.010 5.850 -178.720 ;
        RECT 11.410 -179.010 11.730 -178.720 ;
        RECT 15.450 -179.010 15.770 -178.720 ;
        RECT 21.330 -179.010 21.650 -178.720 ;
        RECT 25.370 -179.010 25.690 -178.720 ;
        RECT -287.900 -179.970 -286.960 -179.490 ;
        RECT 26.460 -179.490 26.940 -178.590 ;
        RECT -282.890 -179.890 -281.200 -179.590 ;
        RECT -272.970 -179.890 -271.280 -179.590 ;
        RECT -263.050 -179.890 -261.360 -179.590 ;
        RECT -253.130 -179.890 -251.440 -179.590 ;
        RECT -243.210 -179.890 -241.520 -179.590 ;
        RECT -233.290 -179.890 -231.600 -179.590 ;
        RECT -223.370 -179.890 -221.680 -179.590 ;
        RECT -213.450 -179.890 -211.760 -179.590 ;
        RECT -203.530 -179.890 -201.840 -179.590 ;
        RECT -193.610 -179.890 -191.920 -179.590 ;
        RECT -183.690 -179.890 -182.000 -179.590 ;
        RECT -173.770 -179.890 -172.080 -179.590 ;
        RECT -163.850 -179.890 -162.160 -179.590 ;
        RECT -153.930 -179.890 -152.240 -179.590 ;
        RECT -144.010 -179.890 -142.320 -179.590 ;
        RECT -134.090 -179.890 -132.400 -179.590 ;
        RECT -124.170 -179.890 -122.480 -179.590 ;
        RECT -114.250 -179.890 -112.560 -179.590 ;
        RECT -104.330 -179.890 -102.640 -179.590 ;
        RECT -94.410 -179.890 -92.720 -179.590 ;
        RECT -84.490 -179.890 -82.800 -179.590 ;
        RECT -74.570 -179.890 -72.880 -179.590 ;
        RECT -64.650 -179.890 -62.960 -179.590 ;
        RECT -54.730 -179.890 -53.040 -179.590 ;
        RECT -44.810 -179.890 -43.120 -179.590 ;
        RECT -34.890 -179.890 -33.200 -179.590 ;
        RECT -24.970 -179.890 -23.280 -179.590 ;
        RECT -15.050 -179.890 -13.360 -179.590 ;
        RECT -5.130 -179.890 -3.440 -179.590 ;
        RECT 4.790 -179.890 6.480 -179.590 ;
        RECT 14.710 -179.890 16.400 -179.590 ;
        RECT 24.630 -179.890 26.320 -179.590 ;
        RECT -282.380 -180.590 -281.380 -179.890 ;
        RECT -272.460 -180.590 -271.460 -179.890 ;
        RECT -262.540 -180.590 -261.540 -179.890 ;
        RECT -252.620 -180.590 -251.620 -179.890 ;
        RECT -242.700 -180.590 -241.700 -179.890 ;
        RECT -232.780 -180.590 -231.780 -179.890 ;
        RECT -222.860 -180.590 -221.860 -179.890 ;
        RECT -212.940 -180.590 -211.940 -179.890 ;
        RECT -203.020 -180.590 -202.020 -179.890 ;
        RECT -193.100 -180.590 -192.100 -179.890 ;
        RECT -183.180 -180.590 -182.180 -179.890 ;
        RECT -173.260 -180.590 -172.260 -179.890 ;
        RECT -163.340 -180.590 -162.340 -179.890 ;
        RECT -153.420 -180.590 -152.420 -179.890 ;
        RECT -143.500 -180.590 -142.500 -179.890 ;
        RECT -133.580 -180.590 -132.580 -179.890 ;
        RECT -123.660 -180.590 -122.660 -179.890 ;
        RECT -113.740 -180.590 -112.740 -179.890 ;
        RECT -103.820 -180.590 -102.820 -179.890 ;
        RECT -93.900 -180.590 -92.900 -179.890 ;
        RECT -83.980 -180.590 -82.980 -179.890 ;
        RECT -74.060 -180.590 -73.060 -179.890 ;
        RECT -64.140 -180.590 -63.140 -179.890 ;
        RECT -54.220 -180.590 -53.220 -179.890 ;
        RECT -44.300 -180.590 -43.300 -179.890 ;
        RECT -34.380 -180.590 -33.380 -179.890 ;
        RECT -24.460 -180.590 -23.460 -179.890 ;
        RECT -14.540 -180.590 -13.540 -179.890 ;
        RECT -4.620 -180.590 -3.620 -179.890 ;
        RECT 5.300 -180.590 6.300 -179.890 ;
        RECT 15.220 -180.590 16.220 -179.890 ;
        RECT 25.140 -180.590 26.140 -179.890 ;
        RECT 26.460 -179.970 27.400 -179.490 ;
  END
END meta_srlatch_set
END LIBRARY

