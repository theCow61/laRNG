VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO meta_srlatch_singleready_flat
  CLASS BLOCK ;
  FOREIGN meta_srlatch_singleready_flat ;
  ORIGIN 1.860 0.250 ;
  SIZE 5.800 BY 7.640 ;
  SITE unithd ;
  PIN i_srclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.860 3.605 3.195 3.875 ;
        RECT -1.115 3.265 -0.780 3.535 ;
      LAYER mcon ;
        RECT 2.940 3.685 3.110 3.855 ;
        RECT -1.030 3.285 -0.860 3.455 ;
      LAYER met1 ;
        RECT -1.220 3.190 -0.760 3.640 ;
        RECT 2.840 3.500 3.300 3.950 ;
      LAYER via ;
        RECT -1.150 3.240 -0.850 3.540 ;
        RECT 2.930 3.600 3.230 3.900 ;
      LAYER met2 ;
        RECT 0.970 3.640 1.110 4.040 ;
        RECT 2.840 3.640 3.300 3.950 ;
        RECT -1.220 3.500 3.300 3.640 ;
        RECT -1.220 3.190 -0.760 3.500 ;
        RECT 0.970 3.100 1.110 3.500 ;
    END
  END i_srclk
  PIN o_ranQ
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 0.585 6.475 2.795 6.655 ;
        RECT 0.585 6.395 1.090 6.475 ;
        RECT 1.890 6.385 2.795 6.475 ;
      LAYER mcon ;
        RECT 0.775 6.395 0.945 6.565 ;
        RECT 2.140 6.395 2.310 6.565 ;
      LAYER met1 ;
        RECT 0.890 6.660 1.890 7.360 ;
        RECT 0.710 6.360 2.400 6.660 ;
    END
  END o_ranQ
  PIN o_ranNQ
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -0.715 0.665 0.190 0.755 ;
        RECT 0.990 0.665 1.495 0.745 ;
        RECT -0.715 0.485 1.495 0.665 ;
      LAYER mcon ;
        RECT -0.230 0.575 -0.060 0.745 ;
        RECT 1.135 0.575 1.305 0.745 ;
      LAYER met1 ;
        RECT -0.320 0.480 1.370 0.780 ;
        RECT 0.190 -0.220 1.190 0.480 ;
    END
  END o_ranNQ
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 1.635 5.170 3.240 7.390 ;
        RECT -1.860 3.515 0.360 5.120 ;
        RECT 1.720 2.020 3.940 3.625 ;
        RECT -1.160 -0.250 0.445 1.970 ;
      LAYER li1 ;
        RECT 2.965 7.115 3.135 7.200 ;
        RECT 1.800 6.825 3.135 7.115 ;
        RECT 2.965 6.215 3.135 6.825 ;
        RECT 2.205 5.885 3.135 6.215 ;
        RECT 2.965 5.360 3.135 5.885 ;
        RECT -1.670 4.845 0.170 5.015 ;
        RECT -1.585 3.680 -1.295 4.845 ;
        RECT -1.125 3.705 -0.845 4.845 ;
        RECT -0.175 3.705 0.085 4.845 ;
        RECT 1.995 2.295 2.255 3.435 ;
        RECT 2.925 2.295 3.205 3.435 ;
        RECT 3.375 2.295 3.665 3.460 ;
        RECT 1.910 2.125 3.750 2.295 ;
        RECT -1.055 1.255 -0.885 1.780 ;
        RECT -1.055 0.925 -0.125 1.255 ;
        RECT -1.055 0.315 -0.885 0.925 ;
        RECT -1.055 0.025 0.280 0.315 ;
        RECT -1.055 -0.060 -0.885 0.025 ;
      LAYER mcon ;
        RECT 2.965 6.885 3.135 7.055 ;
        RECT 2.965 6.425 3.135 6.595 ;
        RECT 2.965 5.965 3.135 6.135 ;
        RECT 2.965 5.505 3.135 5.675 ;
        RECT -1.525 4.845 -1.355 5.015 ;
        RECT -1.065 4.845 -0.895 5.015 ;
        RECT -0.605 4.845 -0.435 5.015 ;
        RECT -0.145 4.845 0.025 5.015 ;
        RECT 2.055 2.125 2.225 2.295 ;
        RECT 2.515 2.125 2.685 2.295 ;
        RECT 2.975 2.125 3.145 2.295 ;
        RECT 3.435 2.125 3.605 2.295 ;
        RECT -1.055 1.465 -0.885 1.635 ;
        RECT -1.055 1.005 -0.885 1.175 ;
        RECT -1.055 0.545 -0.885 0.715 ;
        RECT -1.055 0.085 -0.885 0.255 ;
      LAYER met1 ;
        RECT 2.810 5.360 3.290 7.200 ;
        RECT -1.670 4.690 0.170 5.170 ;
        RECT 1.910 1.970 3.750 2.450 ;
        RECT -1.210 -0.060 -0.730 1.780 ;
      LAYER via ;
        RECT 2.900 6.820 3.200 7.110 ;
        RECT 2.900 5.870 3.200 6.160 ;
        RECT -1.550 4.770 -1.250 5.060 ;
        RECT -0.640 4.810 -0.340 5.100 ;
        RECT 2.440 2.070 2.740 2.360 ;
        RECT 3.340 2.050 3.640 2.340 ;
        RECT -1.160 1.200 -0.860 1.490 ;
        RECT -1.160 0.540 -0.860 0.830 ;
      LAYER met2 ;
        RECT 2.810 5.360 3.290 7.200 ;
        RECT -1.670 4.690 0.160 5.170 ;
        RECT 1.910 1.970 3.750 2.450 ;
        RECT -1.210 -0.060 -0.730 1.780 ;
      LAYER via2 ;
        RECT 2.900 6.820 3.200 7.110 ;
        RECT 2.900 5.870 3.200 6.160 ;
        RECT -1.550 4.770 -1.250 5.060 ;
        RECT -0.640 4.810 -0.340 5.100 ;
        RECT 2.440 2.070 2.740 2.360 ;
        RECT 3.340 2.050 3.640 2.340 ;
        RECT -1.160 1.200 -0.860 1.490 ;
        RECT -1.160 0.540 -0.860 0.830 ;
      LAYER met3 ;
        RECT -1.670 4.690 0.160 5.170 ;
        RECT -1.210 3.870 -0.730 4.690 ;
        RECT 2.810 3.870 3.290 7.200 ;
        RECT -1.220 3.280 3.300 3.870 ;
        RECT -1.210 -0.060 -0.730 3.280 ;
        RECT 2.810 2.450 3.290 3.280 ;
        RECT 1.910 1.970 3.750 2.450 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.520 7.180 1.305 7.185 ;
        RECT 0.440 6.755 1.305 7.180 ;
        RECT 0.440 6.735 1.210 6.755 ;
        RECT 0.435 5.685 1.215 6.735 ;
        RECT 0.245 5.515 1.215 5.685 ;
        RECT 0.435 5.365 1.215 5.515 ;
        RECT 2.980 4.825 3.150 5.015 ;
        RECT 1.915 4.740 3.265 4.825 ;
        RECT 1.915 3.960 3.740 4.740 ;
        RECT 1.915 3.915 3.265 3.960 ;
        RECT 3.305 3.955 3.735 3.960 ;
        RECT -1.655 3.180 -1.225 3.185 ;
        RECT -1.185 3.180 0.165 3.225 ;
        RECT -1.655 2.400 0.165 3.180 ;
        RECT -1.185 2.315 0.165 2.400 ;
        RECT -1.070 2.125 -0.900 2.315 ;
        RECT 0.865 1.625 1.645 1.775 ;
        RECT 0.865 1.455 1.835 1.625 ;
        RECT 0.865 0.405 1.645 1.455 ;
        RECT 0.870 0.385 1.640 0.405 ;
        RECT 0.775 -0.040 1.640 0.385 ;
        RECT 0.775 -0.045 1.560 -0.040 ;
      LAYER li1 ;
        RECT 0.245 7.115 0.415 7.200 ;
        RECT 0.245 6.825 1.140 7.115 ;
        RECT 0.245 6.215 0.415 6.825 ;
        RECT 0.245 5.885 0.795 6.215 ;
        RECT 0.245 5.360 0.415 5.885 ;
        RECT 1.910 4.845 3.750 5.015 ;
        RECT 2.895 4.045 3.205 4.845 ;
        RECT 3.375 4.120 3.665 4.845 ;
        RECT -1.585 2.295 -1.295 3.020 ;
        RECT -1.125 2.295 -0.815 3.095 ;
        RECT -1.670 2.125 0.170 2.295 ;
        RECT 1.665 1.255 1.835 1.780 ;
        RECT 1.285 0.925 1.835 1.255 ;
        RECT 1.665 0.315 1.835 0.925 ;
        RECT 0.940 0.025 1.835 0.315 ;
        RECT 1.665 -0.060 1.835 0.025 ;
      LAYER mcon ;
        RECT 0.245 6.885 0.415 7.055 ;
        RECT 0.245 6.425 0.415 6.595 ;
        RECT 0.245 5.965 0.415 6.135 ;
        RECT 0.245 5.505 0.415 5.675 ;
        RECT 2.055 4.845 2.225 5.015 ;
        RECT 2.515 4.845 2.685 5.015 ;
        RECT 2.975 4.845 3.145 5.015 ;
        RECT 3.435 4.845 3.605 5.015 ;
        RECT -1.525 2.125 -1.355 2.295 ;
        RECT -1.065 2.125 -0.895 2.295 ;
        RECT -0.605 2.125 -0.435 2.295 ;
        RECT -0.145 2.125 0.025 2.295 ;
        RECT 1.665 1.465 1.835 1.635 ;
        RECT 1.665 1.005 1.835 1.175 ;
        RECT 1.665 0.545 1.835 0.715 ;
        RECT 1.665 0.085 1.835 0.255 ;
      LAYER met1 ;
        RECT 0.090 5.360 0.570 7.200 ;
        RECT 1.910 4.690 3.750 5.170 ;
        RECT -1.670 1.970 0.170 2.450 ;
        RECT 1.510 -0.060 1.990 1.780 ;
      LAYER via ;
        RECT 0.190 5.890 0.490 6.180 ;
        RECT 2.010 4.790 2.310 5.080 ;
        RECT -0.220 2.060 0.080 2.350 ;
        RECT 1.620 0.940 1.920 1.230 ;
      LAYER met2 ;
        RECT 0.080 5.370 0.570 7.200 ;
        RECT 1.910 4.680 3.760 5.160 ;
        RECT -1.670 1.980 0.170 2.440 ;
        RECT 1.500 -0.080 1.990 1.780 ;
      LAYER via2 ;
        RECT 0.190 5.890 0.490 6.180 ;
        RECT 2.010 4.790 2.310 5.080 ;
        RECT -0.260 2.030 0.140 2.380 ;
        RECT 1.620 0.940 1.920 1.230 ;
      LAYER met3 ;
        RECT 0.080 5.490 0.530 7.190 ;
        RECT 1.530 4.700 2.430 5.150 ;
        RECT -0.320 1.970 0.380 2.440 ;
        RECT 1.510 1.550 2.000 1.570 ;
        RECT 1.500 -0.070 2.000 1.550 ;
        RECT 1.500 -0.090 1.990 -0.070 ;
      LAYER via3 ;
        RECT 0.120 5.850 0.520 6.200 ;
        RECT 1.960 4.760 2.360 5.110 ;
        RECT -0.260 2.030 0.140 2.380 ;
        RECT 1.570 0.910 1.970 1.260 ;
      LAYER met4 ;
        RECT 0.080 5.370 0.570 7.200 ;
        RECT 0.090 5.160 0.570 5.370 ;
        RECT 1.500 5.160 3.750 5.170 ;
        RECT 0.090 4.680 3.760 5.160 ;
        RECT 0.090 2.450 0.570 4.680 ;
        RECT 1.500 2.450 1.990 4.680 ;
        RECT -1.670 1.970 2.000 2.450 ;
        RECT 1.500 -0.080 1.990 1.970 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.390 6.200 1.720 6.305 ;
        RECT 0.965 6.030 2.035 6.200 ;
        RECT 0.965 5.705 1.135 6.030 ;
        RECT 0.585 5.535 1.135 5.705 ;
        RECT 1.315 5.465 1.685 5.805 ;
        RECT 1.865 5.705 2.035 6.030 ;
        RECT 1.865 5.525 2.795 5.705 ;
        RECT -0.675 3.695 -0.345 4.675 ;
        RECT 1.995 4.045 2.690 4.675 ;
        RECT -0.610 3.095 -0.440 3.695 ;
        RECT 2.015 3.605 2.350 3.855 ;
        RECT -0.270 3.285 0.065 3.535 ;
        RECT 2.520 3.445 2.690 4.045 ;
        RECT -0.610 2.465 0.085 3.095 ;
        RECT 2.425 2.465 2.755 3.445 ;
        RECT -0.715 1.435 0.215 1.615 ;
        RECT 0.045 1.110 0.215 1.435 ;
        RECT 0.395 1.335 0.765 1.675 ;
        RECT 0.945 1.435 1.495 1.605 ;
        RECT 0.945 1.110 1.115 1.435 ;
        RECT 0.045 0.940 1.115 1.110 ;
        RECT 0.360 0.835 0.690 0.940 ;
      LAYER mcon ;
        RECT 1.405 5.545 1.575 5.715 ;
        RECT 2.085 4.125 2.255 4.295 ;
        RECT 2.100 3.685 2.270 3.855 ;
        RECT -0.190 3.285 -0.020 3.455 ;
        RECT -0.175 2.845 -0.005 3.015 ;
        RECT 0.505 1.425 0.675 1.595 ;
      LAYER met1 ;
        RECT 1.340 5.490 1.660 5.780 ;
        RECT 1.390 4.360 1.580 5.490 ;
        RECT 0.400 4.210 2.340 4.360 ;
        RECT -0.260 3.420 0.060 3.530 ;
        RECT 0.400 3.420 0.560 4.210 ;
        RECT 2.000 4.060 2.340 4.210 ;
        RECT 2.020 3.860 2.340 3.890 ;
        RECT -0.260 3.280 0.560 3.420 ;
        RECT 1.520 3.720 2.340 3.860 ;
        RECT -0.260 3.250 0.060 3.280 ;
        RECT -0.260 2.930 0.080 3.080 ;
        RECT 1.520 2.930 1.680 3.720 ;
        RECT 2.020 3.610 2.340 3.720 ;
        RECT -0.260 2.780 1.680 2.930 ;
        RECT 0.500 1.650 0.690 2.780 ;
        RECT 0.420 1.360 0.740 1.650 ;
  END
END meta_srlatch_singleready_flat
END LIBRARY

