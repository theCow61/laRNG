VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO meta_srlatch_stack
  CLASS BLOCK ;
  FOREIGN meta_srlatch_stack ;
  ORIGIN 339.920 194.560 ;
  SIZE 504.270 BY 304.430 ;
  SITE unithd ;
  PIN o_ranQ[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 18.315 89.065 18.820 89.145 ;
        RECT 19.620 89.065 20.525 89.155 ;
        RECT 18.315 88.885 20.525 89.065 ;
      LAYER mcon ;
        RECT 18.505 88.975 18.675 89.145 ;
        RECT 19.870 88.975 20.040 89.145 ;
      LAYER met1 ;
        RECT 18.440 88.880 20.130 89.180 ;
        RECT 18.620 88.180 19.620 88.880 ;
    END
  END o_ranQ[1]
  PIN o_ranQ[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 13.355 94.875 15.565 95.055 ;
        RECT 13.355 94.795 13.860 94.875 ;
        RECT 14.660 94.785 15.565 94.875 ;
      LAYER mcon ;
        RECT 13.545 94.795 13.715 94.965 ;
        RECT 14.910 94.795 15.080 94.965 ;
      LAYER met1 ;
        RECT 13.660 95.060 14.660 95.760 ;
        RECT 13.480 94.760 15.170 95.060 ;
    END
  END o_ranQ[2]
  PIN o_ranQ[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 8.395 89.065 8.900 89.145 ;
        RECT 9.700 89.065 10.605 89.155 ;
        RECT 8.395 88.885 10.605 89.065 ;
      LAYER mcon ;
        RECT 8.585 88.975 8.755 89.145 ;
        RECT 9.950 88.975 10.120 89.145 ;
      LAYER met1 ;
        RECT 8.520 88.880 10.210 89.180 ;
        RECT 8.700 88.180 9.700 88.880 ;
    END
  END o_ranQ[3]
  PIN o_ranQ[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 23.275 94.875 25.485 95.055 ;
        RECT 23.275 94.795 23.780 94.875 ;
        RECT 24.580 94.785 25.485 94.875 ;
      LAYER mcon ;
        RECT 23.465 94.795 23.635 94.965 ;
        RECT 24.830 94.795 25.000 94.965 ;
      LAYER met1 ;
        RECT 23.580 95.060 24.580 95.760 ;
        RECT 23.400 94.760 25.090 95.060 ;
    END
  END o_ranQ[0]
  PIN o_ranQ[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 3.435 94.875 5.645 95.055 ;
        RECT 3.435 94.795 3.940 94.875 ;
        RECT 4.740 94.785 5.645 94.875 ;
      LAYER mcon ;
        RECT 3.625 94.795 3.795 94.965 ;
        RECT 4.990 94.795 5.160 94.965 ;
      LAYER met1 ;
        RECT 3.740 95.060 4.740 95.760 ;
        RECT 3.560 94.760 5.250 95.060 ;
    END
  END o_ranQ[4]
  PIN o_ranQ[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -1.525 89.065 -1.020 89.145 ;
        RECT -0.220 89.065 0.685 89.155 ;
        RECT -1.525 88.885 0.685 89.065 ;
      LAYER mcon ;
        RECT -1.335 88.975 -1.165 89.145 ;
        RECT 0.030 88.975 0.200 89.145 ;
      LAYER met1 ;
        RECT -1.400 88.880 0.290 89.180 ;
        RECT -1.220 88.180 -0.220 88.880 ;
    END
  END o_ranQ[5]
  PIN o_ranQ[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -6.485 94.875 -4.275 95.055 ;
        RECT -6.485 94.795 -5.980 94.875 ;
        RECT -5.180 94.785 -4.275 94.875 ;
      LAYER mcon ;
        RECT -6.295 94.795 -6.125 94.965 ;
        RECT -4.930 94.795 -4.760 94.965 ;
      LAYER met1 ;
        RECT -6.180 95.060 -5.180 95.760 ;
        RECT -6.360 94.760 -4.670 95.060 ;
    END
  END o_ranQ[6]
  PIN o_ranQ[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -11.445 89.065 -10.940 89.145 ;
        RECT -10.140 89.065 -9.235 89.155 ;
        RECT -11.445 88.885 -9.235 89.065 ;
      LAYER mcon ;
        RECT -11.255 88.975 -11.085 89.145 ;
        RECT -9.890 88.975 -9.720 89.145 ;
      LAYER met1 ;
        RECT -11.320 88.880 -9.630 89.180 ;
        RECT -11.140 88.180 -10.140 88.880 ;
    END
  END o_ranQ[7]
  PIN o_ranQ[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -16.405 94.875 -14.195 95.055 ;
        RECT -16.405 94.795 -15.900 94.875 ;
        RECT -15.100 94.785 -14.195 94.875 ;
      LAYER mcon ;
        RECT -16.215 94.795 -16.045 94.965 ;
        RECT -14.850 94.795 -14.680 94.965 ;
      LAYER met1 ;
        RECT -16.100 95.060 -15.100 95.760 ;
        RECT -16.280 94.760 -14.590 95.060 ;
    END
  END o_ranQ[8]
  PIN o_ranQ[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -21.365 89.065 -20.860 89.145 ;
        RECT -20.060 89.065 -19.155 89.155 ;
        RECT -21.365 88.885 -19.155 89.065 ;
      LAYER mcon ;
        RECT -21.175 88.975 -21.005 89.145 ;
        RECT -19.810 88.975 -19.640 89.145 ;
      LAYER met1 ;
        RECT -21.240 88.880 -19.550 89.180 ;
        RECT -21.060 88.180 -20.060 88.880 ;
    END
  END o_ranQ[9]
  PIN o_ranQ[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -26.325 94.875 -24.115 95.055 ;
        RECT -26.325 94.795 -25.820 94.875 ;
        RECT -25.020 94.785 -24.115 94.875 ;
      LAYER mcon ;
        RECT -26.135 94.795 -25.965 94.965 ;
        RECT -24.770 94.795 -24.600 94.965 ;
      LAYER met1 ;
        RECT -26.020 95.060 -25.020 95.760 ;
        RECT -26.200 94.760 -24.510 95.060 ;
    END
  END o_ranQ[10]
  PIN o_ranQ[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -31.285 89.065 -30.780 89.145 ;
        RECT -29.980 89.065 -29.075 89.155 ;
        RECT -31.285 88.885 -29.075 89.065 ;
      LAYER mcon ;
        RECT -31.095 88.975 -30.925 89.145 ;
        RECT -29.730 88.975 -29.560 89.145 ;
      LAYER met1 ;
        RECT -31.160 88.880 -29.470 89.180 ;
        RECT -30.980 88.180 -29.980 88.880 ;
    END
  END o_ranQ[11]
  PIN o_ranQ[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -36.245 94.875 -34.035 95.055 ;
        RECT -36.245 94.795 -35.740 94.875 ;
        RECT -34.940 94.785 -34.035 94.875 ;
      LAYER mcon ;
        RECT -36.055 94.795 -35.885 94.965 ;
        RECT -34.690 94.795 -34.520 94.965 ;
      LAYER met1 ;
        RECT -35.940 95.060 -34.940 95.760 ;
        RECT -36.120 94.760 -34.430 95.060 ;
    END
  END o_ranQ[12]
  PIN o_ranQ[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -41.205 89.065 -40.700 89.145 ;
        RECT -39.900 89.065 -38.995 89.155 ;
        RECT -41.205 88.885 -38.995 89.065 ;
      LAYER mcon ;
        RECT -41.015 88.975 -40.845 89.145 ;
        RECT -39.650 88.975 -39.480 89.145 ;
      LAYER met1 ;
        RECT -41.080 88.880 -39.390 89.180 ;
        RECT -40.900 88.180 -39.900 88.880 ;
    END
  END o_ranQ[13]
  PIN o_ranQ[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -46.165 94.875 -43.955 95.055 ;
        RECT -46.165 94.795 -45.660 94.875 ;
        RECT -44.860 94.785 -43.955 94.875 ;
      LAYER mcon ;
        RECT -45.975 94.795 -45.805 94.965 ;
        RECT -44.610 94.795 -44.440 94.965 ;
      LAYER met1 ;
        RECT -45.860 95.060 -44.860 95.760 ;
        RECT -46.040 94.760 -44.350 95.060 ;
    END
  END o_ranQ[14]
  PIN o_ranQ[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -51.125 89.065 -50.620 89.145 ;
        RECT -49.820 89.065 -48.915 89.155 ;
        RECT -51.125 88.885 -48.915 89.065 ;
      LAYER mcon ;
        RECT -50.935 88.975 -50.765 89.145 ;
        RECT -49.570 88.975 -49.400 89.145 ;
      LAYER met1 ;
        RECT -51.000 88.880 -49.310 89.180 ;
        RECT -50.820 88.180 -49.820 88.880 ;
    END
  END o_ranQ[15]
  PIN o_ranQ[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -61.045 89.065 -60.540 89.145 ;
        RECT -59.740 89.065 -58.835 89.155 ;
        RECT -61.045 88.885 -58.835 89.065 ;
      LAYER mcon ;
        RECT -60.855 88.975 -60.685 89.145 ;
        RECT -59.490 88.975 -59.320 89.145 ;
      LAYER met1 ;
        RECT -60.920 88.880 -59.230 89.180 ;
        RECT -60.740 88.180 -59.740 88.880 ;
    END
  END o_ranQ[17]
  PIN o_ranQ[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -66.005 94.875 -63.795 95.055 ;
        RECT -66.005 94.795 -65.500 94.875 ;
        RECT -64.700 94.785 -63.795 94.875 ;
      LAYER mcon ;
        RECT -65.815 94.795 -65.645 94.965 ;
        RECT -64.450 94.795 -64.280 94.965 ;
      LAYER met1 ;
        RECT -65.700 95.060 -64.700 95.760 ;
        RECT -65.880 94.760 -64.190 95.060 ;
    END
  END o_ranQ[18]
  PIN o_ranQ[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -70.965 89.065 -70.460 89.145 ;
        RECT -69.660 89.065 -68.755 89.155 ;
        RECT -70.965 88.885 -68.755 89.065 ;
      LAYER mcon ;
        RECT -70.775 88.975 -70.605 89.145 ;
        RECT -69.410 88.975 -69.240 89.145 ;
      LAYER met1 ;
        RECT -70.840 88.880 -69.150 89.180 ;
        RECT -70.660 88.180 -69.660 88.880 ;
    END
  END o_ranQ[19]
  PIN o_ranQ[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -56.085 94.875 -53.875 95.055 ;
        RECT -56.085 94.795 -55.580 94.875 ;
        RECT -54.780 94.785 -53.875 94.875 ;
      LAYER mcon ;
        RECT -55.895 94.795 -55.725 94.965 ;
        RECT -54.530 94.795 -54.360 94.965 ;
      LAYER met1 ;
        RECT -55.780 95.060 -54.780 95.760 ;
        RECT -55.960 94.760 -54.270 95.060 ;
    END
  END o_ranQ[16]
  PIN o_ranQ[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -75.925 94.875 -73.715 95.055 ;
        RECT -75.925 94.795 -75.420 94.875 ;
        RECT -74.620 94.785 -73.715 94.875 ;
      LAYER mcon ;
        RECT -75.735 94.795 -75.565 94.965 ;
        RECT -74.370 94.795 -74.200 94.965 ;
      LAYER met1 ;
        RECT -75.620 95.060 -74.620 95.760 ;
        RECT -75.800 94.760 -74.110 95.060 ;
    END
  END o_ranQ[20]
  PIN o_ranQ[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -80.885 89.065 -80.380 89.145 ;
        RECT -79.580 89.065 -78.675 89.155 ;
        RECT -80.885 88.885 -78.675 89.065 ;
      LAYER mcon ;
        RECT -80.695 88.975 -80.525 89.145 ;
        RECT -79.330 88.975 -79.160 89.145 ;
      LAYER met1 ;
        RECT -80.760 88.880 -79.070 89.180 ;
        RECT -80.580 88.180 -79.580 88.880 ;
    END
  END o_ranQ[21]
  PIN o_ranQ[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -85.845 94.875 -83.635 95.055 ;
        RECT -85.845 94.795 -85.340 94.875 ;
        RECT -84.540 94.785 -83.635 94.875 ;
      LAYER mcon ;
        RECT -85.655 94.795 -85.485 94.965 ;
        RECT -84.290 94.795 -84.120 94.965 ;
      LAYER met1 ;
        RECT -85.540 95.060 -84.540 95.760 ;
        RECT -85.720 94.760 -84.030 95.060 ;
    END
  END o_ranQ[22]
  PIN o_ranQ[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -90.805 89.065 -90.300 89.145 ;
        RECT -89.500 89.065 -88.595 89.155 ;
        RECT -90.805 88.885 -88.595 89.065 ;
      LAYER mcon ;
        RECT -90.615 88.975 -90.445 89.145 ;
        RECT -89.250 88.975 -89.080 89.145 ;
      LAYER met1 ;
        RECT -90.680 88.880 -88.990 89.180 ;
        RECT -90.500 88.180 -89.500 88.880 ;
    END
  END o_ranQ[23]
  PIN o_ranQ[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -95.765 94.875 -93.555 95.055 ;
        RECT -95.765 94.795 -95.260 94.875 ;
        RECT -94.460 94.785 -93.555 94.875 ;
      LAYER mcon ;
        RECT -95.575 94.795 -95.405 94.965 ;
        RECT -94.210 94.795 -94.040 94.965 ;
      LAYER met1 ;
        RECT -95.460 95.060 -94.460 95.760 ;
        RECT -95.640 94.760 -93.950 95.060 ;
    END
  END o_ranQ[24]
  PIN o_ranQ[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -100.725 89.065 -100.220 89.145 ;
        RECT -99.420 89.065 -98.515 89.155 ;
        RECT -100.725 88.885 -98.515 89.065 ;
      LAYER mcon ;
        RECT -100.535 88.975 -100.365 89.145 ;
        RECT -99.170 88.975 -99.000 89.145 ;
      LAYER met1 ;
        RECT -100.600 88.880 -98.910 89.180 ;
        RECT -100.420 88.180 -99.420 88.880 ;
    END
  END o_ranQ[25]
  PIN o_ranQ[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -105.685 94.875 -103.475 95.055 ;
        RECT -105.685 94.795 -105.180 94.875 ;
        RECT -104.380 94.785 -103.475 94.875 ;
      LAYER mcon ;
        RECT -105.495 94.795 -105.325 94.965 ;
        RECT -104.130 94.795 -103.960 94.965 ;
      LAYER met1 ;
        RECT -105.380 95.060 -104.380 95.760 ;
        RECT -105.560 94.760 -103.870 95.060 ;
    END
  END o_ranQ[26]
  PIN o_ranQ[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -110.645 89.065 -110.140 89.145 ;
        RECT -109.340 89.065 -108.435 89.155 ;
        RECT -110.645 88.885 -108.435 89.065 ;
      LAYER mcon ;
        RECT -110.455 88.975 -110.285 89.145 ;
        RECT -109.090 88.975 -108.920 89.145 ;
      LAYER met1 ;
        RECT -110.520 88.880 -108.830 89.180 ;
        RECT -110.340 88.180 -109.340 88.880 ;
    END
  END o_ranQ[27]
  PIN o_ranQ[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -115.605 94.875 -113.395 95.055 ;
        RECT -115.605 94.795 -115.100 94.875 ;
        RECT -114.300 94.785 -113.395 94.875 ;
      LAYER mcon ;
        RECT -115.415 94.795 -115.245 94.965 ;
        RECT -114.050 94.795 -113.880 94.965 ;
      LAYER met1 ;
        RECT -115.300 95.060 -114.300 95.760 ;
        RECT -115.480 94.760 -113.790 95.060 ;
    END
  END o_ranQ[28]
  PIN o_ranQ[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -120.565 89.065 -120.060 89.145 ;
        RECT -119.260 89.065 -118.355 89.155 ;
        RECT -120.565 88.885 -118.355 89.065 ;
      LAYER mcon ;
        RECT -120.375 88.975 -120.205 89.145 ;
        RECT -119.010 88.975 -118.840 89.145 ;
      LAYER met1 ;
        RECT -120.440 88.880 -118.750 89.180 ;
        RECT -120.260 88.180 -119.260 88.880 ;
    END
  END o_ranQ[29]
  PIN o_ranQ[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -125.525 94.875 -123.315 95.055 ;
        RECT -125.525 94.795 -125.020 94.875 ;
        RECT -124.220 94.785 -123.315 94.875 ;
      LAYER mcon ;
        RECT -125.335 94.795 -125.165 94.965 ;
        RECT -123.970 94.795 -123.800 94.965 ;
      LAYER met1 ;
        RECT -125.220 95.060 -124.220 95.760 ;
        RECT -125.400 94.760 -123.710 95.060 ;
    END
  END o_ranQ[30]
  PIN o_ranQ[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -130.485 89.065 -129.980 89.145 ;
        RECT -129.180 89.065 -128.275 89.155 ;
        RECT -130.485 88.885 -128.275 89.065 ;
      LAYER mcon ;
        RECT -130.295 88.975 -130.125 89.145 ;
        RECT -128.930 88.975 -128.760 89.145 ;
      LAYER met1 ;
        RECT -130.360 88.880 -128.670 89.180 ;
        RECT -130.180 88.180 -129.180 88.880 ;
    END
  END o_ranQ[31]
  PIN o_ranQ[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -140.405 89.065 -139.900 89.145 ;
        RECT -139.100 89.065 -138.195 89.155 ;
        RECT -140.405 88.885 -138.195 89.065 ;
      LAYER mcon ;
        RECT -140.215 88.975 -140.045 89.145 ;
        RECT -138.850 88.975 -138.680 89.145 ;
      LAYER met1 ;
        RECT -140.280 88.880 -138.590 89.180 ;
        RECT -140.100 88.180 -139.100 88.880 ;
    END
  END o_ranQ[33]
  PIN o_ranQ[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -145.365 94.875 -143.155 95.055 ;
        RECT -145.365 94.795 -144.860 94.875 ;
        RECT -144.060 94.785 -143.155 94.875 ;
      LAYER mcon ;
        RECT -145.175 94.795 -145.005 94.965 ;
        RECT -143.810 94.795 -143.640 94.965 ;
      LAYER met1 ;
        RECT -145.060 95.060 -144.060 95.760 ;
        RECT -145.240 94.760 -143.550 95.060 ;
    END
  END o_ranQ[34]
  PIN o_ranQ[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -150.325 89.065 -149.820 89.145 ;
        RECT -149.020 89.065 -148.115 89.155 ;
        RECT -150.325 88.885 -148.115 89.065 ;
      LAYER mcon ;
        RECT -150.135 88.975 -149.965 89.145 ;
        RECT -148.770 88.975 -148.600 89.145 ;
      LAYER met1 ;
        RECT -150.200 88.880 -148.510 89.180 ;
        RECT -150.020 88.180 -149.020 88.880 ;
    END
  END o_ranQ[35]
  PIN o_ranQ[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -135.445 94.875 -133.235 95.055 ;
        RECT -135.445 94.795 -134.940 94.875 ;
        RECT -134.140 94.785 -133.235 94.875 ;
      LAYER mcon ;
        RECT -135.255 94.795 -135.085 94.965 ;
        RECT -133.890 94.795 -133.720 94.965 ;
      LAYER met1 ;
        RECT -135.140 95.060 -134.140 95.760 ;
        RECT -135.320 94.760 -133.630 95.060 ;
    END
  END o_ranQ[32]
  PIN o_ranQ[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -155.285 94.875 -153.075 95.055 ;
        RECT -155.285 94.795 -154.780 94.875 ;
        RECT -153.980 94.785 -153.075 94.875 ;
      LAYER mcon ;
        RECT -155.095 94.795 -154.925 94.965 ;
        RECT -153.730 94.795 -153.560 94.965 ;
      LAYER met1 ;
        RECT -154.980 95.060 -153.980 95.760 ;
        RECT -155.160 94.760 -153.470 95.060 ;
    END
  END o_ranQ[36]
  PIN o_ranQ[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -160.245 89.065 -159.740 89.145 ;
        RECT -158.940 89.065 -158.035 89.155 ;
        RECT -160.245 88.885 -158.035 89.065 ;
      LAYER mcon ;
        RECT -160.055 88.975 -159.885 89.145 ;
        RECT -158.690 88.975 -158.520 89.145 ;
      LAYER met1 ;
        RECT -160.120 88.880 -158.430 89.180 ;
        RECT -159.940 88.180 -158.940 88.880 ;
    END
  END o_ranQ[37]
  PIN o_ranQ[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -165.205 94.875 -162.995 95.055 ;
        RECT -165.205 94.795 -164.700 94.875 ;
        RECT -163.900 94.785 -162.995 94.875 ;
      LAYER mcon ;
        RECT -165.015 94.795 -164.845 94.965 ;
        RECT -163.650 94.795 -163.480 94.965 ;
      LAYER met1 ;
        RECT -164.900 95.060 -163.900 95.760 ;
        RECT -165.080 94.760 -163.390 95.060 ;
    END
  END o_ranQ[38]
  PIN o_ranQ[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -170.165 89.065 -169.660 89.145 ;
        RECT -168.860 89.065 -167.955 89.155 ;
        RECT -170.165 88.885 -167.955 89.065 ;
      LAYER mcon ;
        RECT -169.975 88.975 -169.805 89.145 ;
        RECT -168.610 88.975 -168.440 89.145 ;
      LAYER met1 ;
        RECT -170.040 88.880 -168.350 89.180 ;
        RECT -169.860 88.180 -168.860 88.880 ;
    END
  END o_ranQ[39]
  PIN o_ranQ[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -175.125 94.875 -172.915 95.055 ;
        RECT -175.125 94.795 -174.620 94.875 ;
        RECT -173.820 94.785 -172.915 94.875 ;
      LAYER mcon ;
        RECT -174.935 94.795 -174.765 94.965 ;
        RECT -173.570 94.795 -173.400 94.965 ;
      LAYER met1 ;
        RECT -174.820 95.060 -173.820 95.760 ;
        RECT -175.000 94.760 -173.310 95.060 ;
    END
  END o_ranQ[40]
  PIN o_ranQ[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -180.085 89.065 -179.580 89.145 ;
        RECT -178.780 89.065 -177.875 89.155 ;
        RECT -180.085 88.885 -177.875 89.065 ;
      LAYER mcon ;
        RECT -179.895 88.975 -179.725 89.145 ;
        RECT -178.530 88.975 -178.360 89.145 ;
      LAYER met1 ;
        RECT -179.960 88.880 -178.270 89.180 ;
        RECT -179.780 88.180 -178.780 88.880 ;
    END
  END o_ranQ[41]
  PIN o_ranQ[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -185.045 94.875 -182.835 95.055 ;
        RECT -185.045 94.795 -184.540 94.875 ;
        RECT -183.740 94.785 -182.835 94.875 ;
      LAYER mcon ;
        RECT -184.855 94.795 -184.685 94.965 ;
        RECT -183.490 94.795 -183.320 94.965 ;
      LAYER met1 ;
        RECT -184.740 95.060 -183.740 95.760 ;
        RECT -184.920 94.760 -183.230 95.060 ;
    END
  END o_ranQ[42]
  PIN o_ranQ[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -190.005 89.065 -189.500 89.145 ;
        RECT -188.700 89.065 -187.795 89.155 ;
        RECT -190.005 88.885 -187.795 89.065 ;
      LAYER mcon ;
        RECT -189.815 88.975 -189.645 89.145 ;
        RECT -188.450 88.975 -188.280 89.145 ;
      LAYER met1 ;
        RECT -189.880 88.880 -188.190 89.180 ;
        RECT -189.700 88.180 -188.700 88.880 ;
    END
  END o_ranQ[43]
  PIN o_ranQ[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -194.965 94.875 -192.755 95.055 ;
        RECT -194.965 94.795 -194.460 94.875 ;
        RECT -193.660 94.785 -192.755 94.875 ;
      LAYER mcon ;
        RECT -194.775 94.795 -194.605 94.965 ;
        RECT -193.410 94.795 -193.240 94.965 ;
      LAYER met1 ;
        RECT -194.660 95.060 -193.660 95.760 ;
        RECT -194.840 94.760 -193.150 95.060 ;
    END
  END o_ranQ[44]
  PIN o_ranQ[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -199.925 89.065 -199.420 89.145 ;
        RECT -198.620 89.065 -197.715 89.155 ;
        RECT -199.925 88.885 -197.715 89.065 ;
      LAYER mcon ;
        RECT -199.735 88.975 -199.565 89.145 ;
        RECT -198.370 88.975 -198.200 89.145 ;
      LAYER met1 ;
        RECT -199.800 88.880 -198.110 89.180 ;
        RECT -199.620 88.180 -198.620 88.880 ;
    END
  END o_ranQ[45]
  PIN o_ranQ[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -204.885 94.875 -202.675 95.055 ;
        RECT -204.885 94.795 -204.380 94.875 ;
        RECT -203.580 94.785 -202.675 94.875 ;
      LAYER mcon ;
        RECT -204.695 94.795 -204.525 94.965 ;
        RECT -203.330 94.795 -203.160 94.965 ;
      LAYER met1 ;
        RECT -204.580 95.060 -203.580 95.760 ;
        RECT -204.760 94.760 -203.070 95.060 ;
    END
  END o_ranQ[46]
  PIN o_ranQ[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -209.845 89.065 -209.340 89.145 ;
        RECT -208.540 89.065 -207.635 89.155 ;
        RECT -209.845 88.885 -207.635 89.065 ;
      LAYER mcon ;
        RECT -209.655 88.975 -209.485 89.145 ;
        RECT -208.290 88.975 -208.120 89.145 ;
      LAYER met1 ;
        RECT -209.720 88.880 -208.030 89.180 ;
        RECT -209.540 88.180 -208.540 88.880 ;
    END
  END o_ranQ[47]
  PIN o_ranQ[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -219.765 89.065 -219.260 89.145 ;
        RECT -218.460 89.065 -217.555 89.155 ;
        RECT -219.765 88.885 -217.555 89.065 ;
      LAYER mcon ;
        RECT -219.575 88.975 -219.405 89.145 ;
        RECT -218.210 88.975 -218.040 89.145 ;
      LAYER met1 ;
        RECT -219.640 88.880 -217.950 89.180 ;
        RECT -219.460 88.180 -218.460 88.880 ;
    END
  END o_ranQ[49]
  PIN o_ranQ[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -224.725 94.875 -222.515 95.055 ;
        RECT -224.725 94.795 -224.220 94.875 ;
        RECT -223.420 94.785 -222.515 94.875 ;
      LAYER mcon ;
        RECT -224.535 94.795 -224.365 94.965 ;
        RECT -223.170 94.795 -223.000 94.965 ;
      LAYER met1 ;
        RECT -224.420 95.060 -223.420 95.760 ;
        RECT -224.600 94.760 -222.910 95.060 ;
    END
  END o_ranQ[50]
  PIN o_ranQ[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -229.685 89.065 -229.180 89.145 ;
        RECT -228.380 89.065 -227.475 89.155 ;
        RECT -229.685 88.885 -227.475 89.065 ;
      LAYER mcon ;
        RECT -229.495 88.975 -229.325 89.145 ;
        RECT -228.130 88.975 -227.960 89.145 ;
      LAYER met1 ;
        RECT -229.560 88.880 -227.870 89.180 ;
        RECT -229.380 88.180 -228.380 88.880 ;
    END
  END o_ranQ[51]
  PIN o_ranQ[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -214.805 94.875 -212.595 95.055 ;
        RECT -214.805 94.795 -214.300 94.875 ;
        RECT -213.500 94.785 -212.595 94.875 ;
      LAYER mcon ;
        RECT -214.615 94.795 -214.445 94.965 ;
        RECT -213.250 94.795 -213.080 94.965 ;
      LAYER met1 ;
        RECT -214.500 95.060 -213.500 95.760 ;
        RECT -214.680 94.760 -212.990 95.060 ;
    END
  END o_ranQ[48]
  PIN o_ranQ[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -234.645 94.875 -232.435 95.055 ;
        RECT -234.645 94.795 -234.140 94.875 ;
        RECT -233.340 94.785 -232.435 94.875 ;
      LAYER mcon ;
        RECT -234.455 94.795 -234.285 94.965 ;
        RECT -233.090 94.795 -232.920 94.965 ;
      LAYER met1 ;
        RECT -234.340 95.060 -233.340 95.760 ;
        RECT -234.520 94.760 -232.830 95.060 ;
    END
  END o_ranQ[52]
  PIN o_ranQ[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -239.605 89.065 -239.100 89.145 ;
        RECT -238.300 89.065 -237.395 89.155 ;
        RECT -239.605 88.885 -237.395 89.065 ;
      LAYER mcon ;
        RECT -239.415 88.975 -239.245 89.145 ;
        RECT -238.050 88.975 -237.880 89.145 ;
      LAYER met1 ;
        RECT -239.480 88.880 -237.790 89.180 ;
        RECT -239.300 88.180 -238.300 88.880 ;
    END
  END o_ranQ[53]
  PIN o_ranQ[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -244.565 94.875 -242.355 95.055 ;
        RECT -244.565 94.795 -244.060 94.875 ;
        RECT -243.260 94.785 -242.355 94.875 ;
      LAYER mcon ;
        RECT -244.375 94.795 -244.205 94.965 ;
        RECT -243.010 94.795 -242.840 94.965 ;
      LAYER met1 ;
        RECT -244.260 95.060 -243.260 95.760 ;
        RECT -244.440 94.760 -242.750 95.060 ;
    END
  END o_ranQ[54]
  PIN o_ranQ[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -249.525 89.065 -249.020 89.145 ;
        RECT -248.220 89.065 -247.315 89.155 ;
        RECT -249.525 88.885 -247.315 89.065 ;
      LAYER mcon ;
        RECT -249.335 88.975 -249.165 89.145 ;
        RECT -247.970 88.975 -247.800 89.145 ;
      LAYER met1 ;
        RECT -249.400 88.880 -247.710 89.180 ;
        RECT -249.220 88.180 -248.220 88.880 ;
    END
  END o_ranQ[55]
  PIN o_ranQ[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -254.485 94.875 -252.275 95.055 ;
        RECT -254.485 94.795 -253.980 94.875 ;
        RECT -253.180 94.785 -252.275 94.875 ;
      LAYER mcon ;
        RECT -254.295 94.795 -254.125 94.965 ;
        RECT -252.930 94.795 -252.760 94.965 ;
      LAYER met1 ;
        RECT -254.180 95.060 -253.180 95.760 ;
        RECT -254.360 94.760 -252.670 95.060 ;
    END
  END o_ranQ[56]
  PIN o_ranQ[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -259.445 89.065 -258.940 89.145 ;
        RECT -258.140 89.065 -257.235 89.155 ;
        RECT -259.445 88.885 -257.235 89.065 ;
      LAYER mcon ;
        RECT -259.255 88.975 -259.085 89.145 ;
        RECT -257.890 88.975 -257.720 89.145 ;
      LAYER met1 ;
        RECT -259.320 88.880 -257.630 89.180 ;
        RECT -259.140 88.180 -258.140 88.880 ;
    END
  END o_ranQ[57]
  PIN o_ranQ[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -264.405 94.875 -262.195 95.055 ;
        RECT -264.405 94.795 -263.900 94.875 ;
        RECT -263.100 94.785 -262.195 94.875 ;
      LAYER mcon ;
        RECT -264.215 94.795 -264.045 94.965 ;
        RECT -262.850 94.795 -262.680 94.965 ;
      LAYER met1 ;
        RECT -264.100 95.060 -263.100 95.760 ;
        RECT -264.280 94.760 -262.590 95.060 ;
    END
  END o_ranQ[58]
  PIN o_ranQ[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -269.365 89.065 -268.860 89.145 ;
        RECT -268.060 89.065 -267.155 89.155 ;
        RECT -269.365 88.885 -267.155 89.065 ;
      LAYER mcon ;
        RECT -269.175 88.975 -269.005 89.145 ;
        RECT -267.810 88.975 -267.640 89.145 ;
      LAYER met1 ;
        RECT -269.240 88.880 -267.550 89.180 ;
        RECT -269.060 88.180 -268.060 88.880 ;
    END
  END o_ranQ[59]
  PIN o_ranQ[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -274.325 94.875 -272.115 95.055 ;
        RECT -274.325 94.795 -273.820 94.875 ;
        RECT -273.020 94.785 -272.115 94.875 ;
      LAYER mcon ;
        RECT -274.135 94.795 -273.965 94.965 ;
        RECT -272.770 94.795 -272.600 94.965 ;
      LAYER met1 ;
        RECT -274.020 95.060 -273.020 95.760 ;
        RECT -274.200 94.760 -272.510 95.060 ;
    END
  END o_ranQ[60]
  PIN o_ranQ[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -279.285 89.065 -278.780 89.145 ;
        RECT -277.980 89.065 -277.075 89.155 ;
        RECT -279.285 88.885 -277.075 89.065 ;
      LAYER mcon ;
        RECT -279.095 88.975 -278.925 89.145 ;
        RECT -277.730 88.975 -277.560 89.145 ;
      LAYER met1 ;
        RECT -279.160 88.880 -277.470 89.180 ;
        RECT -278.980 88.180 -277.980 88.880 ;
    END
  END o_ranQ[61]
  PIN o_ranQ[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -284.245 94.875 -282.035 95.055 ;
        RECT -284.245 94.795 -283.740 94.875 ;
        RECT -282.940 94.785 -282.035 94.875 ;
      LAYER mcon ;
        RECT -284.055 94.795 -283.885 94.965 ;
        RECT -282.690 94.795 -282.520 94.965 ;
      LAYER met1 ;
        RECT -283.940 95.060 -282.940 95.760 ;
        RECT -284.120 94.760 -282.430 95.060 ;
    END
  END o_ranQ[62]
  PIN o_ranQ[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -289.205 89.065 -288.700 89.145 ;
        RECT -287.900 89.065 -286.995 89.155 ;
        RECT -289.205 88.885 -286.995 89.065 ;
      LAYER mcon ;
        RECT -289.015 88.975 -288.845 89.145 ;
        RECT -287.650 88.975 -287.480 89.145 ;
      LAYER met1 ;
        RECT -289.080 88.880 -287.390 89.180 ;
        RECT -288.900 88.180 -287.900 88.880 ;
    END
  END o_ranQ[63]
  PIN i_srclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 126.719994 ;
    PORT
      LAYER li1 ;
        RECT -290.905 92.005 -290.570 92.275 ;
        RECT -281.970 92.005 -281.635 92.275 ;
        RECT -280.985 92.005 -280.650 92.275 ;
        RECT -272.050 92.005 -271.715 92.275 ;
        RECT -271.065 92.005 -270.730 92.275 ;
        RECT -262.130 92.005 -261.795 92.275 ;
        RECT -261.145 92.005 -260.810 92.275 ;
        RECT -252.210 92.005 -251.875 92.275 ;
        RECT -251.225 92.005 -250.890 92.275 ;
        RECT -242.290 92.005 -241.955 92.275 ;
        RECT -241.305 92.005 -240.970 92.275 ;
        RECT -232.370 92.005 -232.035 92.275 ;
        RECT -231.385 92.005 -231.050 92.275 ;
        RECT -222.450 92.005 -222.115 92.275 ;
        RECT -221.465 92.005 -221.130 92.275 ;
        RECT -212.530 92.005 -212.195 92.275 ;
        RECT -211.545 92.005 -211.210 92.275 ;
        RECT -202.610 92.005 -202.275 92.275 ;
        RECT -201.625 92.005 -201.290 92.275 ;
        RECT -192.690 92.005 -192.355 92.275 ;
        RECT -191.705 92.005 -191.370 92.275 ;
        RECT -182.770 92.005 -182.435 92.275 ;
        RECT -181.785 92.005 -181.450 92.275 ;
        RECT -172.850 92.005 -172.515 92.275 ;
        RECT -171.865 92.005 -171.530 92.275 ;
        RECT -162.930 92.005 -162.595 92.275 ;
        RECT -161.945 92.005 -161.610 92.275 ;
        RECT -153.010 92.005 -152.675 92.275 ;
        RECT -152.025 92.005 -151.690 92.275 ;
        RECT -143.090 92.005 -142.755 92.275 ;
        RECT -142.105 92.005 -141.770 92.275 ;
        RECT -133.170 92.005 -132.835 92.275 ;
        RECT -132.185 92.005 -131.850 92.275 ;
        RECT -123.250 92.005 -122.915 92.275 ;
        RECT -122.265 92.005 -121.930 92.275 ;
        RECT -113.330 92.005 -112.995 92.275 ;
        RECT -112.345 92.005 -112.010 92.275 ;
        RECT -103.410 92.005 -103.075 92.275 ;
        RECT -102.425 92.005 -102.090 92.275 ;
        RECT -93.490 92.005 -93.155 92.275 ;
        RECT -92.505 92.005 -92.170 92.275 ;
        RECT -83.570 92.005 -83.235 92.275 ;
        RECT -82.585 92.005 -82.250 92.275 ;
        RECT -73.650 92.005 -73.315 92.275 ;
        RECT -72.665 92.005 -72.330 92.275 ;
        RECT -63.730 92.005 -63.395 92.275 ;
        RECT -62.745 92.005 -62.410 92.275 ;
        RECT -53.810 92.005 -53.475 92.275 ;
        RECT -52.825 92.005 -52.490 92.275 ;
        RECT -43.890 92.005 -43.555 92.275 ;
        RECT -42.905 92.005 -42.570 92.275 ;
        RECT -33.970 92.005 -33.635 92.275 ;
        RECT -32.985 92.005 -32.650 92.275 ;
        RECT -24.050 92.005 -23.715 92.275 ;
        RECT -23.065 92.005 -22.730 92.275 ;
        RECT -14.130 92.005 -13.795 92.275 ;
        RECT -13.145 92.005 -12.810 92.275 ;
        RECT -4.210 92.005 -3.875 92.275 ;
        RECT -3.225 92.005 -2.890 92.275 ;
        RECT 5.710 92.005 6.045 92.275 ;
        RECT 6.695 92.005 7.030 92.275 ;
        RECT 15.630 92.005 15.965 92.275 ;
        RECT 16.615 92.005 16.950 92.275 ;
        RECT 25.550 92.005 25.885 92.275 ;
        RECT -286.930 91.665 -286.595 91.935 ;
        RECT -285.945 91.665 -285.610 91.935 ;
        RECT -277.010 91.665 -276.675 91.935 ;
        RECT -276.025 91.665 -275.690 91.935 ;
        RECT -267.090 91.665 -266.755 91.935 ;
        RECT -266.105 91.665 -265.770 91.935 ;
        RECT -257.170 91.665 -256.835 91.935 ;
        RECT -256.185 91.665 -255.850 91.935 ;
        RECT -247.250 91.665 -246.915 91.935 ;
        RECT -246.265 91.665 -245.930 91.935 ;
        RECT -237.330 91.665 -236.995 91.935 ;
        RECT -236.345 91.665 -236.010 91.935 ;
        RECT -227.410 91.665 -227.075 91.935 ;
        RECT -226.425 91.665 -226.090 91.935 ;
        RECT -217.490 91.665 -217.155 91.935 ;
        RECT -216.505 91.665 -216.170 91.935 ;
        RECT -207.570 91.665 -207.235 91.935 ;
        RECT -206.585 91.665 -206.250 91.935 ;
        RECT -197.650 91.665 -197.315 91.935 ;
        RECT -196.665 91.665 -196.330 91.935 ;
        RECT -187.730 91.665 -187.395 91.935 ;
        RECT -186.745 91.665 -186.410 91.935 ;
        RECT -177.810 91.665 -177.475 91.935 ;
        RECT -176.825 91.665 -176.490 91.935 ;
        RECT -167.890 91.665 -167.555 91.935 ;
        RECT -166.905 91.665 -166.570 91.935 ;
        RECT -157.970 91.665 -157.635 91.935 ;
        RECT -156.985 91.665 -156.650 91.935 ;
        RECT -148.050 91.665 -147.715 91.935 ;
        RECT -147.065 91.665 -146.730 91.935 ;
        RECT -138.130 91.665 -137.795 91.935 ;
        RECT -137.145 91.665 -136.810 91.935 ;
        RECT -128.210 91.665 -127.875 91.935 ;
        RECT -127.225 91.665 -126.890 91.935 ;
        RECT -118.290 91.665 -117.955 91.935 ;
        RECT -117.305 91.665 -116.970 91.935 ;
        RECT -108.370 91.665 -108.035 91.935 ;
        RECT -107.385 91.665 -107.050 91.935 ;
        RECT -98.450 91.665 -98.115 91.935 ;
        RECT -97.465 91.665 -97.130 91.935 ;
        RECT -88.530 91.665 -88.195 91.935 ;
        RECT -87.545 91.665 -87.210 91.935 ;
        RECT -78.610 91.665 -78.275 91.935 ;
        RECT -77.625 91.665 -77.290 91.935 ;
        RECT -68.690 91.665 -68.355 91.935 ;
        RECT -67.705 91.665 -67.370 91.935 ;
        RECT -58.770 91.665 -58.435 91.935 ;
        RECT -57.785 91.665 -57.450 91.935 ;
        RECT -48.850 91.665 -48.515 91.935 ;
        RECT -47.865 91.665 -47.530 91.935 ;
        RECT -38.930 91.665 -38.595 91.935 ;
        RECT -37.945 91.665 -37.610 91.935 ;
        RECT -29.010 91.665 -28.675 91.935 ;
        RECT -28.025 91.665 -27.690 91.935 ;
        RECT -19.090 91.665 -18.755 91.935 ;
        RECT -18.105 91.665 -17.770 91.935 ;
        RECT -9.170 91.665 -8.835 91.935 ;
        RECT -8.185 91.665 -7.850 91.935 ;
        RECT 0.750 91.665 1.085 91.935 ;
        RECT 1.735 91.665 2.070 91.935 ;
        RECT 10.670 91.665 11.005 91.935 ;
        RECT 11.655 91.665 11.990 91.935 ;
        RECT 20.590 91.665 20.925 91.935 ;
        RECT 21.575 91.665 21.910 91.935 ;
        RECT -292.925 7.955 -292.590 8.225 ;
        RECT -283.990 7.955 -283.655 8.225 ;
        RECT -283.005 7.955 -282.670 8.225 ;
        RECT -274.070 7.955 -273.735 8.225 ;
        RECT -273.085 7.955 -272.750 8.225 ;
        RECT -264.150 7.955 -263.815 8.225 ;
        RECT -263.165 7.955 -262.830 8.225 ;
        RECT -254.230 7.955 -253.895 8.225 ;
        RECT -253.245 7.955 -252.910 8.225 ;
        RECT -244.310 7.955 -243.975 8.225 ;
        RECT -243.325 7.955 -242.990 8.225 ;
        RECT -234.390 7.955 -234.055 8.225 ;
        RECT -233.405 7.955 -233.070 8.225 ;
        RECT -224.470 7.955 -224.135 8.225 ;
        RECT -223.485 7.955 -223.150 8.225 ;
        RECT -214.550 7.955 -214.215 8.225 ;
        RECT -213.565 7.955 -213.230 8.225 ;
        RECT -204.630 7.955 -204.295 8.225 ;
        RECT -203.645 7.955 -203.310 8.225 ;
        RECT -194.710 7.955 -194.375 8.225 ;
        RECT -193.725 7.955 -193.390 8.225 ;
        RECT -184.790 7.955 -184.455 8.225 ;
        RECT -183.805 7.955 -183.470 8.225 ;
        RECT -174.870 7.955 -174.535 8.225 ;
        RECT -173.885 7.955 -173.550 8.225 ;
        RECT -164.950 7.955 -164.615 8.225 ;
        RECT -163.965 7.955 -163.630 8.225 ;
        RECT -155.030 7.955 -154.695 8.225 ;
        RECT -154.045 7.955 -153.710 8.225 ;
        RECT -145.110 7.955 -144.775 8.225 ;
        RECT -144.125 7.955 -143.790 8.225 ;
        RECT -135.190 7.955 -134.855 8.225 ;
        RECT -134.205 7.955 -133.870 8.225 ;
        RECT -125.270 7.955 -124.935 8.225 ;
        RECT -124.285 7.955 -123.950 8.225 ;
        RECT -115.350 7.955 -115.015 8.225 ;
        RECT -114.365 7.955 -114.030 8.225 ;
        RECT -105.430 7.955 -105.095 8.225 ;
        RECT -104.445 7.955 -104.110 8.225 ;
        RECT -95.510 7.955 -95.175 8.225 ;
        RECT -94.525 7.955 -94.190 8.225 ;
        RECT -85.590 7.955 -85.255 8.225 ;
        RECT -84.605 7.955 -84.270 8.225 ;
        RECT -75.670 7.955 -75.335 8.225 ;
        RECT -74.685 7.955 -74.350 8.225 ;
        RECT -65.750 7.955 -65.415 8.225 ;
        RECT -64.765 7.955 -64.430 8.225 ;
        RECT -55.830 7.955 -55.495 8.225 ;
        RECT -54.845 7.955 -54.510 8.225 ;
        RECT -45.910 7.955 -45.575 8.225 ;
        RECT -44.925 7.955 -44.590 8.225 ;
        RECT -35.990 7.955 -35.655 8.225 ;
        RECT -35.005 7.955 -34.670 8.225 ;
        RECT -26.070 7.955 -25.735 8.225 ;
        RECT -25.085 7.955 -24.750 8.225 ;
        RECT -16.150 7.955 -15.815 8.225 ;
        RECT -15.165 7.955 -14.830 8.225 ;
        RECT -6.230 7.955 -5.895 8.225 ;
        RECT -5.245 7.955 -4.910 8.225 ;
        RECT 3.690 7.955 4.025 8.225 ;
        RECT 4.675 7.955 5.010 8.225 ;
        RECT 13.610 7.955 13.945 8.225 ;
        RECT 14.595 7.955 14.930 8.225 ;
        RECT 23.530 7.955 23.865 8.225 ;
        RECT -288.950 7.615 -288.615 7.885 ;
        RECT -287.965 7.615 -287.630 7.885 ;
        RECT -279.030 7.615 -278.695 7.885 ;
        RECT -278.045 7.615 -277.710 7.885 ;
        RECT -269.110 7.615 -268.775 7.885 ;
        RECT -268.125 7.615 -267.790 7.885 ;
        RECT -259.190 7.615 -258.855 7.885 ;
        RECT -258.205 7.615 -257.870 7.885 ;
        RECT -249.270 7.615 -248.935 7.885 ;
        RECT -248.285 7.615 -247.950 7.885 ;
        RECT -239.350 7.615 -239.015 7.885 ;
        RECT -238.365 7.615 -238.030 7.885 ;
        RECT -229.430 7.615 -229.095 7.885 ;
        RECT -228.445 7.615 -228.110 7.885 ;
        RECT -219.510 7.615 -219.175 7.885 ;
        RECT -218.525 7.615 -218.190 7.885 ;
        RECT -209.590 7.615 -209.255 7.885 ;
        RECT -208.605 7.615 -208.270 7.885 ;
        RECT -199.670 7.615 -199.335 7.885 ;
        RECT -198.685 7.615 -198.350 7.885 ;
        RECT -189.750 7.615 -189.415 7.885 ;
        RECT -188.765 7.615 -188.430 7.885 ;
        RECT -179.830 7.615 -179.495 7.885 ;
        RECT -178.845 7.615 -178.510 7.885 ;
        RECT -169.910 7.615 -169.575 7.885 ;
        RECT -168.925 7.615 -168.590 7.885 ;
        RECT -159.990 7.615 -159.655 7.885 ;
        RECT -159.005 7.615 -158.670 7.885 ;
        RECT -150.070 7.615 -149.735 7.885 ;
        RECT -149.085 7.615 -148.750 7.885 ;
        RECT -140.150 7.615 -139.815 7.885 ;
        RECT -139.165 7.615 -138.830 7.885 ;
        RECT -130.230 7.615 -129.895 7.885 ;
        RECT -129.245 7.615 -128.910 7.885 ;
        RECT -120.310 7.615 -119.975 7.885 ;
        RECT -119.325 7.615 -118.990 7.885 ;
        RECT -110.390 7.615 -110.055 7.885 ;
        RECT -109.405 7.615 -109.070 7.885 ;
        RECT -100.470 7.615 -100.135 7.885 ;
        RECT -99.485 7.615 -99.150 7.885 ;
        RECT -90.550 7.615 -90.215 7.885 ;
        RECT -89.565 7.615 -89.230 7.885 ;
        RECT -80.630 7.615 -80.295 7.885 ;
        RECT -79.645 7.615 -79.310 7.885 ;
        RECT -70.710 7.615 -70.375 7.885 ;
        RECT -69.725 7.615 -69.390 7.885 ;
        RECT -60.790 7.615 -60.455 7.885 ;
        RECT -59.805 7.615 -59.470 7.885 ;
        RECT -50.870 7.615 -50.535 7.885 ;
        RECT -49.885 7.615 -49.550 7.885 ;
        RECT -40.950 7.615 -40.615 7.885 ;
        RECT -39.965 7.615 -39.630 7.885 ;
        RECT -31.030 7.615 -30.695 7.885 ;
        RECT -30.045 7.615 -29.710 7.885 ;
        RECT -21.110 7.615 -20.775 7.885 ;
        RECT -20.125 7.615 -19.790 7.885 ;
        RECT -11.190 7.615 -10.855 7.885 ;
        RECT -10.205 7.615 -9.870 7.885 ;
        RECT -1.270 7.615 -0.935 7.885 ;
        RECT -0.285 7.615 0.050 7.885 ;
        RECT 8.650 7.615 8.985 7.885 ;
        RECT 9.635 7.615 9.970 7.885 ;
        RECT 18.570 7.615 18.905 7.885 ;
        RECT 19.555 7.615 19.890 7.885 ;
        RECT -292.565 -80.995 -292.230 -80.725 ;
        RECT -283.630 -80.995 -283.295 -80.725 ;
        RECT -282.645 -80.995 -282.310 -80.725 ;
        RECT -273.710 -80.995 -273.375 -80.725 ;
        RECT -272.725 -80.995 -272.390 -80.725 ;
        RECT -263.790 -80.995 -263.455 -80.725 ;
        RECT -262.805 -80.995 -262.470 -80.725 ;
        RECT -253.870 -80.995 -253.535 -80.725 ;
        RECT -252.885 -80.995 -252.550 -80.725 ;
        RECT -243.950 -80.995 -243.615 -80.725 ;
        RECT -242.965 -80.995 -242.630 -80.725 ;
        RECT -234.030 -80.995 -233.695 -80.725 ;
        RECT -233.045 -80.995 -232.710 -80.725 ;
        RECT -224.110 -80.995 -223.775 -80.725 ;
        RECT -223.125 -80.995 -222.790 -80.725 ;
        RECT -214.190 -80.995 -213.855 -80.725 ;
        RECT -213.205 -80.995 -212.870 -80.725 ;
        RECT -204.270 -80.995 -203.935 -80.725 ;
        RECT -203.285 -80.995 -202.950 -80.725 ;
        RECT -194.350 -80.995 -194.015 -80.725 ;
        RECT -193.365 -80.995 -193.030 -80.725 ;
        RECT -184.430 -80.995 -184.095 -80.725 ;
        RECT -183.445 -80.995 -183.110 -80.725 ;
        RECT -174.510 -80.995 -174.175 -80.725 ;
        RECT -173.525 -80.995 -173.190 -80.725 ;
        RECT -164.590 -80.995 -164.255 -80.725 ;
        RECT -163.605 -80.995 -163.270 -80.725 ;
        RECT -154.670 -80.995 -154.335 -80.725 ;
        RECT -153.685 -80.995 -153.350 -80.725 ;
        RECT -144.750 -80.995 -144.415 -80.725 ;
        RECT -143.765 -80.995 -143.430 -80.725 ;
        RECT -134.830 -80.995 -134.495 -80.725 ;
        RECT -133.845 -80.995 -133.510 -80.725 ;
        RECT -124.910 -80.995 -124.575 -80.725 ;
        RECT -123.925 -80.995 -123.590 -80.725 ;
        RECT -114.990 -80.995 -114.655 -80.725 ;
        RECT -114.005 -80.995 -113.670 -80.725 ;
        RECT -105.070 -80.995 -104.735 -80.725 ;
        RECT -104.085 -80.995 -103.750 -80.725 ;
        RECT -95.150 -80.995 -94.815 -80.725 ;
        RECT -94.165 -80.995 -93.830 -80.725 ;
        RECT -85.230 -80.995 -84.895 -80.725 ;
        RECT -84.245 -80.995 -83.910 -80.725 ;
        RECT -75.310 -80.995 -74.975 -80.725 ;
        RECT -74.325 -80.995 -73.990 -80.725 ;
        RECT -65.390 -80.995 -65.055 -80.725 ;
        RECT -64.405 -80.995 -64.070 -80.725 ;
        RECT -55.470 -80.995 -55.135 -80.725 ;
        RECT -54.485 -80.995 -54.150 -80.725 ;
        RECT -45.550 -80.995 -45.215 -80.725 ;
        RECT -44.565 -80.995 -44.230 -80.725 ;
        RECT -35.630 -80.995 -35.295 -80.725 ;
        RECT -34.645 -80.995 -34.310 -80.725 ;
        RECT -25.710 -80.995 -25.375 -80.725 ;
        RECT -24.725 -80.995 -24.390 -80.725 ;
        RECT -15.790 -80.995 -15.455 -80.725 ;
        RECT -14.805 -80.995 -14.470 -80.725 ;
        RECT -5.870 -80.995 -5.535 -80.725 ;
        RECT -4.885 -80.995 -4.550 -80.725 ;
        RECT 4.050 -80.995 4.385 -80.725 ;
        RECT 5.035 -80.995 5.370 -80.725 ;
        RECT 13.970 -80.995 14.305 -80.725 ;
        RECT 14.955 -80.995 15.290 -80.725 ;
        RECT 23.890 -80.995 24.225 -80.725 ;
        RECT -288.590 -81.335 -288.255 -81.065 ;
        RECT -287.605 -81.335 -287.270 -81.065 ;
        RECT -278.670 -81.335 -278.335 -81.065 ;
        RECT -277.685 -81.335 -277.350 -81.065 ;
        RECT -268.750 -81.335 -268.415 -81.065 ;
        RECT -267.765 -81.335 -267.430 -81.065 ;
        RECT -258.830 -81.335 -258.495 -81.065 ;
        RECT -257.845 -81.335 -257.510 -81.065 ;
        RECT -248.910 -81.335 -248.575 -81.065 ;
        RECT -247.925 -81.335 -247.590 -81.065 ;
        RECT -238.990 -81.335 -238.655 -81.065 ;
        RECT -238.005 -81.335 -237.670 -81.065 ;
        RECT -229.070 -81.335 -228.735 -81.065 ;
        RECT -228.085 -81.335 -227.750 -81.065 ;
        RECT -219.150 -81.335 -218.815 -81.065 ;
        RECT -218.165 -81.335 -217.830 -81.065 ;
        RECT -209.230 -81.335 -208.895 -81.065 ;
        RECT -208.245 -81.335 -207.910 -81.065 ;
        RECT -199.310 -81.335 -198.975 -81.065 ;
        RECT -198.325 -81.335 -197.990 -81.065 ;
        RECT -189.390 -81.335 -189.055 -81.065 ;
        RECT -188.405 -81.335 -188.070 -81.065 ;
        RECT -179.470 -81.335 -179.135 -81.065 ;
        RECT -178.485 -81.335 -178.150 -81.065 ;
        RECT -169.550 -81.335 -169.215 -81.065 ;
        RECT -168.565 -81.335 -168.230 -81.065 ;
        RECT -159.630 -81.335 -159.295 -81.065 ;
        RECT -158.645 -81.335 -158.310 -81.065 ;
        RECT -149.710 -81.335 -149.375 -81.065 ;
        RECT -148.725 -81.335 -148.390 -81.065 ;
        RECT -139.790 -81.335 -139.455 -81.065 ;
        RECT -138.805 -81.335 -138.470 -81.065 ;
        RECT -129.870 -81.335 -129.535 -81.065 ;
        RECT -128.885 -81.335 -128.550 -81.065 ;
        RECT -119.950 -81.335 -119.615 -81.065 ;
        RECT -118.965 -81.335 -118.630 -81.065 ;
        RECT -110.030 -81.335 -109.695 -81.065 ;
        RECT -109.045 -81.335 -108.710 -81.065 ;
        RECT -100.110 -81.335 -99.775 -81.065 ;
        RECT -99.125 -81.335 -98.790 -81.065 ;
        RECT -90.190 -81.335 -89.855 -81.065 ;
        RECT -89.205 -81.335 -88.870 -81.065 ;
        RECT -80.270 -81.335 -79.935 -81.065 ;
        RECT -79.285 -81.335 -78.950 -81.065 ;
        RECT -70.350 -81.335 -70.015 -81.065 ;
        RECT -69.365 -81.335 -69.030 -81.065 ;
        RECT -60.430 -81.335 -60.095 -81.065 ;
        RECT -59.445 -81.335 -59.110 -81.065 ;
        RECT -50.510 -81.335 -50.175 -81.065 ;
        RECT -49.525 -81.335 -49.190 -81.065 ;
        RECT -40.590 -81.335 -40.255 -81.065 ;
        RECT -39.605 -81.335 -39.270 -81.065 ;
        RECT -30.670 -81.335 -30.335 -81.065 ;
        RECT -29.685 -81.335 -29.350 -81.065 ;
        RECT -20.750 -81.335 -20.415 -81.065 ;
        RECT -19.765 -81.335 -19.430 -81.065 ;
        RECT -10.830 -81.335 -10.495 -81.065 ;
        RECT -9.845 -81.335 -9.510 -81.065 ;
        RECT -0.910 -81.335 -0.575 -81.065 ;
        RECT 0.075 -81.335 0.410 -81.065 ;
        RECT 9.010 -81.335 9.345 -81.065 ;
        RECT 9.995 -81.335 10.330 -81.065 ;
        RECT 18.930 -81.335 19.265 -81.065 ;
        RECT 19.915 -81.335 20.250 -81.065 ;
        RECT -294.325 -175.575 -293.990 -175.305 ;
        RECT -285.390 -175.575 -285.055 -175.305 ;
        RECT -284.405 -175.575 -284.070 -175.305 ;
        RECT -275.470 -175.575 -275.135 -175.305 ;
        RECT -274.485 -175.575 -274.150 -175.305 ;
        RECT -265.550 -175.575 -265.215 -175.305 ;
        RECT -264.565 -175.575 -264.230 -175.305 ;
        RECT -255.630 -175.575 -255.295 -175.305 ;
        RECT -254.645 -175.575 -254.310 -175.305 ;
        RECT -245.710 -175.575 -245.375 -175.305 ;
        RECT -244.725 -175.575 -244.390 -175.305 ;
        RECT -235.790 -175.575 -235.455 -175.305 ;
        RECT -234.805 -175.575 -234.470 -175.305 ;
        RECT -225.870 -175.575 -225.535 -175.305 ;
        RECT -224.885 -175.575 -224.550 -175.305 ;
        RECT -215.950 -175.575 -215.615 -175.305 ;
        RECT -214.965 -175.575 -214.630 -175.305 ;
        RECT -206.030 -175.575 -205.695 -175.305 ;
        RECT -205.045 -175.575 -204.710 -175.305 ;
        RECT -196.110 -175.575 -195.775 -175.305 ;
        RECT -195.125 -175.575 -194.790 -175.305 ;
        RECT -186.190 -175.575 -185.855 -175.305 ;
        RECT -185.205 -175.575 -184.870 -175.305 ;
        RECT -176.270 -175.575 -175.935 -175.305 ;
        RECT -175.285 -175.575 -174.950 -175.305 ;
        RECT -166.350 -175.575 -166.015 -175.305 ;
        RECT -165.365 -175.575 -165.030 -175.305 ;
        RECT -156.430 -175.575 -156.095 -175.305 ;
        RECT -155.445 -175.575 -155.110 -175.305 ;
        RECT -146.510 -175.575 -146.175 -175.305 ;
        RECT -145.525 -175.575 -145.190 -175.305 ;
        RECT -136.590 -175.575 -136.255 -175.305 ;
        RECT -135.605 -175.575 -135.270 -175.305 ;
        RECT -126.670 -175.575 -126.335 -175.305 ;
        RECT -125.685 -175.575 -125.350 -175.305 ;
        RECT -116.750 -175.575 -116.415 -175.305 ;
        RECT -115.765 -175.575 -115.430 -175.305 ;
        RECT -106.830 -175.575 -106.495 -175.305 ;
        RECT -105.845 -175.575 -105.510 -175.305 ;
        RECT -96.910 -175.575 -96.575 -175.305 ;
        RECT -95.925 -175.575 -95.590 -175.305 ;
        RECT -86.990 -175.575 -86.655 -175.305 ;
        RECT -86.005 -175.575 -85.670 -175.305 ;
        RECT -77.070 -175.575 -76.735 -175.305 ;
        RECT -76.085 -175.575 -75.750 -175.305 ;
        RECT -67.150 -175.575 -66.815 -175.305 ;
        RECT -66.165 -175.575 -65.830 -175.305 ;
        RECT -57.230 -175.575 -56.895 -175.305 ;
        RECT -56.245 -175.575 -55.910 -175.305 ;
        RECT -47.310 -175.575 -46.975 -175.305 ;
        RECT -46.325 -175.575 -45.990 -175.305 ;
        RECT -37.390 -175.575 -37.055 -175.305 ;
        RECT -36.405 -175.575 -36.070 -175.305 ;
        RECT -27.470 -175.575 -27.135 -175.305 ;
        RECT -26.485 -175.575 -26.150 -175.305 ;
        RECT -17.550 -175.575 -17.215 -175.305 ;
        RECT -16.565 -175.575 -16.230 -175.305 ;
        RECT -7.630 -175.575 -7.295 -175.305 ;
        RECT -6.645 -175.575 -6.310 -175.305 ;
        RECT 2.290 -175.575 2.625 -175.305 ;
        RECT 3.275 -175.575 3.610 -175.305 ;
        RECT 12.210 -175.575 12.545 -175.305 ;
        RECT 13.195 -175.575 13.530 -175.305 ;
        RECT 22.130 -175.575 22.465 -175.305 ;
        RECT -290.350 -175.915 -290.015 -175.645 ;
        RECT -289.365 -175.915 -289.030 -175.645 ;
        RECT -280.430 -175.915 -280.095 -175.645 ;
        RECT -279.445 -175.915 -279.110 -175.645 ;
        RECT -270.510 -175.915 -270.175 -175.645 ;
        RECT -269.525 -175.915 -269.190 -175.645 ;
        RECT -260.590 -175.915 -260.255 -175.645 ;
        RECT -259.605 -175.915 -259.270 -175.645 ;
        RECT -250.670 -175.915 -250.335 -175.645 ;
        RECT -249.685 -175.915 -249.350 -175.645 ;
        RECT -240.750 -175.915 -240.415 -175.645 ;
        RECT -239.765 -175.915 -239.430 -175.645 ;
        RECT -230.830 -175.915 -230.495 -175.645 ;
        RECT -229.845 -175.915 -229.510 -175.645 ;
        RECT -220.910 -175.915 -220.575 -175.645 ;
        RECT -219.925 -175.915 -219.590 -175.645 ;
        RECT -210.990 -175.915 -210.655 -175.645 ;
        RECT -210.005 -175.915 -209.670 -175.645 ;
        RECT -201.070 -175.915 -200.735 -175.645 ;
        RECT -200.085 -175.915 -199.750 -175.645 ;
        RECT -191.150 -175.915 -190.815 -175.645 ;
        RECT -190.165 -175.915 -189.830 -175.645 ;
        RECT -181.230 -175.915 -180.895 -175.645 ;
        RECT -180.245 -175.915 -179.910 -175.645 ;
        RECT -171.310 -175.915 -170.975 -175.645 ;
        RECT -170.325 -175.915 -169.990 -175.645 ;
        RECT -161.390 -175.915 -161.055 -175.645 ;
        RECT -160.405 -175.915 -160.070 -175.645 ;
        RECT -151.470 -175.915 -151.135 -175.645 ;
        RECT -150.485 -175.915 -150.150 -175.645 ;
        RECT -141.550 -175.915 -141.215 -175.645 ;
        RECT -140.565 -175.915 -140.230 -175.645 ;
        RECT -131.630 -175.915 -131.295 -175.645 ;
        RECT -130.645 -175.915 -130.310 -175.645 ;
        RECT -121.710 -175.915 -121.375 -175.645 ;
        RECT -120.725 -175.915 -120.390 -175.645 ;
        RECT -111.790 -175.915 -111.455 -175.645 ;
        RECT -110.805 -175.915 -110.470 -175.645 ;
        RECT -101.870 -175.915 -101.535 -175.645 ;
        RECT -100.885 -175.915 -100.550 -175.645 ;
        RECT -91.950 -175.915 -91.615 -175.645 ;
        RECT -90.965 -175.915 -90.630 -175.645 ;
        RECT -82.030 -175.915 -81.695 -175.645 ;
        RECT -81.045 -175.915 -80.710 -175.645 ;
        RECT -72.110 -175.915 -71.775 -175.645 ;
        RECT -71.125 -175.915 -70.790 -175.645 ;
        RECT -62.190 -175.915 -61.855 -175.645 ;
        RECT -61.205 -175.915 -60.870 -175.645 ;
        RECT -52.270 -175.915 -51.935 -175.645 ;
        RECT -51.285 -175.915 -50.950 -175.645 ;
        RECT -42.350 -175.915 -42.015 -175.645 ;
        RECT -41.365 -175.915 -41.030 -175.645 ;
        RECT -32.430 -175.915 -32.095 -175.645 ;
        RECT -31.445 -175.915 -31.110 -175.645 ;
        RECT -22.510 -175.915 -22.175 -175.645 ;
        RECT -21.525 -175.915 -21.190 -175.645 ;
        RECT -12.590 -175.915 -12.255 -175.645 ;
        RECT -11.605 -175.915 -11.270 -175.645 ;
        RECT -2.670 -175.915 -2.335 -175.645 ;
        RECT -1.685 -175.915 -1.350 -175.645 ;
        RECT 7.250 -175.915 7.585 -175.645 ;
        RECT 8.235 -175.915 8.570 -175.645 ;
        RECT 17.170 -175.915 17.505 -175.645 ;
        RECT 18.155 -175.915 18.490 -175.645 ;
      LAYER mcon ;
        RECT -290.820 92.085 -290.650 92.255 ;
        RECT -281.890 92.085 -281.720 92.255 ;
        RECT -280.900 92.085 -280.730 92.255 ;
        RECT -271.970 92.085 -271.800 92.255 ;
        RECT -270.980 92.085 -270.810 92.255 ;
        RECT -262.050 92.085 -261.880 92.255 ;
        RECT -261.060 92.085 -260.890 92.255 ;
        RECT -252.130 92.085 -251.960 92.255 ;
        RECT -251.140 92.085 -250.970 92.255 ;
        RECT -242.210 92.085 -242.040 92.255 ;
        RECT -241.220 92.085 -241.050 92.255 ;
        RECT -232.290 92.085 -232.120 92.255 ;
        RECT -231.300 92.085 -231.130 92.255 ;
        RECT -222.370 92.085 -222.200 92.255 ;
        RECT -221.380 92.085 -221.210 92.255 ;
        RECT -212.450 92.085 -212.280 92.255 ;
        RECT -211.460 92.085 -211.290 92.255 ;
        RECT -202.530 92.085 -202.360 92.255 ;
        RECT -201.540 92.085 -201.370 92.255 ;
        RECT -192.610 92.085 -192.440 92.255 ;
        RECT -191.620 92.085 -191.450 92.255 ;
        RECT -182.690 92.085 -182.520 92.255 ;
        RECT -181.700 92.085 -181.530 92.255 ;
        RECT -172.770 92.085 -172.600 92.255 ;
        RECT -171.780 92.085 -171.610 92.255 ;
        RECT -162.850 92.085 -162.680 92.255 ;
        RECT -161.860 92.085 -161.690 92.255 ;
        RECT -152.930 92.085 -152.760 92.255 ;
        RECT -151.940 92.085 -151.770 92.255 ;
        RECT -143.010 92.085 -142.840 92.255 ;
        RECT -142.020 92.085 -141.850 92.255 ;
        RECT -133.090 92.085 -132.920 92.255 ;
        RECT -132.100 92.085 -131.930 92.255 ;
        RECT -123.170 92.085 -123.000 92.255 ;
        RECT -122.180 92.085 -122.010 92.255 ;
        RECT -113.250 92.085 -113.080 92.255 ;
        RECT -112.260 92.085 -112.090 92.255 ;
        RECT -103.330 92.085 -103.160 92.255 ;
        RECT -102.340 92.085 -102.170 92.255 ;
        RECT -93.410 92.085 -93.240 92.255 ;
        RECT -92.420 92.085 -92.250 92.255 ;
        RECT -83.490 92.085 -83.320 92.255 ;
        RECT -82.500 92.085 -82.330 92.255 ;
        RECT -73.570 92.085 -73.400 92.255 ;
        RECT -72.580 92.085 -72.410 92.255 ;
        RECT -63.650 92.085 -63.480 92.255 ;
        RECT -62.660 92.085 -62.490 92.255 ;
        RECT -53.730 92.085 -53.560 92.255 ;
        RECT -52.740 92.085 -52.570 92.255 ;
        RECT -43.810 92.085 -43.640 92.255 ;
        RECT -42.820 92.085 -42.650 92.255 ;
        RECT -33.890 92.085 -33.720 92.255 ;
        RECT -32.900 92.085 -32.730 92.255 ;
        RECT -23.970 92.085 -23.800 92.255 ;
        RECT -22.980 92.085 -22.810 92.255 ;
        RECT -14.050 92.085 -13.880 92.255 ;
        RECT -13.060 92.085 -12.890 92.255 ;
        RECT -4.130 92.085 -3.960 92.255 ;
        RECT -3.140 92.085 -2.970 92.255 ;
        RECT 5.790 92.085 5.960 92.255 ;
        RECT 6.780 92.085 6.950 92.255 ;
        RECT 15.710 92.085 15.880 92.255 ;
        RECT 16.700 92.085 16.870 92.255 ;
        RECT 25.630 92.085 25.800 92.255 ;
        RECT -286.850 91.685 -286.680 91.855 ;
        RECT -285.860 91.685 -285.690 91.855 ;
        RECT -276.930 91.685 -276.760 91.855 ;
        RECT -275.940 91.685 -275.770 91.855 ;
        RECT -267.010 91.685 -266.840 91.855 ;
        RECT -266.020 91.685 -265.850 91.855 ;
        RECT -257.090 91.685 -256.920 91.855 ;
        RECT -256.100 91.685 -255.930 91.855 ;
        RECT -247.170 91.685 -247.000 91.855 ;
        RECT -246.180 91.685 -246.010 91.855 ;
        RECT -237.250 91.685 -237.080 91.855 ;
        RECT -236.260 91.685 -236.090 91.855 ;
        RECT -227.330 91.685 -227.160 91.855 ;
        RECT -226.340 91.685 -226.170 91.855 ;
        RECT -217.410 91.685 -217.240 91.855 ;
        RECT -216.420 91.685 -216.250 91.855 ;
        RECT -207.490 91.685 -207.320 91.855 ;
        RECT -206.500 91.685 -206.330 91.855 ;
        RECT -197.570 91.685 -197.400 91.855 ;
        RECT -196.580 91.685 -196.410 91.855 ;
        RECT -187.650 91.685 -187.480 91.855 ;
        RECT -186.660 91.685 -186.490 91.855 ;
        RECT -177.730 91.685 -177.560 91.855 ;
        RECT -176.740 91.685 -176.570 91.855 ;
        RECT -167.810 91.685 -167.640 91.855 ;
        RECT -166.820 91.685 -166.650 91.855 ;
        RECT -157.890 91.685 -157.720 91.855 ;
        RECT -156.900 91.685 -156.730 91.855 ;
        RECT -147.970 91.685 -147.800 91.855 ;
        RECT -146.980 91.685 -146.810 91.855 ;
        RECT -138.050 91.685 -137.880 91.855 ;
        RECT -137.060 91.685 -136.890 91.855 ;
        RECT -128.130 91.685 -127.960 91.855 ;
        RECT -127.140 91.685 -126.970 91.855 ;
        RECT -118.210 91.685 -118.040 91.855 ;
        RECT -117.220 91.685 -117.050 91.855 ;
        RECT -108.290 91.685 -108.120 91.855 ;
        RECT -107.300 91.685 -107.130 91.855 ;
        RECT -98.370 91.685 -98.200 91.855 ;
        RECT -97.380 91.685 -97.210 91.855 ;
        RECT -88.450 91.685 -88.280 91.855 ;
        RECT -87.460 91.685 -87.290 91.855 ;
        RECT -78.530 91.685 -78.360 91.855 ;
        RECT -77.540 91.685 -77.370 91.855 ;
        RECT -68.610 91.685 -68.440 91.855 ;
        RECT -67.620 91.685 -67.450 91.855 ;
        RECT -58.690 91.685 -58.520 91.855 ;
        RECT -57.700 91.685 -57.530 91.855 ;
        RECT -48.770 91.685 -48.600 91.855 ;
        RECT -47.780 91.685 -47.610 91.855 ;
        RECT -38.850 91.685 -38.680 91.855 ;
        RECT -37.860 91.685 -37.690 91.855 ;
        RECT -28.930 91.685 -28.760 91.855 ;
        RECT -27.940 91.685 -27.770 91.855 ;
        RECT -19.010 91.685 -18.840 91.855 ;
        RECT -18.020 91.685 -17.850 91.855 ;
        RECT -9.090 91.685 -8.920 91.855 ;
        RECT -8.100 91.685 -7.930 91.855 ;
        RECT 0.830 91.685 1.000 91.855 ;
        RECT 1.820 91.685 1.990 91.855 ;
        RECT 10.750 91.685 10.920 91.855 ;
        RECT 11.740 91.685 11.910 91.855 ;
        RECT 20.670 91.685 20.840 91.855 ;
        RECT 21.660 91.685 21.830 91.855 ;
        RECT -292.840 8.035 -292.670 8.205 ;
        RECT -283.910 8.035 -283.740 8.205 ;
        RECT -282.920 8.035 -282.750 8.205 ;
        RECT -273.990 8.035 -273.820 8.205 ;
        RECT -273.000 8.035 -272.830 8.205 ;
        RECT -264.070 8.035 -263.900 8.205 ;
        RECT -263.080 8.035 -262.910 8.205 ;
        RECT -254.150 8.035 -253.980 8.205 ;
        RECT -253.160 8.035 -252.990 8.205 ;
        RECT -244.230 8.035 -244.060 8.205 ;
        RECT -243.240 8.035 -243.070 8.205 ;
        RECT -234.310 8.035 -234.140 8.205 ;
        RECT -233.320 8.035 -233.150 8.205 ;
        RECT -224.390 8.035 -224.220 8.205 ;
        RECT -223.400 8.035 -223.230 8.205 ;
        RECT -214.470 8.035 -214.300 8.205 ;
        RECT -213.480 8.035 -213.310 8.205 ;
        RECT -204.550 8.035 -204.380 8.205 ;
        RECT -203.560 8.035 -203.390 8.205 ;
        RECT -194.630 8.035 -194.460 8.205 ;
        RECT -193.640 8.035 -193.470 8.205 ;
        RECT -184.710 8.035 -184.540 8.205 ;
        RECT -183.720 8.035 -183.550 8.205 ;
        RECT -174.790 8.035 -174.620 8.205 ;
        RECT -173.800 8.035 -173.630 8.205 ;
        RECT -164.870 8.035 -164.700 8.205 ;
        RECT -163.880 8.035 -163.710 8.205 ;
        RECT -154.950 8.035 -154.780 8.205 ;
        RECT -153.960 8.035 -153.790 8.205 ;
        RECT -145.030 8.035 -144.860 8.205 ;
        RECT -144.040 8.035 -143.870 8.205 ;
        RECT -135.110 8.035 -134.940 8.205 ;
        RECT -134.120 8.035 -133.950 8.205 ;
        RECT -125.190 8.035 -125.020 8.205 ;
        RECT -124.200 8.035 -124.030 8.205 ;
        RECT -115.270 8.035 -115.100 8.205 ;
        RECT -114.280 8.035 -114.110 8.205 ;
        RECT -105.350 8.035 -105.180 8.205 ;
        RECT -104.360 8.035 -104.190 8.205 ;
        RECT -95.430 8.035 -95.260 8.205 ;
        RECT -94.440 8.035 -94.270 8.205 ;
        RECT -85.510 8.035 -85.340 8.205 ;
        RECT -84.520 8.035 -84.350 8.205 ;
        RECT -75.590 8.035 -75.420 8.205 ;
        RECT -74.600 8.035 -74.430 8.205 ;
        RECT -65.670 8.035 -65.500 8.205 ;
        RECT -64.680 8.035 -64.510 8.205 ;
        RECT -55.750 8.035 -55.580 8.205 ;
        RECT -54.760 8.035 -54.590 8.205 ;
        RECT -45.830 8.035 -45.660 8.205 ;
        RECT -44.840 8.035 -44.670 8.205 ;
        RECT -35.910 8.035 -35.740 8.205 ;
        RECT -34.920 8.035 -34.750 8.205 ;
        RECT -25.990 8.035 -25.820 8.205 ;
        RECT -25.000 8.035 -24.830 8.205 ;
        RECT -16.070 8.035 -15.900 8.205 ;
        RECT -15.080 8.035 -14.910 8.205 ;
        RECT -6.150 8.035 -5.980 8.205 ;
        RECT -5.160 8.035 -4.990 8.205 ;
        RECT 3.770 8.035 3.940 8.205 ;
        RECT 4.760 8.035 4.930 8.205 ;
        RECT 13.690 8.035 13.860 8.205 ;
        RECT 14.680 8.035 14.850 8.205 ;
        RECT 23.610 8.035 23.780 8.205 ;
        RECT -288.870 7.635 -288.700 7.805 ;
        RECT -287.880 7.635 -287.710 7.805 ;
        RECT -278.950 7.635 -278.780 7.805 ;
        RECT -277.960 7.635 -277.790 7.805 ;
        RECT -269.030 7.635 -268.860 7.805 ;
        RECT -268.040 7.635 -267.870 7.805 ;
        RECT -259.110 7.635 -258.940 7.805 ;
        RECT -258.120 7.635 -257.950 7.805 ;
        RECT -249.190 7.635 -249.020 7.805 ;
        RECT -248.200 7.635 -248.030 7.805 ;
        RECT -239.270 7.635 -239.100 7.805 ;
        RECT -238.280 7.635 -238.110 7.805 ;
        RECT -229.350 7.635 -229.180 7.805 ;
        RECT -228.360 7.635 -228.190 7.805 ;
        RECT -219.430 7.635 -219.260 7.805 ;
        RECT -218.440 7.635 -218.270 7.805 ;
        RECT -209.510 7.635 -209.340 7.805 ;
        RECT -208.520 7.635 -208.350 7.805 ;
        RECT -199.590 7.635 -199.420 7.805 ;
        RECT -198.600 7.635 -198.430 7.805 ;
        RECT -189.670 7.635 -189.500 7.805 ;
        RECT -188.680 7.635 -188.510 7.805 ;
        RECT -179.750 7.635 -179.580 7.805 ;
        RECT -178.760 7.635 -178.590 7.805 ;
        RECT -169.830 7.635 -169.660 7.805 ;
        RECT -168.840 7.635 -168.670 7.805 ;
        RECT -159.910 7.635 -159.740 7.805 ;
        RECT -158.920 7.635 -158.750 7.805 ;
        RECT -149.990 7.635 -149.820 7.805 ;
        RECT -149.000 7.635 -148.830 7.805 ;
        RECT -140.070 7.635 -139.900 7.805 ;
        RECT -139.080 7.635 -138.910 7.805 ;
        RECT -130.150 7.635 -129.980 7.805 ;
        RECT -129.160 7.635 -128.990 7.805 ;
        RECT -120.230 7.635 -120.060 7.805 ;
        RECT -119.240 7.635 -119.070 7.805 ;
        RECT -110.310 7.635 -110.140 7.805 ;
        RECT -109.320 7.635 -109.150 7.805 ;
        RECT -100.390 7.635 -100.220 7.805 ;
        RECT -99.400 7.635 -99.230 7.805 ;
        RECT -90.470 7.635 -90.300 7.805 ;
        RECT -89.480 7.635 -89.310 7.805 ;
        RECT -80.550 7.635 -80.380 7.805 ;
        RECT -79.560 7.635 -79.390 7.805 ;
        RECT -70.630 7.635 -70.460 7.805 ;
        RECT -69.640 7.635 -69.470 7.805 ;
        RECT -60.710 7.635 -60.540 7.805 ;
        RECT -59.720 7.635 -59.550 7.805 ;
        RECT -50.790 7.635 -50.620 7.805 ;
        RECT -49.800 7.635 -49.630 7.805 ;
        RECT -40.870 7.635 -40.700 7.805 ;
        RECT -39.880 7.635 -39.710 7.805 ;
        RECT -30.950 7.635 -30.780 7.805 ;
        RECT -29.960 7.635 -29.790 7.805 ;
        RECT -21.030 7.635 -20.860 7.805 ;
        RECT -20.040 7.635 -19.870 7.805 ;
        RECT -11.110 7.635 -10.940 7.805 ;
        RECT -10.120 7.635 -9.950 7.805 ;
        RECT -1.190 7.635 -1.020 7.805 ;
        RECT -0.200 7.635 -0.030 7.805 ;
        RECT 8.730 7.635 8.900 7.805 ;
        RECT 9.720 7.635 9.890 7.805 ;
        RECT 18.650 7.635 18.820 7.805 ;
        RECT 19.640 7.635 19.810 7.805 ;
        RECT -292.480 -80.915 -292.310 -80.745 ;
        RECT -283.550 -80.915 -283.380 -80.745 ;
        RECT -282.560 -80.915 -282.390 -80.745 ;
        RECT -273.630 -80.915 -273.460 -80.745 ;
        RECT -272.640 -80.915 -272.470 -80.745 ;
        RECT -263.710 -80.915 -263.540 -80.745 ;
        RECT -262.720 -80.915 -262.550 -80.745 ;
        RECT -253.790 -80.915 -253.620 -80.745 ;
        RECT -252.800 -80.915 -252.630 -80.745 ;
        RECT -243.870 -80.915 -243.700 -80.745 ;
        RECT -242.880 -80.915 -242.710 -80.745 ;
        RECT -233.950 -80.915 -233.780 -80.745 ;
        RECT -232.960 -80.915 -232.790 -80.745 ;
        RECT -224.030 -80.915 -223.860 -80.745 ;
        RECT -223.040 -80.915 -222.870 -80.745 ;
        RECT -214.110 -80.915 -213.940 -80.745 ;
        RECT -213.120 -80.915 -212.950 -80.745 ;
        RECT -204.190 -80.915 -204.020 -80.745 ;
        RECT -203.200 -80.915 -203.030 -80.745 ;
        RECT -194.270 -80.915 -194.100 -80.745 ;
        RECT -193.280 -80.915 -193.110 -80.745 ;
        RECT -184.350 -80.915 -184.180 -80.745 ;
        RECT -183.360 -80.915 -183.190 -80.745 ;
        RECT -174.430 -80.915 -174.260 -80.745 ;
        RECT -173.440 -80.915 -173.270 -80.745 ;
        RECT -164.510 -80.915 -164.340 -80.745 ;
        RECT -163.520 -80.915 -163.350 -80.745 ;
        RECT -154.590 -80.915 -154.420 -80.745 ;
        RECT -153.600 -80.915 -153.430 -80.745 ;
        RECT -144.670 -80.915 -144.500 -80.745 ;
        RECT -143.680 -80.915 -143.510 -80.745 ;
        RECT -134.750 -80.915 -134.580 -80.745 ;
        RECT -133.760 -80.915 -133.590 -80.745 ;
        RECT -124.830 -80.915 -124.660 -80.745 ;
        RECT -123.840 -80.915 -123.670 -80.745 ;
        RECT -114.910 -80.915 -114.740 -80.745 ;
        RECT -113.920 -80.915 -113.750 -80.745 ;
        RECT -104.990 -80.915 -104.820 -80.745 ;
        RECT -104.000 -80.915 -103.830 -80.745 ;
        RECT -95.070 -80.915 -94.900 -80.745 ;
        RECT -94.080 -80.915 -93.910 -80.745 ;
        RECT -85.150 -80.915 -84.980 -80.745 ;
        RECT -84.160 -80.915 -83.990 -80.745 ;
        RECT -75.230 -80.915 -75.060 -80.745 ;
        RECT -74.240 -80.915 -74.070 -80.745 ;
        RECT -65.310 -80.915 -65.140 -80.745 ;
        RECT -64.320 -80.915 -64.150 -80.745 ;
        RECT -55.390 -80.915 -55.220 -80.745 ;
        RECT -54.400 -80.915 -54.230 -80.745 ;
        RECT -45.470 -80.915 -45.300 -80.745 ;
        RECT -44.480 -80.915 -44.310 -80.745 ;
        RECT -35.550 -80.915 -35.380 -80.745 ;
        RECT -34.560 -80.915 -34.390 -80.745 ;
        RECT -25.630 -80.915 -25.460 -80.745 ;
        RECT -24.640 -80.915 -24.470 -80.745 ;
        RECT -15.710 -80.915 -15.540 -80.745 ;
        RECT -14.720 -80.915 -14.550 -80.745 ;
        RECT -5.790 -80.915 -5.620 -80.745 ;
        RECT -4.800 -80.915 -4.630 -80.745 ;
        RECT 4.130 -80.915 4.300 -80.745 ;
        RECT 5.120 -80.915 5.290 -80.745 ;
        RECT 14.050 -80.915 14.220 -80.745 ;
        RECT 15.040 -80.915 15.210 -80.745 ;
        RECT 23.970 -80.915 24.140 -80.745 ;
        RECT -288.510 -81.315 -288.340 -81.145 ;
        RECT -287.520 -81.315 -287.350 -81.145 ;
        RECT -278.590 -81.315 -278.420 -81.145 ;
        RECT -277.600 -81.315 -277.430 -81.145 ;
        RECT -268.670 -81.315 -268.500 -81.145 ;
        RECT -267.680 -81.315 -267.510 -81.145 ;
        RECT -258.750 -81.315 -258.580 -81.145 ;
        RECT -257.760 -81.315 -257.590 -81.145 ;
        RECT -248.830 -81.315 -248.660 -81.145 ;
        RECT -247.840 -81.315 -247.670 -81.145 ;
        RECT -238.910 -81.315 -238.740 -81.145 ;
        RECT -237.920 -81.315 -237.750 -81.145 ;
        RECT -228.990 -81.315 -228.820 -81.145 ;
        RECT -228.000 -81.315 -227.830 -81.145 ;
        RECT -219.070 -81.315 -218.900 -81.145 ;
        RECT -218.080 -81.315 -217.910 -81.145 ;
        RECT -209.150 -81.315 -208.980 -81.145 ;
        RECT -208.160 -81.315 -207.990 -81.145 ;
        RECT -199.230 -81.315 -199.060 -81.145 ;
        RECT -198.240 -81.315 -198.070 -81.145 ;
        RECT -189.310 -81.315 -189.140 -81.145 ;
        RECT -188.320 -81.315 -188.150 -81.145 ;
        RECT -179.390 -81.315 -179.220 -81.145 ;
        RECT -178.400 -81.315 -178.230 -81.145 ;
        RECT -169.470 -81.315 -169.300 -81.145 ;
        RECT -168.480 -81.315 -168.310 -81.145 ;
        RECT -159.550 -81.315 -159.380 -81.145 ;
        RECT -158.560 -81.315 -158.390 -81.145 ;
        RECT -149.630 -81.315 -149.460 -81.145 ;
        RECT -148.640 -81.315 -148.470 -81.145 ;
        RECT -139.710 -81.315 -139.540 -81.145 ;
        RECT -138.720 -81.315 -138.550 -81.145 ;
        RECT -129.790 -81.315 -129.620 -81.145 ;
        RECT -128.800 -81.315 -128.630 -81.145 ;
        RECT -119.870 -81.315 -119.700 -81.145 ;
        RECT -118.880 -81.315 -118.710 -81.145 ;
        RECT -109.950 -81.315 -109.780 -81.145 ;
        RECT -108.960 -81.315 -108.790 -81.145 ;
        RECT -100.030 -81.315 -99.860 -81.145 ;
        RECT -99.040 -81.315 -98.870 -81.145 ;
        RECT -90.110 -81.315 -89.940 -81.145 ;
        RECT -89.120 -81.315 -88.950 -81.145 ;
        RECT -80.190 -81.315 -80.020 -81.145 ;
        RECT -79.200 -81.315 -79.030 -81.145 ;
        RECT -70.270 -81.315 -70.100 -81.145 ;
        RECT -69.280 -81.315 -69.110 -81.145 ;
        RECT -60.350 -81.315 -60.180 -81.145 ;
        RECT -59.360 -81.315 -59.190 -81.145 ;
        RECT -50.430 -81.315 -50.260 -81.145 ;
        RECT -49.440 -81.315 -49.270 -81.145 ;
        RECT -40.510 -81.315 -40.340 -81.145 ;
        RECT -39.520 -81.315 -39.350 -81.145 ;
        RECT -30.590 -81.315 -30.420 -81.145 ;
        RECT -29.600 -81.315 -29.430 -81.145 ;
        RECT -20.670 -81.315 -20.500 -81.145 ;
        RECT -19.680 -81.315 -19.510 -81.145 ;
        RECT -10.750 -81.315 -10.580 -81.145 ;
        RECT -9.760 -81.315 -9.590 -81.145 ;
        RECT -0.830 -81.315 -0.660 -81.145 ;
        RECT 0.160 -81.315 0.330 -81.145 ;
        RECT 9.090 -81.315 9.260 -81.145 ;
        RECT 10.080 -81.315 10.250 -81.145 ;
        RECT 19.010 -81.315 19.180 -81.145 ;
        RECT 20.000 -81.315 20.170 -81.145 ;
        RECT -294.240 -175.495 -294.070 -175.325 ;
        RECT -285.310 -175.495 -285.140 -175.325 ;
        RECT -284.320 -175.495 -284.150 -175.325 ;
        RECT -275.390 -175.495 -275.220 -175.325 ;
        RECT -274.400 -175.495 -274.230 -175.325 ;
        RECT -265.470 -175.495 -265.300 -175.325 ;
        RECT -264.480 -175.495 -264.310 -175.325 ;
        RECT -255.550 -175.495 -255.380 -175.325 ;
        RECT -254.560 -175.495 -254.390 -175.325 ;
        RECT -245.630 -175.495 -245.460 -175.325 ;
        RECT -244.640 -175.495 -244.470 -175.325 ;
        RECT -235.710 -175.495 -235.540 -175.325 ;
        RECT -234.720 -175.495 -234.550 -175.325 ;
        RECT -225.790 -175.495 -225.620 -175.325 ;
        RECT -224.800 -175.495 -224.630 -175.325 ;
        RECT -215.870 -175.495 -215.700 -175.325 ;
        RECT -214.880 -175.495 -214.710 -175.325 ;
        RECT -205.950 -175.495 -205.780 -175.325 ;
        RECT -204.960 -175.495 -204.790 -175.325 ;
        RECT -196.030 -175.495 -195.860 -175.325 ;
        RECT -195.040 -175.495 -194.870 -175.325 ;
        RECT -186.110 -175.495 -185.940 -175.325 ;
        RECT -185.120 -175.495 -184.950 -175.325 ;
        RECT -176.190 -175.495 -176.020 -175.325 ;
        RECT -175.200 -175.495 -175.030 -175.325 ;
        RECT -166.270 -175.495 -166.100 -175.325 ;
        RECT -165.280 -175.495 -165.110 -175.325 ;
        RECT -156.350 -175.495 -156.180 -175.325 ;
        RECT -155.360 -175.495 -155.190 -175.325 ;
        RECT -146.430 -175.495 -146.260 -175.325 ;
        RECT -145.440 -175.495 -145.270 -175.325 ;
        RECT -136.510 -175.495 -136.340 -175.325 ;
        RECT -135.520 -175.495 -135.350 -175.325 ;
        RECT -126.590 -175.495 -126.420 -175.325 ;
        RECT -125.600 -175.495 -125.430 -175.325 ;
        RECT -116.670 -175.495 -116.500 -175.325 ;
        RECT -115.680 -175.495 -115.510 -175.325 ;
        RECT -106.750 -175.495 -106.580 -175.325 ;
        RECT -105.760 -175.495 -105.590 -175.325 ;
        RECT -96.830 -175.495 -96.660 -175.325 ;
        RECT -95.840 -175.495 -95.670 -175.325 ;
        RECT -86.910 -175.495 -86.740 -175.325 ;
        RECT -85.920 -175.495 -85.750 -175.325 ;
        RECT -76.990 -175.495 -76.820 -175.325 ;
        RECT -76.000 -175.495 -75.830 -175.325 ;
        RECT -67.070 -175.495 -66.900 -175.325 ;
        RECT -66.080 -175.495 -65.910 -175.325 ;
        RECT -57.150 -175.495 -56.980 -175.325 ;
        RECT -56.160 -175.495 -55.990 -175.325 ;
        RECT -47.230 -175.495 -47.060 -175.325 ;
        RECT -46.240 -175.495 -46.070 -175.325 ;
        RECT -37.310 -175.495 -37.140 -175.325 ;
        RECT -36.320 -175.495 -36.150 -175.325 ;
        RECT -27.390 -175.495 -27.220 -175.325 ;
        RECT -26.400 -175.495 -26.230 -175.325 ;
        RECT -17.470 -175.495 -17.300 -175.325 ;
        RECT -16.480 -175.495 -16.310 -175.325 ;
        RECT -7.550 -175.495 -7.380 -175.325 ;
        RECT -6.560 -175.495 -6.390 -175.325 ;
        RECT 2.370 -175.495 2.540 -175.325 ;
        RECT 3.360 -175.495 3.530 -175.325 ;
        RECT 12.290 -175.495 12.460 -175.325 ;
        RECT 13.280 -175.495 13.450 -175.325 ;
        RECT 22.210 -175.495 22.380 -175.325 ;
        RECT -290.270 -175.895 -290.100 -175.725 ;
        RECT -289.280 -175.895 -289.110 -175.725 ;
        RECT -280.350 -175.895 -280.180 -175.725 ;
        RECT -279.360 -175.895 -279.190 -175.725 ;
        RECT -270.430 -175.895 -270.260 -175.725 ;
        RECT -269.440 -175.895 -269.270 -175.725 ;
        RECT -260.510 -175.895 -260.340 -175.725 ;
        RECT -259.520 -175.895 -259.350 -175.725 ;
        RECT -250.590 -175.895 -250.420 -175.725 ;
        RECT -249.600 -175.895 -249.430 -175.725 ;
        RECT -240.670 -175.895 -240.500 -175.725 ;
        RECT -239.680 -175.895 -239.510 -175.725 ;
        RECT -230.750 -175.895 -230.580 -175.725 ;
        RECT -229.760 -175.895 -229.590 -175.725 ;
        RECT -220.830 -175.895 -220.660 -175.725 ;
        RECT -219.840 -175.895 -219.670 -175.725 ;
        RECT -210.910 -175.895 -210.740 -175.725 ;
        RECT -209.920 -175.895 -209.750 -175.725 ;
        RECT -200.990 -175.895 -200.820 -175.725 ;
        RECT -200.000 -175.895 -199.830 -175.725 ;
        RECT -191.070 -175.895 -190.900 -175.725 ;
        RECT -190.080 -175.895 -189.910 -175.725 ;
        RECT -181.150 -175.895 -180.980 -175.725 ;
        RECT -180.160 -175.895 -179.990 -175.725 ;
        RECT -171.230 -175.895 -171.060 -175.725 ;
        RECT -170.240 -175.895 -170.070 -175.725 ;
        RECT -161.310 -175.895 -161.140 -175.725 ;
        RECT -160.320 -175.895 -160.150 -175.725 ;
        RECT -151.390 -175.895 -151.220 -175.725 ;
        RECT -150.400 -175.895 -150.230 -175.725 ;
        RECT -141.470 -175.895 -141.300 -175.725 ;
        RECT -140.480 -175.895 -140.310 -175.725 ;
        RECT -131.550 -175.895 -131.380 -175.725 ;
        RECT -130.560 -175.895 -130.390 -175.725 ;
        RECT -121.630 -175.895 -121.460 -175.725 ;
        RECT -120.640 -175.895 -120.470 -175.725 ;
        RECT -111.710 -175.895 -111.540 -175.725 ;
        RECT -110.720 -175.895 -110.550 -175.725 ;
        RECT -101.790 -175.895 -101.620 -175.725 ;
        RECT -100.800 -175.895 -100.630 -175.725 ;
        RECT -91.870 -175.895 -91.700 -175.725 ;
        RECT -90.880 -175.895 -90.710 -175.725 ;
        RECT -81.950 -175.895 -81.780 -175.725 ;
        RECT -80.960 -175.895 -80.790 -175.725 ;
        RECT -72.030 -175.895 -71.860 -175.725 ;
        RECT -71.040 -175.895 -70.870 -175.725 ;
        RECT -62.110 -175.895 -61.940 -175.725 ;
        RECT -61.120 -175.895 -60.950 -175.725 ;
        RECT -52.190 -175.895 -52.020 -175.725 ;
        RECT -51.200 -175.895 -51.030 -175.725 ;
        RECT -42.270 -175.895 -42.100 -175.725 ;
        RECT -41.280 -175.895 -41.110 -175.725 ;
        RECT -32.350 -175.895 -32.180 -175.725 ;
        RECT -31.360 -175.895 -31.190 -175.725 ;
        RECT -22.430 -175.895 -22.260 -175.725 ;
        RECT -21.440 -175.895 -21.270 -175.725 ;
        RECT -12.510 -175.895 -12.340 -175.725 ;
        RECT -11.520 -175.895 -11.350 -175.725 ;
        RECT -2.590 -175.895 -2.420 -175.725 ;
        RECT -1.600 -175.895 -1.430 -175.725 ;
        RECT 7.330 -175.895 7.500 -175.725 ;
        RECT 8.320 -175.895 8.490 -175.725 ;
        RECT 17.250 -175.895 17.420 -175.725 ;
        RECT 18.240 -175.895 18.410 -175.725 ;
      LAYER met1 ;
        RECT -291.010 91.900 -290.550 92.350 ;
        RECT -286.950 91.590 -286.490 92.040 ;
        RECT -286.050 91.590 -285.590 92.040 ;
        RECT -281.990 91.900 -281.530 92.350 ;
        RECT -281.090 91.900 -280.630 92.350 ;
        RECT -277.030 91.590 -276.570 92.040 ;
        RECT -276.130 91.590 -275.670 92.040 ;
        RECT -272.070 91.900 -271.610 92.350 ;
        RECT -271.170 91.900 -270.710 92.350 ;
        RECT -267.110 91.590 -266.650 92.040 ;
        RECT -266.210 91.590 -265.750 92.040 ;
        RECT -262.150 91.900 -261.690 92.350 ;
        RECT -261.250 91.900 -260.790 92.350 ;
        RECT -257.190 91.590 -256.730 92.040 ;
        RECT -256.290 91.590 -255.830 92.040 ;
        RECT -252.230 91.900 -251.770 92.350 ;
        RECT -251.330 91.900 -250.870 92.350 ;
        RECT -247.270 91.590 -246.810 92.040 ;
        RECT -246.370 91.590 -245.910 92.040 ;
        RECT -242.310 91.900 -241.850 92.350 ;
        RECT -241.410 91.900 -240.950 92.350 ;
        RECT -237.350 91.590 -236.890 92.040 ;
        RECT -236.450 91.590 -235.990 92.040 ;
        RECT -232.390 91.900 -231.930 92.350 ;
        RECT -231.490 91.900 -231.030 92.350 ;
        RECT -227.430 91.590 -226.970 92.040 ;
        RECT -226.530 91.590 -226.070 92.040 ;
        RECT -222.470 91.900 -222.010 92.350 ;
        RECT -221.570 91.900 -221.110 92.350 ;
        RECT -217.510 91.590 -217.050 92.040 ;
        RECT -216.610 91.590 -216.150 92.040 ;
        RECT -212.550 91.900 -212.090 92.350 ;
        RECT -211.650 91.900 -211.190 92.350 ;
        RECT -207.590 91.590 -207.130 92.040 ;
        RECT -206.690 91.590 -206.230 92.040 ;
        RECT -202.630 91.900 -202.170 92.350 ;
        RECT -201.730 91.900 -201.270 92.350 ;
        RECT -197.670 91.590 -197.210 92.040 ;
        RECT -196.770 91.590 -196.310 92.040 ;
        RECT -192.710 91.900 -192.250 92.350 ;
        RECT -191.810 91.900 -191.350 92.350 ;
        RECT -187.750 91.590 -187.290 92.040 ;
        RECT -186.850 91.590 -186.390 92.040 ;
        RECT -182.790 91.900 -182.330 92.350 ;
        RECT -181.890 91.900 -181.430 92.350 ;
        RECT -177.830 91.590 -177.370 92.040 ;
        RECT -176.930 91.590 -176.470 92.040 ;
        RECT -172.870 91.900 -172.410 92.350 ;
        RECT -171.970 91.900 -171.510 92.350 ;
        RECT -167.910 91.590 -167.450 92.040 ;
        RECT -167.010 91.590 -166.550 92.040 ;
        RECT -162.950 91.900 -162.490 92.350 ;
        RECT -162.050 91.900 -161.590 92.350 ;
        RECT -157.990 91.590 -157.530 92.040 ;
        RECT -157.090 91.590 -156.630 92.040 ;
        RECT -153.030 91.900 -152.570 92.350 ;
        RECT -152.130 91.900 -151.670 92.350 ;
        RECT -148.070 91.590 -147.610 92.040 ;
        RECT -147.170 91.590 -146.710 92.040 ;
        RECT -143.110 91.900 -142.650 92.350 ;
        RECT -142.210 91.900 -141.750 92.350 ;
        RECT -138.150 91.590 -137.690 92.040 ;
        RECT -137.250 91.590 -136.790 92.040 ;
        RECT -133.190 91.900 -132.730 92.350 ;
        RECT -132.290 91.900 -131.830 92.350 ;
        RECT -128.230 91.590 -127.770 92.040 ;
        RECT -127.330 91.590 -126.870 92.040 ;
        RECT -123.270 91.900 -122.810 92.350 ;
        RECT -122.370 91.900 -121.910 92.350 ;
        RECT -118.310 91.590 -117.850 92.040 ;
        RECT -117.410 91.590 -116.950 92.040 ;
        RECT -113.350 91.900 -112.890 92.350 ;
        RECT -112.450 91.900 -111.990 92.350 ;
        RECT -108.390 91.590 -107.930 92.040 ;
        RECT -107.490 91.590 -107.030 92.040 ;
        RECT -103.430 91.900 -102.970 92.350 ;
        RECT -102.530 91.900 -102.070 92.350 ;
        RECT -98.470 91.590 -98.010 92.040 ;
        RECT -97.570 91.590 -97.110 92.040 ;
        RECT -93.510 91.900 -93.050 92.350 ;
        RECT -92.610 91.900 -92.150 92.350 ;
        RECT -88.550 91.590 -88.090 92.040 ;
        RECT -87.650 91.590 -87.190 92.040 ;
        RECT -83.590 91.900 -83.130 92.350 ;
        RECT -82.690 91.900 -82.230 92.350 ;
        RECT -78.630 91.590 -78.170 92.040 ;
        RECT -77.730 91.590 -77.270 92.040 ;
        RECT -73.670 91.900 -73.210 92.350 ;
        RECT -72.770 91.900 -72.310 92.350 ;
        RECT -68.710 91.590 -68.250 92.040 ;
        RECT -67.810 91.590 -67.350 92.040 ;
        RECT -63.750 91.900 -63.290 92.350 ;
        RECT -62.850 91.900 -62.390 92.350 ;
        RECT -58.790 91.590 -58.330 92.040 ;
        RECT -57.890 91.590 -57.430 92.040 ;
        RECT -53.830 91.900 -53.370 92.350 ;
        RECT -52.930 91.900 -52.470 92.350 ;
        RECT -48.870 91.590 -48.410 92.040 ;
        RECT -47.970 91.590 -47.510 92.040 ;
        RECT -43.910 91.900 -43.450 92.350 ;
        RECT -43.010 91.900 -42.550 92.350 ;
        RECT -38.950 91.590 -38.490 92.040 ;
        RECT -38.050 91.590 -37.590 92.040 ;
        RECT -33.990 91.900 -33.530 92.350 ;
        RECT -33.090 91.900 -32.630 92.350 ;
        RECT -29.030 91.590 -28.570 92.040 ;
        RECT -28.130 91.590 -27.670 92.040 ;
        RECT -24.070 91.900 -23.610 92.350 ;
        RECT -23.170 91.900 -22.710 92.350 ;
        RECT -19.110 91.590 -18.650 92.040 ;
        RECT -18.210 91.590 -17.750 92.040 ;
        RECT -14.150 91.900 -13.690 92.350 ;
        RECT -13.250 91.900 -12.790 92.350 ;
        RECT -9.190 91.590 -8.730 92.040 ;
        RECT -8.290 91.590 -7.830 92.040 ;
        RECT -4.230 91.900 -3.770 92.350 ;
        RECT -3.330 91.900 -2.870 92.350 ;
        RECT 0.730 91.590 1.190 92.040 ;
        RECT 1.630 91.590 2.090 92.040 ;
        RECT 5.690 91.900 6.150 92.350 ;
        RECT 6.590 91.900 7.050 92.350 ;
        RECT 10.650 91.590 11.110 92.040 ;
        RECT 11.550 91.590 12.010 92.040 ;
        RECT 15.610 91.900 16.070 92.350 ;
        RECT 16.510 91.900 16.970 92.350 ;
        RECT 20.570 91.590 21.030 92.040 ;
        RECT 21.470 91.590 21.930 92.040 ;
        RECT 25.530 91.900 25.990 92.350 ;
        RECT -293.030 7.850 -292.570 8.300 ;
        RECT -288.970 7.540 -288.510 7.990 ;
        RECT -288.070 7.540 -287.610 7.990 ;
        RECT -284.010 7.850 -283.550 8.300 ;
        RECT -283.110 7.850 -282.650 8.300 ;
        RECT -279.050 7.540 -278.590 7.990 ;
        RECT -278.150 7.540 -277.690 7.990 ;
        RECT -274.090 7.850 -273.630 8.300 ;
        RECT -273.190 7.850 -272.730 8.300 ;
        RECT -269.130 7.540 -268.670 7.990 ;
        RECT -268.230 7.540 -267.770 7.990 ;
        RECT -264.170 7.850 -263.710 8.300 ;
        RECT -263.270 7.850 -262.810 8.300 ;
        RECT -259.210 7.540 -258.750 7.990 ;
        RECT -258.310 7.540 -257.850 7.990 ;
        RECT -254.250 7.850 -253.790 8.300 ;
        RECT -253.350 7.850 -252.890 8.300 ;
        RECT -249.290 7.540 -248.830 7.990 ;
        RECT -248.390 7.540 -247.930 7.990 ;
        RECT -244.330 7.850 -243.870 8.300 ;
        RECT -243.430 7.850 -242.970 8.300 ;
        RECT -239.370 7.540 -238.910 7.990 ;
        RECT -238.470 7.540 -238.010 7.990 ;
        RECT -234.410 7.850 -233.950 8.300 ;
        RECT -233.510 7.850 -233.050 8.300 ;
        RECT -229.450 7.540 -228.990 7.990 ;
        RECT -228.550 7.540 -228.090 7.990 ;
        RECT -224.490 7.850 -224.030 8.300 ;
        RECT -223.590 7.850 -223.130 8.300 ;
        RECT -219.530 7.540 -219.070 7.990 ;
        RECT -218.630 7.540 -218.170 7.990 ;
        RECT -214.570 7.850 -214.110 8.300 ;
        RECT -213.670 7.850 -213.210 8.300 ;
        RECT -209.610 7.540 -209.150 7.990 ;
        RECT -208.710 7.540 -208.250 7.990 ;
        RECT -204.650 7.850 -204.190 8.300 ;
        RECT -203.750 7.850 -203.290 8.300 ;
        RECT -199.690 7.540 -199.230 7.990 ;
        RECT -198.790 7.540 -198.330 7.990 ;
        RECT -194.730 7.850 -194.270 8.300 ;
        RECT -193.830 7.850 -193.370 8.300 ;
        RECT -189.770 7.540 -189.310 7.990 ;
        RECT -188.870 7.540 -188.410 7.990 ;
        RECT -184.810 7.850 -184.350 8.300 ;
        RECT -183.910 7.850 -183.450 8.300 ;
        RECT -179.850 7.540 -179.390 7.990 ;
        RECT -178.950 7.540 -178.490 7.990 ;
        RECT -174.890 7.850 -174.430 8.300 ;
        RECT -173.990 7.850 -173.530 8.300 ;
        RECT -169.930 7.540 -169.470 7.990 ;
        RECT -169.030 7.540 -168.570 7.990 ;
        RECT -164.970 7.850 -164.510 8.300 ;
        RECT -164.070 7.850 -163.610 8.300 ;
        RECT -160.010 7.540 -159.550 7.990 ;
        RECT -159.110 7.540 -158.650 7.990 ;
        RECT -155.050 7.850 -154.590 8.300 ;
        RECT -154.150 7.850 -153.690 8.300 ;
        RECT -150.090 7.540 -149.630 7.990 ;
        RECT -149.190 7.540 -148.730 7.990 ;
        RECT -145.130 7.850 -144.670 8.300 ;
        RECT -144.230 7.850 -143.770 8.300 ;
        RECT -140.170 7.540 -139.710 7.990 ;
        RECT -139.270 7.540 -138.810 7.990 ;
        RECT -135.210 7.850 -134.750 8.300 ;
        RECT -134.310 7.850 -133.850 8.300 ;
        RECT -130.250 7.540 -129.790 7.990 ;
        RECT -129.350 7.540 -128.890 7.990 ;
        RECT -125.290 7.850 -124.830 8.300 ;
        RECT -124.390 7.850 -123.930 8.300 ;
        RECT -120.330 7.540 -119.870 7.990 ;
        RECT -119.430 7.540 -118.970 7.990 ;
        RECT -115.370 7.850 -114.910 8.300 ;
        RECT -114.470 7.850 -114.010 8.300 ;
        RECT -110.410 7.540 -109.950 7.990 ;
        RECT -109.510 7.540 -109.050 7.990 ;
        RECT -105.450 7.850 -104.990 8.300 ;
        RECT -104.550 7.850 -104.090 8.300 ;
        RECT -100.490 7.540 -100.030 7.990 ;
        RECT -99.590 7.540 -99.130 7.990 ;
        RECT -95.530 7.850 -95.070 8.300 ;
        RECT -94.630 7.850 -94.170 8.300 ;
        RECT -90.570 7.540 -90.110 7.990 ;
        RECT -89.670 7.540 -89.210 7.990 ;
        RECT -85.610 7.850 -85.150 8.300 ;
        RECT -84.710 7.850 -84.250 8.300 ;
        RECT -80.650 7.540 -80.190 7.990 ;
        RECT -79.750 7.540 -79.290 7.990 ;
        RECT -75.690 7.850 -75.230 8.300 ;
        RECT -74.790 7.850 -74.330 8.300 ;
        RECT -70.730 7.540 -70.270 7.990 ;
        RECT -69.830 7.540 -69.370 7.990 ;
        RECT -65.770 7.850 -65.310 8.300 ;
        RECT -64.870 7.850 -64.410 8.300 ;
        RECT -60.810 7.540 -60.350 7.990 ;
        RECT -59.910 7.540 -59.450 7.990 ;
        RECT -55.850 7.850 -55.390 8.300 ;
        RECT -54.950 7.850 -54.490 8.300 ;
        RECT -50.890 7.540 -50.430 7.990 ;
        RECT -49.990 7.540 -49.530 7.990 ;
        RECT -45.930 7.850 -45.470 8.300 ;
        RECT -45.030 7.850 -44.570 8.300 ;
        RECT -40.970 7.540 -40.510 7.990 ;
        RECT -40.070 7.540 -39.610 7.990 ;
        RECT -36.010 7.850 -35.550 8.300 ;
        RECT -35.110 7.850 -34.650 8.300 ;
        RECT -31.050 7.540 -30.590 7.990 ;
        RECT -30.150 7.540 -29.690 7.990 ;
        RECT -26.090 7.850 -25.630 8.300 ;
        RECT -25.190 7.850 -24.730 8.300 ;
        RECT -21.130 7.540 -20.670 7.990 ;
        RECT -20.230 7.540 -19.770 7.990 ;
        RECT -16.170 7.850 -15.710 8.300 ;
        RECT -15.270 7.850 -14.810 8.300 ;
        RECT -11.210 7.540 -10.750 7.990 ;
        RECT -10.310 7.540 -9.850 7.990 ;
        RECT -6.250 7.850 -5.790 8.300 ;
        RECT -5.350 7.850 -4.890 8.300 ;
        RECT -1.290 7.540 -0.830 7.990 ;
        RECT -0.390 7.540 0.070 7.990 ;
        RECT 3.670 7.850 4.130 8.300 ;
        RECT 4.570 7.850 5.030 8.300 ;
        RECT 8.630 7.540 9.090 7.990 ;
        RECT 9.530 7.540 9.990 7.990 ;
        RECT 13.590 7.850 14.050 8.300 ;
        RECT 14.490 7.850 14.950 8.300 ;
        RECT 18.550 7.540 19.010 7.990 ;
        RECT 19.450 7.540 19.910 7.990 ;
        RECT 23.510 7.850 23.970 8.300 ;
        RECT -292.670 -81.100 -292.210 -80.650 ;
        RECT -288.610 -81.410 -288.150 -80.960 ;
        RECT -287.710 -81.410 -287.250 -80.960 ;
        RECT -283.650 -81.100 -283.190 -80.650 ;
        RECT -282.750 -81.100 -282.290 -80.650 ;
        RECT -278.690 -81.410 -278.230 -80.960 ;
        RECT -277.790 -81.410 -277.330 -80.960 ;
        RECT -273.730 -81.100 -273.270 -80.650 ;
        RECT -272.830 -81.100 -272.370 -80.650 ;
        RECT -268.770 -81.410 -268.310 -80.960 ;
        RECT -267.870 -81.410 -267.410 -80.960 ;
        RECT -263.810 -81.100 -263.350 -80.650 ;
        RECT -262.910 -81.100 -262.450 -80.650 ;
        RECT -258.850 -81.410 -258.390 -80.960 ;
        RECT -257.950 -81.410 -257.490 -80.960 ;
        RECT -253.890 -81.100 -253.430 -80.650 ;
        RECT -252.990 -81.100 -252.530 -80.650 ;
        RECT -248.930 -81.410 -248.470 -80.960 ;
        RECT -248.030 -81.410 -247.570 -80.960 ;
        RECT -243.970 -81.100 -243.510 -80.650 ;
        RECT -243.070 -81.100 -242.610 -80.650 ;
        RECT -239.010 -81.410 -238.550 -80.960 ;
        RECT -238.110 -81.410 -237.650 -80.960 ;
        RECT -234.050 -81.100 -233.590 -80.650 ;
        RECT -233.150 -81.100 -232.690 -80.650 ;
        RECT -229.090 -81.410 -228.630 -80.960 ;
        RECT -228.190 -81.410 -227.730 -80.960 ;
        RECT -224.130 -81.100 -223.670 -80.650 ;
        RECT -223.230 -81.100 -222.770 -80.650 ;
        RECT -219.170 -81.410 -218.710 -80.960 ;
        RECT -218.270 -81.410 -217.810 -80.960 ;
        RECT -214.210 -81.100 -213.750 -80.650 ;
        RECT -213.310 -81.100 -212.850 -80.650 ;
        RECT -209.250 -81.410 -208.790 -80.960 ;
        RECT -208.350 -81.410 -207.890 -80.960 ;
        RECT -204.290 -81.100 -203.830 -80.650 ;
        RECT -203.390 -81.100 -202.930 -80.650 ;
        RECT -199.330 -81.410 -198.870 -80.960 ;
        RECT -198.430 -81.410 -197.970 -80.960 ;
        RECT -194.370 -81.100 -193.910 -80.650 ;
        RECT -193.470 -81.100 -193.010 -80.650 ;
        RECT -189.410 -81.410 -188.950 -80.960 ;
        RECT -188.510 -81.410 -188.050 -80.960 ;
        RECT -184.450 -81.100 -183.990 -80.650 ;
        RECT -183.550 -81.100 -183.090 -80.650 ;
        RECT -179.490 -81.410 -179.030 -80.960 ;
        RECT -178.590 -81.410 -178.130 -80.960 ;
        RECT -174.530 -81.100 -174.070 -80.650 ;
        RECT -173.630 -81.100 -173.170 -80.650 ;
        RECT -169.570 -81.410 -169.110 -80.960 ;
        RECT -168.670 -81.410 -168.210 -80.960 ;
        RECT -164.610 -81.100 -164.150 -80.650 ;
        RECT -163.710 -81.100 -163.250 -80.650 ;
        RECT -159.650 -81.410 -159.190 -80.960 ;
        RECT -158.750 -81.410 -158.290 -80.960 ;
        RECT -154.690 -81.100 -154.230 -80.650 ;
        RECT -153.790 -81.100 -153.330 -80.650 ;
        RECT -149.730 -81.410 -149.270 -80.960 ;
        RECT -148.830 -81.410 -148.370 -80.960 ;
        RECT -144.770 -81.100 -144.310 -80.650 ;
        RECT -143.870 -81.100 -143.410 -80.650 ;
        RECT -139.810 -81.410 -139.350 -80.960 ;
        RECT -138.910 -81.410 -138.450 -80.960 ;
        RECT -134.850 -81.100 -134.390 -80.650 ;
        RECT -133.950 -81.100 -133.490 -80.650 ;
        RECT -129.890 -81.410 -129.430 -80.960 ;
        RECT -128.990 -81.410 -128.530 -80.960 ;
        RECT -124.930 -81.100 -124.470 -80.650 ;
        RECT -124.030 -81.100 -123.570 -80.650 ;
        RECT -119.970 -81.410 -119.510 -80.960 ;
        RECT -119.070 -81.410 -118.610 -80.960 ;
        RECT -115.010 -81.100 -114.550 -80.650 ;
        RECT -114.110 -81.100 -113.650 -80.650 ;
        RECT -110.050 -81.410 -109.590 -80.960 ;
        RECT -109.150 -81.410 -108.690 -80.960 ;
        RECT -105.090 -81.100 -104.630 -80.650 ;
        RECT -104.190 -81.100 -103.730 -80.650 ;
        RECT -100.130 -81.410 -99.670 -80.960 ;
        RECT -99.230 -81.410 -98.770 -80.960 ;
        RECT -95.170 -81.100 -94.710 -80.650 ;
        RECT -94.270 -81.100 -93.810 -80.650 ;
        RECT -90.210 -81.410 -89.750 -80.960 ;
        RECT -89.310 -81.410 -88.850 -80.960 ;
        RECT -85.250 -81.100 -84.790 -80.650 ;
        RECT -84.350 -81.100 -83.890 -80.650 ;
        RECT -80.290 -81.410 -79.830 -80.960 ;
        RECT -79.390 -81.410 -78.930 -80.960 ;
        RECT -75.330 -81.100 -74.870 -80.650 ;
        RECT -74.430 -81.100 -73.970 -80.650 ;
        RECT -70.370 -81.410 -69.910 -80.960 ;
        RECT -69.470 -81.410 -69.010 -80.960 ;
        RECT -65.410 -81.100 -64.950 -80.650 ;
        RECT -64.510 -81.100 -64.050 -80.650 ;
        RECT -60.450 -81.410 -59.990 -80.960 ;
        RECT -59.550 -81.410 -59.090 -80.960 ;
        RECT -55.490 -81.100 -55.030 -80.650 ;
        RECT -54.590 -81.100 -54.130 -80.650 ;
        RECT -50.530 -81.410 -50.070 -80.960 ;
        RECT -49.630 -81.410 -49.170 -80.960 ;
        RECT -45.570 -81.100 -45.110 -80.650 ;
        RECT -44.670 -81.100 -44.210 -80.650 ;
        RECT -40.610 -81.410 -40.150 -80.960 ;
        RECT -39.710 -81.410 -39.250 -80.960 ;
        RECT -35.650 -81.100 -35.190 -80.650 ;
        RECT -34.750 -81.100 -34.290 -80.650 ;
        RECT -30.690 -81.410 -30.230 -80.960 ;
        RECT -29.790 -81.410 -29.330 -80.960 ;
        RECT -25.730 -81.100 -25.270 -80.650 ;
        RECT -24.830 -81.100 -24.370 -80.650 ;
        RECT -20.770 -81.410 -20.310 -80.960 ;
        RECT -19.870 -81.410 -19.410 -80.960 ;
        RECT -15.810 -81.100 -15.350 -80.650 ;
        RECT -14.910 -81.100 -14.450 -80.650 ;
        RECT -10.850 -81.410 -10.390 -80.960 ;
        RECT -9.950 -81.410 -9.490 -80.960 ;
        RECT -5.890 -81.100 -5.430 -80.650 ;
        RECT -4.990 -81.100 -4.530 -80.650 ;
        RECT -0.930 -81.410 -0.470 -80.960 ;
        RECT -0.030 -81.410 0.430 -80.960 ;
        RECT 4.030 -81.100 4.490 -80.650 ;
        RECT 4.930 -81.100 5.390 -80.650 ;
        RECT 8.990 -81.410 9.450 -80.960 ;
        RECT 9.890 -81.410 10.350 -80.960 ;
        RECT 13.950 -81.100 14.410 -80.650 ;
        RECT 14.850 -81.100 15.310 -80.650 ;
        RECT 18.910 -81.410 19.370 -80.960 ;
        RECT 19.810 -81.410 20.270 -80.960 ;
        RECT 23.870 -81.100 24.330 -80.650 ;
        RECT -294.430 -175.680 -293.970 -175.230 ;
        RECT -290.370 -175.990 -289.910 -175.540 ;
        RECT -289.470 -175.990 -289.010 -175.540 ;
        RECT -285.410 -175.680 -284.950 -175.230 ;
        RECT -284.510 -175.680 -284.050 -175.230 ;
        RECT -280.450 -175.990 -279.990 -175.540 ;
        RECT -279.550 -175.990 -279.090 -175.540 ;
        RECT -275.490 -175.680 -275.030 -175.230 ;
        RECT -274.590 -175.680 -274.130 -175.230 ;
        RECT -270.530 -175.990 -270.070 -175.540 ;
        RECT -269.630 -175.990 -269.170 -175.540 ;
        RECT -265.570 -175.680 -265.110 -175.230 ;
        RECT -264.670 -175.680 -264.210 -175.230 ;
        RECT -260.610 -175.990 -260.150 -175.540 ;
        RECT -259.710 -175.990 -259.250 -175.540 ;
        RECT -255.650 -175.680 -255.190 -175.230 ;
        RECT -254.750 -175.680 -254.290 -175.230 ;
        RECT -250.690 -175.990 -250.230 -175.540 ;
        RECT -249.790 -175.990 -249.330 -175.540 ;
        RECT -245.730 -175.680 -245.270 -175.230 ;
        RECT -244.830 -175.680 -244.370 -175.230 ;
        RECT -240.770 -175.990 -240.310 -175.540 ;
        RECT -239.870 -175.990 -239.410 -175.540 ;
        RECT -235.810 -175.680 -235.350 -175.230 ;
        RECT -234.910 -175.680 -234.450 -175.230 ;
        RECT -230.850 -175.990 -230.390 -175.540 ;
        RECT -229.950 -175.990 -229.490 -175.540 ;
        RECT -225.890 -175.680 -225.430 -175.230 ;
        RECT -224.990 -175.680 -224.530 -175.230 ;
        RECT -220.930 -175.990 -220.470 -175.540 ;
        RECT -220.030 -175.990 -219.570 -175.540 ;
        RECT -215.970 -175.680 -215.510 -175.230 ;
        RECT -215.070 -175.680 -214.610 -175.230 ;
        RECT -211.010 -175.990 -210.550 -175.540 ;
        RECT -210.110 -175.990 -209.650 -175.540 ;
        RECT -206.050 -175.680 -205.590 -175.230 ;
        RECT -205.150 -175.680 -204.690 -175.230 ;
        RECT -201.090 -175.990 -200.630 -175.540 ;
        RECT -200.190 -175.990 -199.730 -175.540 ;
        RECT -196.130 -175.680 -195.670 -175.230 ;
        RECT -195.230 -175.680 -194.770 -175.230 ;
        RECT -191.170 -175.990 -190.710 -175.540 ;
        RECT -190.270 -175.990 -189.810 -175.540 ;
        RECT -186.210 -175.680 -185.750 -175.230 ;
        RECT -185.310 -175.680 -184.850 -175.230 ;
        RECT -181.250 -175.990 -180.790 -175.540 ;
        RECT -180.350 -175.990 -179.890 -175.540 ;
        RECT -176.290 -175.680 -175.830 -175.230 ;
        RECT -175.390 -175.680 -174.930 -175.230 ;
        RECT -171.330 -175.990 -170.870 -175.540 ;
        RECT -170.430 -175.990 -169.970 -175.540 ;
        RECT -166.370 -175.680 -165.910 -175.230 ;
        RECT -165.470 -175.680 -165.010 -175.230 ;
        RECT -161.410 -175.990 -160.950 -175.540 ;
        RECT -160.510 -175.990 -160.050 -175.540 ;
        RECT -156.450 -175.680 -155.990 -175.230 ;
        RECT -155.550 -175.680 -155.090 -175.230 ;
        RECT -151.490 -175.990 -151.030 -175.540 ;
        RECT -150.590 -175.990 -150.130 -175.540 ;
        RECT -146.530 -175.680 -146.070 -175.230 ;
        RECT -145.630 -175.680 -145.170 -175.230 ;
        RECT -141.570 -175.990 -141.110 -175.540 ;
        RECT -140.670 -175.990 -140.210 -175.540 ;
        RECT -136.610 -175.680 -136.150 -175.230 ;
        RECT -135.710 -175.680 -135.250 -175.230 ;
        RECT -131.650 -175.990 -131.190 -175.540 ;
        RECT -130.750 -175.990 -130.290 -175.540 ;
        RECT -126.690 -175.680 -126.230 -175.230 ;
        RECT -125.790 -175.680 -125.330 -175.230 ;
        RECT -121.730 -175.990 -121.270 -175.540 ;
        RECT -120.830 -175.990 -120.370 -175.540 ;
        RECT -116.770 -175.680 -116.310 -175.230 ;
        RECT -115.870 -175.680 -115.410 -175.230 ;
        RECT -111.810 -175.990 -111.350 -175.540 ;
        RECT -110.910 -175.990 -110.450 -175.540 ;
        RECT -106.850 -175.680 -106.390 -175.230 ;
        RECT -105.950 -175.680 -105.490 -175.230 ;
        RECT -101.890 -175.990 -101.430 -175.540 ;
        RECT -100.990 -175.990 -100.530 -175.540 ;
        RECT -96.930 -175.680 -96.470 -175.230 ;
        RECT -96.030 -175.680 -95.570 -175.230 ;
        RECT -91.970 -175.990 -91.510 -175.540 ;
        RECT -91.070 -175.990 -90.610 -175.540 ;
        RECT -87.010 -175.680 -86.550 -175.230 ;
        RECT -86.110 -175.680 -85.650 -175.230 ;
        RECT -82.050 -175.990 -81.590 -175.540 ;
        RECT -81.150 -175.990 -80.690 -175.540 ;
        RECT -77.090 -175.680 -76.630 -175.230 ;
        RECT -76.190 -175.680 -75.730 -175.230 ;
        RECT -72.130 -175.990 -71.670 -175.540 ;
        RECT -71.230 -175.990 -70.770 -175.540 ;
        RECT -67.170 -175.680 -66.710 -175.230 ;
        RECT -66.270 -175.680 -65.810 -175.230 ;
        RECT -62.210 -175.990 -61.750 -175.540 ;
        RECT -61.310 -175.990 -60.850 -175.540 ;
        RECT -57.250 -175.680 -56.790 -175.230 ;
        RECT -56.350 -175.680 -55.890 -175.230 ;
        RECT -52.290 -175.990 -51.830 -175.540 ;
        RECT -51.390 -175.990 -50.930 -175.540 ;
        RECT -47.330 -175.680 -46.870 -175.230 ;
        RECT -46.430 -175.680 -45.970 -175.230 ;
        RECT -42.370 -175.990 -41.910 -175.540 ;
        RECT -41.470 -175.990 -41.010 -175.540 ;
        RECT -37.410 -175.680 -36.950 -175.230 ;
        RECT -36.510 -175.680 -36.050 -175.230 ;
        RECT -32.450 -175.990 -31.990 -175.540 ;
        RECT -31.550 -175.990 -31.090 -175.540 ;
        RECT -27.490 -175.680 -27.030 -175.230 ;
        RECT -26.590 -175.680 -26.130 -175.230 ;
        RECT -22.530 -175.990 -22.070 -175.540 ;
        RECT -21.630 -175.990 -21.170 -175.540 ;
        RECT -17.570 -175.680 -17.110 -175.230 ;
        RECT -16.670 -175.680 -16.210 -175.230 ;
        RECT -12.610 -175.990 -12.150 -175.540 ;
        RECT -11.710 -175.990 -11.250 -175.540 ;
        RECT -7.650 -175.680 -7.190 -175.230 ;
        RECT -6.750 -175.680 -6.290 -175.230 ;
        RECT -2.690 -175.990 -2.230 -175.540 ;
        RECT -1.790 -175.990 -1.330 -175.540 ;
        RECT 2.270 -175.680 2.730 -175.230 ;
        RECT 3.170 -175.680 3.630 -175.230 ;
        RECT 7.230 -175.990 7.690 -175.540 ;
        RECT 8.130 -175.990 8.590 -175.540 ;
        RECT 12.190 -175.680 12.650 -175.230 ;
        RECT 13.090 -175.680 13.550 -175.230 ;
        RECT 17.150 -175.990 17.610 -175.540 ;
        RECT 18.050 -175.990 18.510 -175.540 ;
        RECT 22.110 -175.680 22.570 -175.230 ;
      LAYER via ;
        RECT -290.940 92.000 -290.640 92.300 ;
        RECT -286.860 91.640 -286.560 91.940 ;
        RECT -285.980 91.640 -285.680 91.940 ;
        RECT -281.900 92.000 -281.600 92.300 ;
        RECT -281.020 92.000 -280.720 92.300 ;
        RECT -276.940 91.640 -276.640 91.940 ;
        RECT -276.060 91.640 -275.760 91.940 ;
        RECT -271.980 92.000 -271.680 92.300 ;
        RECT -271.100 92.000 -270.800 92.300 ;
        RECT -267.020 91.640 -266.720 91.940 ;
        RECT -266.140 91.640 -265.840 91.940 ;
        RECT -262.060 92.000 -261.760 92.300 ;
        RECT -261.180 92.000 -260.880 92.300 ;
        RECT -257.100 91.640 -256.800 91.940 ;
        RECT -256.220 91.640 -255.920 91.940 ;
        RECT -252.140 92.000 -251.840 92.300 ;
        RECT -251.260 92.000 -250.960 92.300 ;
        RECT -247.180 91.640 -246.880 91.940 ;
        RECT -246.300 91.640 -246.000 91.940 ;
        RECT -242.220 92.000 -241.920 92.300 ;
        RECT -241.340 92.000 -241.040 92.300 ;
        RECT -237.260 91.640 -236.960 91.940 ;
        RECT -236.380 91.640 -236.080 91.940 ;
        RECT -232.300 92.000 -232.000 92.300 ;
        RECT -231.420 92.000 -231.120 92.300 ;
        RECT -227.340 91.640 -227.040 91.940 ;
        RECT -226.460 91.640 -226.160 91.940 ;
        RECT -222.380 92.000 -222.080 92.300 ;
        RECT -221.500 92.000 -221.200 92.300 ;
        RECT -217.420 91.640 -217.120 91.940 ;
        RECT -216.540 91.640 -216.240 91.940 ;
        RECT -212.460 92.000 -212.160 92.300 ;
        RECT -211.580 92.000 -211.280 92.300 ;
        RECT -207.500 91.640 -207.200 91.940 ;
        RECT -206.620 91.640 -206.320 91.940 ;
        RECT -202.540 92.000 -202.240 92.300 ;
        RECT -201.660 92.000 -201.360 92.300 ;
        RECT -197.580 91.640 -197.280 91.940 ;
        RECT -196.700 91.640 -196.400 91.940 ;
        RECT -192.620 92.000 -192.320 92.300 ;
        RECT -191.740 92.000 -191.440 92.300 ;
        RECT -187.660 91.640 -187.360 91.940 ;
        RECT -186.780 91.640 -186.480 91.940 ;
        RECT -182.700 92.000 -182.400 92.300 ;
        RECT -181.820 92.000 -181.520 92.300 ;
        RECT -177.740 91.640 -177.440 91.940 ;
        RECT -176.860 91.640 -176.560 91.940 ;
        RECT -172.780 92.000 -172.480 92.300 ;
        RECT -171.900 92.000 -171.600 92.300 ;
        RECT -167.820 91.640 -167.520 91.940 ;
        RECT -166.940 91.640 -166.640 91.940 ;
        RECT -162.860 92.000 -162.560 92.300 ;
        RECT -161.980 92.000 -161.680 92.300 ;
        RECT -157.900 91.640 -157.600 91.940 ;
        RECT -157.020 91.640 -156.720 91.940 ;
        RECT -152.940 92.000 -152.640 92.300 ;
        RECT -152.060 92.000 -151.760 92.300 ;
        RECT -147.980 91.640 -147.680 91.940 ;
        RECT -147.100 91.640 -146.800 91.940 ;
        RECT -143.020 92.000 -142.720 92.300 ;
        RECT -142.140 92.000 -141.840 92.300 ;
        RECT -138.060 91.640 -137.760 91.940 ;
        RECT -137.180 91.640 -136.880 91.940 ;
        RECT -133.100 92.000 -132.800 92.300 ;
        RECT -132.220 92.000 -131.920 92.300 ;
        RECT -128.140 91.640 -127.840 91.940 ;
        RECT -127.260 91.640 -126.960 91.940 ;
        RECT -123.180 92.000 -122.880 92.300 ;
        RECT -122.300 92.000 -122.000 92.300 ;
        RECT -118.220 91.640 -117.920 91.940 ;
        RECT -117.340 91.640 -117.040 91.940 ;
        RECT -113.260 92.000 -112.960 92.300 ;
        RECT -112.380 92.000 -112.080 92.300 ;
        RECT -108.300 91.640 -108.000 91.940 ;
        RECT -107.420 91.640 -107.120 91.940 ;
        RECT -103.340 92.000 -103.040 92.300 ;
        RECT -102.460 92.000 -102.160 92.300 ;
        RECT -98.380 91.640 -98.080 91.940 ;
        RECT -97.500 91.640 -97.200 91.940 ;
        RECT -93.420 92.000 -93.120 92.300 ;
        RECT -92.540 92.000 -92.240 92.300 ;
        RECT -88.460 91.640 -88.160 91.940 ;
        RECT -87.580 91.640 -87.280 91.940 ;
        RECT -83.500 92.000 -83.200 92.300 ;
        RECT -82.620 92.000 -82.320 92.300 ;
        RECT -78.540 91.640 -78.240 91.940 ;
        RECT -77.660 91.640 -77.360 91.940 ;
        RECT -73.580 92.000 -73.280 92.300 ;
        RECT -72.700 92.000 -72.400 92.300 ;
        RECT -68.620 91.640 -68.320 91.940 ;
        RECT -67.740 91.640 -67.440 91.940 ;
        RECT -63.660 92.000 -63.360 92.300 ;
        RECT -62.780 92.000 -62.480 92.300 ;
        RECT -58.700 91.640 -58.400 91.940 ;
        RECT -57.820 91.640 -57.520 91.940 ;
        RECT -53.740 92.000 -53.440 92.300 ;
        RECT -52.860 92.000 -52.560 92.300 ;
        RECT -48.780 91.640 -48.480 91.940 ;
        RECT -47.900 91.640 -47.600 91.940 ;
        RECT -43.820 92.000 -43.520 92.300 ;
        RECT -42.940 92.000 -42.640 92.300 ;
        RECT -38.860 91.640 -38.560 91.940 ;
        RECT -37.980 91.640 -37.680 91.940 ;
        RECT -33.900 92.000 -33.600 92.300 ;
        RECT -33.020 92.000 -32.720 92.300 ;
        RECT -28.940 91.640 -28.640 91.940 ;
        RECT -28.060 91.640 -27.760 91.940 ;
        RECT -23.980 92.000 -23.680 92.300 ;
        RECT -23.100 92.000 -22.800 92.300 ;
        RECT -19.020 91.640 -18.720 91.940 ;
        RECT -18.140 91.640 -17.840 91.940 ;
        RECT -14.060 92.000 -13.760 92.300 ;
        RECT -13.180 92.000 -12.880 92.300 ;
        RECT -9.100 91.640 -8.800 91.940 ;
        RECT -8.220 91.640 -7.920 91.940 ;
        RECT -4.140 92.000 -3.840 92.300 ;
        RECT -3.260 92.000 -2.960 92.300 ;
        RECT 0.820 91.640 1.120 91.940 ;
        RECT 1.700 91.640 2.000 91.940 ;
        RECT 5.780 92.000 6.080 92.300 ;
        RECT 6.660 92.000 6.960 92.300 ;
        RECT 10.740 91.640 11.040 91.940 ;
        RECT 11.620 91.640 11.920 91.940 ;
        RECT 15.700 92.000 16.000 92.300 ;
        RECT 16.580 92.000 16.880 92.300 ;
        RECT 20.660 91.640 20.960 91.940 ;
        RECT 21.540 91.640 21.840 91.940 ;
        RECT 25.620 92.000 25.920 92.300 ;
        RECT -292.960 7.950 -292.660 8.250 ;
        RECT -288.880 7.590 -288.580 7.890 ;
        RECT -288.000 7.590 -287.700 7.890 ;
        RECT -283.920 7.950 -283.620 8.250 ;
        RECT -283.040 7.950 -282.740 8.250 ;
        RECT -278.960 7.590 -278.660 7.890 ;
        RECT -278.080 7.590 -277.780 7.890 ;
        RECT -274.000 7.950 -273.700 8.250 ;
        RECT -273.120 7.950 -272.820 8.250 ;
        RECT -269.040 7.590 -268.740 7.890 ;
        RECT -268.160 7.590 -267.860 7.890 ;
        RECT -264.080 7.950 -263.780 8.250 ;
        RECT -263.200 7.950 -262.900 8.250 ;
        RECT -259.120 7.590 -258.820 7.890 ;
        RECT -258.240 7.590 -257.940 7.890 ;
        RECT -254.160 7.950 -253.860 8.250 ;
        RECT -253.280 7.950 -252.980 8.250 ;
        RECT -249.200 7.590 -248.900 7.890 ;
        RECT -248.320 7.590 -248.020 7.890 ;
        RECT -244.240 7.950 -243.940 8.250 ;
        RECT -243.360 7.950 -243.060 8.250 ;
        RECT -239.280 7.590 -238.980 7.890 ;
        RECT -238.400 7.590 -238.100 7.890 ;
        RECT -234.320 7.950 -234.020 8.250 ;
        RECT -233.440 7.950 -233.140 8.250 ;
        RECT -229.360 7.590 -229.060 7.890 ;
        RECT -228.480 7.590 -228.180 7.890 ;
        RECT -224.400 7.950 -224.100 8.250 ;
        RECT -223.520 7.950 -223.220 8.250 ;
        RECT -219.440 7.590 -219.140 7.890 ;
        RECT -218.560 7.590 -218.260 7.890 ;
        RECT -214.480 7.950 -214.180 8.250 ;
        RECT -213.600 7.950 -213.300 8.250 ;
        RECT -209.520 7.590 -209.220 7.890 ;
        RECT -208.640 7.590 -208.340 7.890 ;
        RECT -204.560 7.950 -204.260 8.250 ;
        RECT -203.680 7.950 -203.380 8.250 ;
        RECT -199.600 7.590 -199.300 7.890 ;
        RECT -198.720 7.590 -198.420 7.890 ;
        RECT -194.640 7.950 -194.340 8.250 ;
        RECT -193.760 7.950 -193.460 8.250 ;
        RECT -189.680 7.590 -189.380 7.890 ;
        RECT -188.800 7.590 -188.500 7.890 ;
        RECT -184.720 7.950 -184.420 8.250 ;
        RECT -183.840 7.950 -183.540 8.250 ;
        RECT -179.760 7.590 -179.460 7.890 ;
        RECT -178.880 7.590 -178.580 7.890 ;
        RECT -174.800 7.950 -174.500 8.250 ;
        RECT -173.920 7.950 -173.620 8.250 ;
        RECT -169.840 7.590 -169.540 7.890 ;
        RECT -168.960 7.590 -168.660 7.890 ;
        RECT -164.880 7.950 -164.580 8.250 ;
        RECT -164.000 7.950 -163.700 8.250 ;
        RECT -159.920 7.590 -159.620 7.890 ;
        RECT -159.040 7.590 -158.740 7.890 ;
        RECT -154.960 7.950 -154.660 8.250 ;
        RECT -154.080 7.950 -153.780 8.250 ;
        RECT -150.000 7.590 -149.700 7.890 ;
        RECT -149.120 7.590 -148.820 7.890 ;
        RECT -145.040 7.950 -144.740 8.250 ;
        RECT -144.160 7.950 -143.860 8.250 ;
        RECT -140.080 7.590 -139.780 7.890 ;
        RECT -139.200 7.590 -138.900 7.890 ;
        RECT -135.120 7.950 -134.820 8.250 ;
        RECT -134.240 7.950 -133.940 8.250 ;
        RECT -130.160 7.590 -129.860 7.890 ;
        RECT -129.280 7.590 -128.980 7.890 ;
        RECT -125.200 7.950 -124.900 8.250 ;
        RECT -124.320 7.950 -124.020 8.250 ;
        RECT -120.240 7.590 -119.940 7.890 ;
        RECT -119.360 7.590 -119.060 7.890 ;
        RECT -115.280 7.950 -114.980 8.250 ;
        RECT -114.400 7.950 -114.100 8.250 ;
        RECT -110.320 7.590 -110.020 7.890 ;
        RECT -109.440 7.590 -109.140 7.890 ;
        RECT -105.360 7.950 -105.060 8.250 ;
        RECT -104.480 7.950 -104.180 8.250 ;
        RECT -100.400 7.590 -100.100 7.890 ;
        RECT -99.520 7.590 -99.220 7.890 ;
        RECT -95.440 7.950 -95.140 8.250 ;
        RECT -94.560 7.950 -94.260 8.250 ;
        RECT -90.480 7.590 -90.180 7.890 ;
        RECT -89.600 7.590 -89.300 7.890 ;
        RECT -85.520 7.950 -85.220 8.250 ;
        RECT -84.640 7.950 -84.340 8.250 ;
        RECT -80.560 7.590 -80.260 7.890 ;
        RECT -79.680 7.590 -79.380 7.890 ;
        RECT -75.600 7.950 -75.300 8.250 ;
        RECT -74.720 7.950 -74.420 8.250 ;
        RECT -70.640 7.590 -70.340 7.890 ;
        RECT -69.760 7.590 -69.460 7.890 ;
        RECT -65.680 7.950 -65.380 8.250 ;
        RECT -64.800 7.950 -64.500 8.250 ;
        RECT -60.720 7.590 -60.420 7.890 ;
        RECT -59.840 7.590 -59.540 7.890 ;
        RECT -55.760 7.950 -55.460 8.250 ;
        RECT -54.880 7.950 -54.580 8.250 ;
        RECT -50.800 7.590 -50.500 7.890 ;
        RECT -49.920 7.590 -49.620 7.890 ;
        RECT -45.840 7.950 -45.540 8.250 ;
        RECT -44.960 7.950 -44.660 8.250 ;
        RECT -40.880 7.590 -40.580 7.890 ;
        RECT -40.000 7.590 -39.700 7.890 ;
        RECT -35.920 7.950 -35.620 8.250 ;
        RECT -35.040 7.950 -34.740 8.250 ;
        RECT -30.960 7.590 -30.660 7.890 ;
        RECT -30.080 7.590 -29.780 7.890 ;
        RECT -26.000 7.950 -25.700 8.250 ;
        RECT -25.120 7.950 -24.820 8.250 ;
        RECT -21.040 7.590 -20.740 7.890 ;
        RECT -20.160 7.590 -19.860 7.890 ;
        RECT -16.080 7.950 -15.780 8.250 ;
        RECT -15.200 7.950 -14.900 8.250 ;
        RECT -11.120 7.590 -10.820 7.890 ;
        RECT -10.240 7.590 -9.940 7.890 ;
        RECT -6.160 7.950 -5.860 8.250 ;
        RECT -5.280 7.950 -4.980 8.250 ;
        RECT -1.200 7.590 -0.900 7.890 ;
        RECT -0.320 7.590 -0.020 7.890 ;
        RECT 3.760 7.950 4.060 8.250 ;
        RECT 4.640 7.950 4.940 8.250 ;
        RECT 8.720 7.590 9.020 7.890 ;
        RECT 9.600 7.590 9.900 7.890 ;
        RECT 13.680 7.950 13.980 8.250 ;
        RECT 14.560 7.950 14.860 8.250 ;
        RECT 18.640 7.590 18.940 7.890 ;
        RECT 19.520 7.590 19.820 7.890 ;
        RECT 23.600 7.950 23.900 8.250 ;
        RECT -292.600 -81.000 -292.300 -80.700 ;
        RECT -288.520 -81.360 -288.220 -81.060 ;
        RECT -287.640 -81.360 -287.340 -81.060 ;
        RECT -283.560 -81.000 -283.260 -80.700 ;
        RECT -282.680 -81.000 -282.380 -80.700 ;
        RECT -278.600 -81.360 -278.300 -81.060 ;
        RECT -277.720 -81.360 -277.420 -81.060 ;
        RECT -273.640 -81.000 -273.340 -80.700 ;
        RECT -272.760 -81.000 -272.460 -80.700 ;
        RECT -268.680 -81.360 -268.380 -81.060 ;
        RECT -267.800 -81.360 -267.500 -81.060 ;
        RECT -263.720 -81.000 -263.420 -80.700 ;
        RECT -262.840 -81.000 -262.540 -80.700 ;
        RECT -258.760 -81.360 -258.460 -81.060 ;
        RECT -257.880 -81.360 -257.580 -81.060 ;
        RECT -253.800 -81.000 -253.500 -80.700 ;
        RECT -252.920 -81.000 -252.620 -80.700 ;
        RECT -248.840 -81.360 -248.540 -81.060 ;
        RECT -247.960 -81.360 -247.660 -81.060 ;
        RECT -243.880 -81.000 -243.580 -80.700 ;
        RECT -243.000 -81.000 -242.700 -80.700 ;
        RECT -238.920 -81.360 -238.620 -81.060 ;
        RECT -238.040 -81.360 -237.740 -81.060 ;
        RECT -233.960 -81.000 -233.660 -80.700 ;
        RECT -233.080 -81.000 -232.780 -80.700 ;
        RECT -229.000 -81.360 -228.700 -81.060 ;
        RECT -228.120 -81.360 -227.820 -81.060 ;
        RECT -224.040 -81.000 -223.740 -80.700 ;
        RECT -223.160 -81.000 -222.860 -80.700 ;
        RECT -219.080 -81.360 -218.780 -81.060 ;
        RECT -218.200 -81.360 -217.900 -81.060 ;
        RECT -214.120 -81.000 -213.820 -80.700 ;
        RECT -213.240 -81.000 -212.940 -80.700 ;
        RECT -209.160 -81.360 -208.860 -81.060 ;
        RECT -208.280 -81.360 -207.980 -81.060 ;
        RECT -204.200 -81.000 -203.900 -80.700 ;
        RECT -203.320 -81.000 -203.020 -80.700 ;
        RECT -199.240 -81.360 -198.940 -81.060 ;
        RECT -198.360 -81.360 -198.060 -81.060 ;
        RECT -194.280 -81.000 -193.980 -80.700 ;
        RECT -193.400 -81.000 -193.100 -80.700 ;
        RECT -189.320 -81.360 -189.020 -81.060 ;
        RECT -188.440 -81.360 -188.140 -81.060 ;
        RECT -184.360 -81.000 -184.060 -80.700 ;
        RECT -183.480 -81.000 -183.180 -80.700 ;
        RECT -179.400 -81.360 -179.100 -81.060 ;
        RECT -178.520 -81.360 -178.220 -81.060 ;
        RECT -174.440 -81.000 -174.140 -80.700 ;
        RECT -173.560 -81.000 -173.260 -80.700 ;
        RECT -169.480 -81.360 -169.180 -81.060 ;
        RECT -168.600 -81.360 -168.300 -81.060 ;
        RECT -164.520 -81.000 -164.220 -80.700 ;
        RECT -163.640 -81.000 -163.340 -80.700 ;
        RECT -159.560 -81.360 -159.260 -81.060 ;
        RECT -158.680 -81.360 -158.380 -81.060 ;
        RECT -154.600 -81.000 -154.300 -80.700 ;
        RECT -153.720 -81.000 -153.420 -80.700 ;
        RECT -149.640 -81.360 -149.340 -81.060 ;
        RECT -148.760 -81.360 -148.460 -81.060 ;
        RECT -144.680 -81.000 -144.380 -80.700 ;
        RECT -143.800 -81.000 -143.500 -80.700 ;
        RECT -139.720 -81.360 -139.420 -81.060 ;
        RECT -138.840 -81.360 -138.540 -81.060 ;
        RECT -134.760 -81.000 -134.460 -80.700 ;
        RECT -133.880 -81.000 -133.580 -80.700 ;
        RECT -129.800 -81.360 -129.500 -81.060 ;
        RECT -128.920 -81.360 -128.620 -81.060 ;
        RECT -124.840 -81.000 -124.540 -80.700 ;
        RECT -123.960 -81.000 -123.660 -80.700 ;
        RECT -119.880 -81.360 -119.580 -81.060 ;
        RECT -119.000 -81.360 -118.700 -81.060 ;
        RECT -114.920 -81.000 -114.620 -80.700 ;
        RECT -114.040 -81.000 -113.740 -80.700 ;
        RECT -109.960 -81.360 -109.660 -81.060 ;
        RECT -109.080 -81.360 -108.780 -81.060 ;
        RECT -105.000 -81.000 -104.700 -80.700 ;
        RECT -104.120 -81.000 -103.820 -80.700 ;
        RECT -100.040 -81.360 -99.740 -81.060 ;
        RECT -99.160 -81.360 -98.860 -81.060 ;
        RECT -95.080 -81.000 -94.780 -80.700 ;
        RECT -94.200 -81.000 -93.900 -80.700 ;
        RECT -90.120 -81.360 -89.820 -81.060 ;
        RECT -89.240 -81.360 -88.940 -81.060 ;
        RECT -85.160 -81.000 -84.860 -80.700 ;
        RECT -84.280 -81.000 -83.980 -80.700 ;
        RECT -80.200 -81.360 -79.900 -81.060 ;
        RECT -79.320 -81.360 -79.020 -81.060 ;
        RECT -75.240 -81.000 -74.940 -80.700 ;
        RECT -74.360 -81.000 -74.060 -80.700 ;
        RECT -70.280 -81.360 -69.980 -81.060 ;
        RECT -69.400 -81.360 -69.100 -81.060 ;
        RECT -65.320 -81.000 -65.020 -80.700 ;
        RECT -64.440 -81.000 -64.140 -80.700 ;
        RECT -60.360 -81.360 -60.060 -81.060 ;
        RECT -59.480 -81.360 -59.180 -81.060 ;
        RECT -55.400 -81.000 -55.100 -80.700 ;
        RECT -54.520 -81.000 -54.220 -80.700 ;
        RECT -50.440 -81.360 -50.140 -81.060 ;
        RECT -49.560 -81.360 -49.260 -81.060 ;
        RECT -45.480 -81.000 -45.180 -80.700 ;
        RECT -44.600 -81.000 -44.300 -80.700 ;
        RECT -40.520 -81.360 -40.220 -81.060 ;
        RECT -39.640 -81.360 -39.340 -81.060 ;
        RECT -35.560 -81.000 -35.260 -80.700 ;
        RECT -34.680 -81.000 -34.380 -80.700 ;
        RECT -30.600 -81.360 -30.300 -81.060 ;
        RECT -29.720 -81.360 -29.420 -81.060 ;
        RECT -25.640 -81.000 -25.340 -80.700 ;
        RECT -24.760 -81.000 -24.460 -80.700 ;
        RECT -20.680 -81.360 -20.380 -81.060 ;
        RECT -19.800 -81.360 -19.500 -81.060 ;
        RECT -15.720 -81.000 -15.420 -80.700 ;
        RECT -14.840 -81.000 -14.540 -80.700 ;
        RECT -10.760 -81.360 -10.460 -81.060 ;
        RECT -9.880 -81.360 -9.580 -81.060 ;
        RECT -5.800 -81.000 -5.500 -80.700 ;
        RECT -4.920 -81.000 -4.620 -80.700 ;
        RECT -0.840 -81.360 -0.540 -81.060 ;
        RECT 0.040 -81.360 0.340 -81.060 ;
        RECT 4.120 -81.000 4.420 -80.700 ;
        RECT 5.000 -81.000 5.300 -80.700 ;
        RECT 9.080 -81.360 9.380 -81.060 ;
        RECT 9.960 -81.360 10.260 -81.060 ;
        RECT 14.040 -81.000 14.340 -80.700 ;
        RECT 14.920 -81.000 15.220 -80.700 ;
        RECT 19.000 -81.360 19.300 -81.060 ;
        RECT 19.880 -81.360 20.180 -81.060 ;
        RECT 23.960 -81.000 24.260 -80.700 ;
        RECT -294.360 -175.580 -294.060 -175.280 ;
        RECT -290.280 -175.940 -289.980 -175.640 ;
        RECT -289.400 -175.940 -289.100 -175.640 ;
        RECT -285.320 -175.580 -285.020 -175.280 ;
        RECT -284.440 -175.580 -284.140 -175.280 ;
        RECT -280.360 -175.940 -280.060 -175.640 ;
        RECT -279.480 -175.940 -279.180 -175.640 ;
        RECT -275.400 -175.580 -275.100 -175.280 ;
        RECT -274.520 -175.580 -274.220 -175.280 ;
        RECT -270.440 -175.940 -270.140 -175.640 ;
        RECT -269.560 -175.940 -269.260 -175.640 ;
        RECT -265.480 -175.580 -265.180 -175.280 ;
        RECT -264.600 -175.580 -264.300 -175.280 ;
        RECT -260.520 -175.940 -260.220 -175.640 ;
        RECT -259.640 -175.940 -259.340 -175.640 ;
        RECT -255.560 -175.580 -255.260 -175.280 ;
        RECT -254.680 -175.580 -254.380 -175.280 ;
        RECT -250.600 -175.940 -250.300 -175.640 ;
        RECT -249.720 -175.940 -249.420 -175.640 ;
        RECT -245.640 -175.580 -245.340 -175.280 ;
        RECT -244.760 -175.580 -244.460 -175.280 ;
        RECT -240.680 -175.940 -240.380 -175.640 ;
        RECT -239.800 -175.940 -239.500 -175.640 ;
        RECT -235.720 -175.580 -235.420 -175.280 ;
        RECT -234.840 -175.580 -234.540 -175.280 ;
        RECT -230.760 -175.940 -230.460 -175.640 ;
        RECT -229.880 -175.940 -229.580 -175.640 ;
        RECT -225.800 -175.580 -225.500 -175.280 ;
        RECT -224.920 -175.580 -224.620 -175.280 ;
        RECT -220.840 -175.940 -220.540 -175.640 ;
        RECT -219.960 -175.940 -219.660 -175.640 ;
        RECT -215.880 -175.580 -215.580 -175.280 ;
        RECT -215.000 -175.580 -214.700 -175.280 ;
        RECT -210.920 -175.940 -210.620 -175.640 ;
        RECT -210.040 -175.940 -209.740 -175.640 ;
        RECT -205.960 -175.580 -205.660 -175.280 ;
        RECT -205.080 -175.580 -204.780 -175.280 ;
        RECT -201.000 -175.940 -200.700 -175.640 ;
        RECT -200.120 -175.940 -199.820 -175.640 ;
        RECT -196.040 -175.580 -195.740 -175.280 ;
        RECT -195.160 -175.580 -194.860 -175.280 ;
        RECT -191.080 -175.940 -190.780 -175.640 ;
        RECT -190.200 -175.940 -189.900 -175.640 ;
        RECT -186.120 -175.580 -185.820 -175.280 ;
        RECT -185.240 -175.580 -184.940 -175.280 ;
        RECT -181.160 -175.940 -180.860 -175.640 ;
        RECT -180.280 -175.940 -179.980 -175.640 ;
        RECT -176.200 -175.580 -175.900 -175.280 ;
        RECT -175.320 -175.580 -175.020 -175.280 ;
        RECT -171.240 -175.940 -170.940 -175.640 ;
        RECT -170.360 -175.940 -170.060 -175.640 ;
        RECT -166.280 -175.580 -165.980 -175.280 ;
        RECT -165.400 -175.580 -165.100 -175.280 ;
        RECT -161.320 -175.940 -161.020 -175.640 ;
        RECT -160.440 -175.940 -160.140 -175.640 ;
        RECT -156.360 -175.580 -156.060 -175.280 ;
        RECT -155.480 -175.580 -155.180 -175.280 ;
        RECT -151.400 -175.940 -151.100 -175.640 ;
        RECT -150.520 -175.940 -150.220 -175.640 ;
        RECT -146.440 -175.580 -146.140 -175.280 ;
        RECT -145.560 -175.580 -145.260 -175.280 ;
        RECT -141.480 -175.940 -141.180 -175.640 ;
        RECT -140.600 -175.940 -140.300 -175.640 ;
        RECT -136.520 -175.580 -136.220 -175.280 ;
        RECT -135.640 -175.580 -135.340 -175.280 ;
        RECT -131.560 -175.940 -131.260 -175.640 ;
        RECT -130.680 -175.940 -130.380 -175.640 ;
        RECT -126.600 -175.580 -126.300 -175.280 ;
        RECT -125.720 -175.580 -125.420 -175.280 ;
        RECT -121.640 -175.940 -121.340 -175.640 ;
        RECT -120.760 -175.940 -120.460 -175.640 ;
        RECT -116.680 -175.580 -116.380 -175.280 ;
        RECT -115.800 -175.580 -115.500 -175.280 ;
        RECT -111.720 -175.940 -111.420 -175.640 ;
        RECT -110.840 -175.940 -110.540 -175.640 ;
        RECT -106.760 -175.580 -106.460 -175.280 ;
        RECT -105.880 -175.580 -105.580 -175.280 ;
        RECT -101.800 -175.940 -101.500 -175.640 ;
        RECT -100.920 -175.940 -100.620 -175.640 ;
        RECT -96.840 -175.580 -96.540 -175.280 ;
        RECT -95.960 -175.580 -95.660 -175.280 ;
        RECT -91.880 -175.940 -91.580 -175.640 ;
        RECT -91.000 -175.940 -90.700 -175.640 ;
        RECT -86.920 -175.580 -86.620 -175.280 ;
        RECT -86.040 -175.580 -85.740 -175.280 ;
        RECT -81.960 -175.940 -81.660 -175.640 ;
        RECT -81.080 -175.940 -80.780 -175.640 ;
        RECT -77.000 -175.580 -76.700 -175.280 ;
        RECT -76.120 -175.580 -75.820 -175.280 ;
        RECT -72.040 -175.940 -71.740 -175.640 ;
        RECT -71.160 -175.940 -70.860 -175.640 ;
        RECT -67.080 -175.580 -66.780 -175.280 ;
        RECT -66.200 -175.580 -65.900 -175.280 ;
        RECT -62.120 -175.940 -61.820 -175.640 ;
        RECT -61.240 -175.940 -60.940 -175.640 ;
        RECT -57.160 -175.580 -56.860 -175.280 ;
        RECT -56.280 -175.580 -55.980 -175.280 ;
        RECT -52.200 -175.940 -51.900 -175.640 ;
        RECT -51.320 -175.940 -51.020 -175.640 ;
        RECT -47.240 -175.580 -46.940 -175.280 ;
        RECT -46.360 -175.580 -46.060 -175.280 ;
        RECT -42.280 -175.940 -41.980 -175.640 ;
        RECT -41.400 -175.940 -41.100 -175.640 ;
        RECT -37.320 -175.580 -37.020 -175.280 ;
        RECT -36.440 -175.580 -36.140 -175.280 ;
        RECT -32.360 -175.940 -32.060 -175.640 ;
        RECT -31.480 -175.940 -31.180 -175.640 ;
        RECT -27.400 -175.580 -27.100 -175.280 ;
        RECT -26.520 -175.580 -26.220 -175.280 ;
        RECT -22.440 -175.940 -22.140 -175.640 ;
        RECT -21.560 -175.940 -21.260 -175.640 ;
        RECT -17.480 -175.580 -17.180 -175.280 ;
        RECT -16.600 -175.580 -16.300 -175.280 ;
        RECT -12.520 -175.940 -12.220 -175.640 ;
        RECT -11.640 -175.940 -11.340 -175.640 ;
        RECT -7.560 -175.580 -7.260 -175.280 ;
        RECT -6.680 -175.580 -6.380 -175.280 ;
        RECT -2.600 -175.940 -2.300 -175.640 ;
        RECT -1.720 -175.940 -1.420 -175.640 ;
        RECT 2.360 -175.580 2.660 -175.280 ;
        RECT 3.240 -175.580 3.540 -175.280 ;
        RECT 7.320 -175.940 7.620 -175.640 ;
        RECT 8.200 -175.940 8.500 -175.640 ;
        RECT 12.280 -175.580 12.580 -175.280 ;
        RECT 13.160 -175.580 13.460 -175.280 ;
        RECT 17.240 -175.940 17.540 -175.640 ;
        RECT 18.120 -175.940 18.420 -175.640 ;
        RECT 22.200 -175.580 22.500 -175.280 ;
      LAYER met2 ;
        RECT -291.010 92.040 -290.550 92.350 ;
        RECT -288.820 92.040 -288.680 92.440 ;
        RECT -283.860 92.040 -283.720 92.440 ;
        RECT -281.990 92.040 -280.630 92.350 ;
        RECT -278.900 92.040 -278.760 92.440 ;
        RECT -273.940 92.040 -273.800 92.440 ;
        RECT -272.070 92.040 -270.710 92.350 ;
        RECT -268.980 92.040 -268.840 92.440 ;
        RECT -264.020 92.040 -263.880 92.440 ;
        RECT -262.150 92.040 -260.790 92.350 ;
        RECT -259.060 92.040 -258.920 92.440 ;
        RECT -254.100 92.040 -253.960 92.440 ;
        RECT -252.230 92.040 -250.870 92.350 ;
        RECT -249.140 92.040 -249.000 92.440 ;
        RECT -244.180 92.040 -244.040 92.440 ;
        RECT -242.310 92.040 -240.950 92.350 ;
        RECT -239.220 92.040 -239.080 92.440 ;
        RECT -234.260 92.040 -234.120 92.440 ;
        RECT -232.390 92.040 -231.030 92.350 ;
        RECT -229.300 92.040 -229.160 92.440 ;
        RECT -224.340 92.040 -224.200 92.440 ;
        RECT -222.470 92.040 -221.110 92.350 ;
        RECT -219.380 92.040 -219.240 92.440 ;
        RECT -214.420 92.040 -214.280 92.440 ;
        RECT -212.550 92.040 -211.190 92.350 ;
        RECT -209.460 92.040 -209.320 92.440 ;
        RECT -204.500 92.040 -204.360 92.440 ;
        RECT -202.630 92.040 -201.270 92.350 ;
        RECT -199.540 92.040 -199.400 92.440 ;
        RECT -194.580 92.040 -194.440 92.440 ;
        RECT -192.710 92.040 -191.350 92.350 ;
        RECT -189.620 92.040 -189.480 92.440 ;
        RECT -184.660 92.040 -184.520 92.440 ;
        RECT -182.790 92.040 -181.430 92.350 ;
        RECT -179.700 92.040 -179.560 92.440 ;
        RECT -174.740 92.040 -174.600 92.440 ;
        RECT -172.870 92.040 -171.510 92.350 ;
        RECT -169.780 92.040 -169.640 92.440 ;
        RECT -164.820 92.040 -164.680 92.440 ;
        RECT -162.950 92.040 -161.590 92.350 ;
        RECT -159.860 92.040 -159.720 92.440 ;
        RECT -154.900 92.040 -154.760 92.440 ;
        RECT -153.030 92.040 -151.670 92.350 ;
        RECT -149.940 92.040 -149.800 92.440 ;
        RECT -144.980 92.040 -144.840 92.440 ;
        RECT -143.110 92.040 -141.750 92.350 ;
        RECT -140.020 92.040 -139.880 92.440 ;
        RECT -135.060 92.040 -134.920 92.440 ;
        RECT -133.190 92.040 -131.830 92.350 ;
        RECT -130.100 92.040 -129.960 92.440 ;
        RECT -125.140 92.040 -125.000 92.440 ;
        RECT -123.270 92.040 -121.910 92.350 ;
        RECT -120.180 92.040 -120.040 92.440 ;
        RECT -115.220 92.040 -115.080 92.440 ;
        RECT -113.350 92.040 -111.990 92.350 ;
        RECT -110.260 92.040 -110.120 92.440 ;
        RECT -105.300 92.040 -105.160 92.440 ;
        RECT -103.430 92.040 -102.070 92.350 ;
        RECT -100.340 92.040 -100.200 92.440 ;
        RECT -95.380 92.040 -95.240 92.440 ;
        RECT -93.510 92.040 -92.150 92.350 ;
        RECT -90.420 92.040 -90.280 92.440 ;
        RECT -85.460 92.040 -85.320 92.440 ;
        RECT -83.590 92.040 -82.230 92.350 ;
        RECT -80.500 92.040 -80.360 92.440 ;
        RECT -75.540 92.040 -75.400 92.440 ;
        RECT -73.670 92.040 -72.310 92.350 ;
        RECT -70.580 92.040 -70.440 92.440 ;
        RECT -65.620 92.040 -65.480 92.440 ;
        RECT -63.750 92.040 -62.390 92.350 ;
        RECT -60.660 92.040 -60.520 92.440 ;
        RECT -55.700 92.040 -55.560 92.440 ;
        RECT -53.830 92.040 -52.470 92.350 ;
        RECT -50.740 92.040 -50.600 92.440 ;
        RECT -45.780 92.040 -45.640 92.440 ;
        RECT -43.910 92.040 -42.550 92.350 ;
        RECT -40.820 92.040 -40.680 92.440 ;
        RECT -35.860 92.040 -35.720 92.440 ;
        RECT -33.990 92.040 -32.630 92.350 ;
        RECT -30.900 92.040 -30.760 92.440 ;
        RECT -25.940 92.040 -25.800 92.440 ;
        RECT -24.070 92.040 -22.710 92.350 ;
        RECT -20.980 92.040 -20.840 92.440 ;
        RECT -16.020 92.040 -15.880 92.440 ;
        RECT -14.150 92.040 -12.790 92.350 ;
        RECT -11.060 92.040 -10.920 92.440 ;
        RECT -6.100 92.040 -5.960 92.440 ;
        RECT -4.230 92.040 -2.870 92.350 ;
        RECT -1.140 92.040 -1.000 92.440 ;
        RECT 3.820 92.040 3.960 92.440 ;
        RECT 5.690 92.040 7.050 92.350 ;
        RECT 8.780 92.040 8.920 92.440 ;
        RECT 13.740 92.040 13.880 92.440 ;
        RECT 15.610 92.040 16.970 92.350 ;
        RECT 18.700 92.040 18.840 92.440 ;
        RECT 23.660 92.040 23.800 92.440 ;
        RECT 37.260 92.370 37.720 96.680 ;
        RECT 32.950 92.360 37.720 92.370 ;
        RECT 25.530 92.040 37.720 92.360 ;
        RECT -291.010 91.910 37.720 92.040 ;
        RECT -291.010 91.900 34.270 91.910 ;
        RECT -288.820 91.500 -288.680 91.900 ;
        RECT -286.950 91.590 -285.590 91.900 ;
        RECT -283.860 91.500 -283.720 91.900 ;
        RECT -278.900 91.500 -278.760 91.900 ;
        RECT -277.030 91.590 -275.670 91.900 ;
        RECT -273.940 91.500 -273.800 91.900 ;
        RECT -268.980 91.500 -268.840 91.900 ;
        RECT -267.110 91.590 -265.750 91.900 ;
        RECT -264.020 91.500 -263.880 91.900 ;
        RECT -259.060 91.500 -258.920 91.900 ;
        RECT -257.190 91.590 -255.830 91.900 ;
        RECT -254.100 91.500 -253.960 91.900 ;
        RECT -249.140 91.500 -249.000 91.900 ;
        RECT -247.270 91.590 -245.910 91.900 ;
        RECT -244.180 91.500 -244.040 91.900 ;
        RECT -239.220 91.500 -239.080 91.900 ;
        RECT -237.350 91.590 -235.990 91.900 ;
        RECT -234.260 91.500 -234.120 91.900 ;
        RECT -229.300 91.500 -229.160 91.900 ;
        RECT -227.430 91.590 -226.070 91.900 ;
        RECT -224.340 91.500 -224.200 91.900 ;
        RECT -219.380 91.500 -219.240 91.900 ;
        RECT -217.510 91.590 -216.150 91.900 ;
        RECT -214.420 91.500 -214.280 91.900 ;
        RECT -209.460 91.500 -209.320 91.900 ;
        RECT -207.590 91.590 -206.230 91.900 ;
        RECT -204.500 91.500 -204.360 91.900 ;
        RECT -199.540 91.500 -199.400 91.900 ;
        RECT -197.670 91.590 -196.310 91.900 ;
        RECT -194.580 91.500 -194.440 91.900 ;
        RECT -189.620 91.500 -189.480 91.900 ;
        RECT -187.750 91.590 -186.390 91.900 ;
        RECT -184.660 91.500 -184.520 91.900 ;
        RECT -179.700 91.500 -179.560 91.900 ;
        RECT -177.830 91.590 -176.470 91.900 ;
        RECT -174.740 91.500 -174.600 91.900 ;
        RECT -169.780 91.500 -169.640 91.900 ;
        RECT -167.910 91.590 -166.550 91.900 ;
        RECT -164.820 91.500 -164.680 91.900 ;
        RECT -159.860 91.500 -159.720 91.900 ;
        RECT -157.990 91.590 -156.630 91.900 ;
        RECT -154.900 91.500 -154.760 91.900 ;
        RECT -149.940 91.500 -149.800 91.900 ;
        RECT -148.070 91.590 -146.710 91.900 ;
        RECT -144.980 91.500 -144.840 91.900 ;
        RECT -140.020 91.500 -139.880 91.900 ;
        RECT -138.150 91.590 -136.790 91.900 ;
        RECT -135.060 91.500 -134.920 91.900 ;
        RECT -130.100 91.500 -129.960 91.900 ;
        RECT -128.230 91.590 -126.870 91.900 ;
        RECT -125.140 91.500 -125.000 91.900 ;
        RECT -120.180 91.500 -120.040 91.900 ;
        RECT -118.310 91.590 -116.950 91.900 ;
        RECT -115.220 91.500 -115.080 91.900 ;
        RECT -110.260 91.500 -110.120 91.900 ;
        RECT -108.390 91.590 -107.030 91.900 ;
        RECT -105.300 91.500 -105.160 91.900 ;
        RECT -100.340 91.500 -100.200 91.900 ;
        RECT -98.470 91.590 -97.110 91.900 ;
        RECT -95.380 91.500 -95.240 91.900 ;
        RECT -90.420 91.500 -90.280 91.900 ;
        RECT -88.550 91.590 -87.190 91.900 ;
        RECT -85.460 91.500 -85.320 91.900 ;
        RECT -80.500 91.500 -80.360 91.900 ;
        RECT -78.630 91.590 -77.270 91.900 ;
        RECT -75.540 91.500 -75.400 91.900 ;
        RECT -70.580 91.500 -70.440 91.900 ;
        RECT -68.710 91.590 -67.350 91.900 ;
        RECT -65.620 91.500 -65.480 91.900 ;
        RECT -60.660 91.500 -60.520 91.900 ;
        RECT -58.790 91.590 -57.430 91.900 ;
        RECT -55.700 91.500 -55.560 91.900 ;
        RECT -50.740 91.500 -50.600 91.900 ;
        RECT -48.870 91.590 -47.510 91.900 ;
        RECT -45.780 91.500 -45.640 91.900 ;
        RECT -40.820 91.500 -40.680 91.900 ;
        RECT -38.950 91.590 -37.590 91.900 ;
        RECT -35.860 91.500 -35.720 91.900 ;
        RECT -30.900 91.500 -30.760 91.900 ;
        RECT -29.030 91.590 -27.670 91.900 ;
        RECT -25.940 91.500 -25.800 91.900 ;
        RECT -20.980 91.500 -20.840 91.900 ;
        RECT -19.110 91.590 -17.750 91.900 ;
        RECT -16.020 91.500 -15.880 91.900 ;
        RECT -11.060 91.500 -10.920 91.900 ;
        RECT -9.190 91.590 -7.830 91.900 ;
        RECT -6.100 91.500 -5.960 91.900 ;
        RECT -1.140 91.500 -1.000 91.900 ;
        RECT 0.730 91.590 2.090 91.900 ;
        RECT 3.820 91.500 3.960 91.900 ;
        RECT 8.780 91.500 8.920 91.900 ;
        RECT 10.650 91.590 12.010 91.900 ;
        RECT 13.740 91.500 13.880 91.900 ;
        RECT 18.700 91.500 18.840 91.900 ;
        RECT 20.570 91.590 21.930 91.900 ;
        RECT 23.660 91.500 23.800 91.900 ;
        RECT -293.030 7.990 -292.570 8.300 ;
        RECT -290.840 7.990 -290.700 8.390 ;
        RECT -285.880 7.990 -285.740 8.390 ;
        RECT -284.010 7.990 -282.650 8.300 ;
        RECT -280.920 7.990 -280.780 8.390 ;
        RECT -275.960 7.990 -275.820 8.390 ;
        RECT -274.090 7.990 -272.730 8.300 ;
        RECT -271.000 7.990 -270.860 8.390 ;
        RECT -266.040 7.990 -265.900 8.390 ;
        RECT -264.170 7.990 -262.810 8.300 ;
        RECT -261.080 7.990 -260.940 8.390 ;
        RECT -256.120 7.990 -255.980 8.390 ;
        RECT -254.250 7.990 -252.890 8.300 ;
        RECT -251.160 7.990 -251.020 8.390 ;
        RECT -246.200 7.990 -246.060 8.390 ;
        RECT -244.330 7.990 -242.970 8.300 ;
        RECT -241.240 7.990 -241.100 8.390 ;
        RECT -236.280 7.990 -236.140 8.390 ;
        RECT -234.410 7.990 -233.050 8.300 ;
        RECT -231.320 7.990 -231.180 8.390 ;
        RECT -226.360 7.990 -226.220 8.390 ;
        RECT -224.490 7.990 -223.130 8.300 ;
        RECT -221.400 7.990 -221.260 8.390 ;
        RECT -216.440 7.990 -216.300 8.390 ;
        RECT -214.570 7.990 -213.210 8.300 ;
        RECT -211.480 7.990 -211.340 8.390 ;
        RECT -206.520 7.990 -206.380 8.390 ;
        RECT -204.650 7.990 -203.290 8.300 ;
        RECT -201.560 7.990 -201.420 8.390 ;
        RECT -196.600 7.990 -196.460 8.390 ;
        RECT -194.730 7.990 -193.370 8.300 ;
        RECT -191.640 7.990 -191.500 8.390 ;
        RECT -186.680 7.990 -186.540 8.390 ;
        RECT -184.810 7.990 -183.450 8.300 ;
        RECT -181.720 7.990 -181.580 8.390 ;
        RECT -176.760 7.990 -176.620 8.390 ;
        RECT -174.890 7.990 -173.530 8.300 ;
        RECT -171.800 7.990 -171.660 8.390 ;
        RECT -166.840 7.990 -166.700 8.390 ;
        RECT -164.970 7.990 -163.610 8.300 ;
        RECT -161.880 7.990 -161.740 8.390 ;
        RECT -156.920 7.990 -156.780 8.390 ;
        RECT -155.050 7.990 -153.690 8.300 ;
        RECT -151.960 7.990 -151.820 8.390 ;
        RECT -147.000 7.990 -146.860 8.390 ;
        RECT -145.130 7.990 -143.770 8.300 ;
        RECT -142.040 7.990 -141.900 8.390 ;
        RECT -137.080 7.990 -136.940 8.390 ;
        RECT -135.210 7.990 -133.850 8.300 ;
        RECT -132.120 7.990 -131.980 8.390 ;
        RECT -127.160 7.990 -127.020 8.390 ;
        RECT -125.290 7.990 -123.930 8.300 ;
        RECT -122.200 7.990 -122.060 8.390 ;
        RECT -117.240 7.990 -117.100 8.390 ;
        RECT -115.370 7.990 -114.010 8.300 ;
        RECT -112.280 7.990 -112.140 8.390 ;
        RECT -107.320 7.990 -107.180 8.390 ;
        RECT -105.450 7.990 -104.090 8.300 ;
        RECT -102.360 7.990 -102.220 8.390 ;
        RECT -97.400 7.990 -97.260 8.390 ;
        RECT -95.530 7.990 -94.170 8.300 ;
        RECT -92.440 7.990 -92.300 8.390 ;
        RECT -87.480 7.990 -87.340 8.390 ;
        RECT -85.610 7.990 -84.250 8.300 ;
        RECT -82.520 7.990 -82.380 8.390 ;
        RECT -77.560 7.990 -77.420 8.390 ;
        RECT -75.690 7.990 -74.330 8.300 ;
        RECT -72.600 7.990 -72.460 8.390 ;
        RECT -67.640 7.990 -67.500 8.390 ;
        RECT -65.770 7.990 -64.410 8.300 ;
        RECT -62.680 7.990 -62.540 8.390 ;
        RECT -57.720 7.990 -57.580 8.390 ;
        RECT -55.850 7.990 -54.490 8.300 ;
        RECT -52.760 7.990 -52.620 8.390 ;
        RECT -47.800 7.990 -47.660 8.390 ;
        RECT -45.930 7.990 -44.570 8.300 ;
        RECT -42.840 7.990 -42.700 8.390 ;
        RECT -37.880 7.990 -37.740 8.390 ;
        RECT -36.010 7.990 -34.650 8.300 ;
        RECT -32.920 7.990 -32.780 8.390 ;
        RECT -27.960 7.990 -27.820 8.390 ;
        RECT -26.090 7.990 -24.730 8.300 ;
        RECT -23.000 7.990 -22.860 8.390 ;
        RECT -18.040 7.990 -17.900 8.390 ;
        RECT -16.170 7.990 -14.810 8.300 ;
        RECT -13.080 7.990 -12.940 8.390 ;
        RECT -8.120 7.990 -7.980 8.390 ;
        RECT -6.250 7.990 -4.890 8.300 ;
        RECT -3.160 7.990 -3.020 8.390 ;
        RECT 1.800 7.990 1.940 8.390 ;
        RECT 3.670 7.990 5.030 8.300 ;
        RECT 6.760 7.990 6.900 8.390 ;
        RECT 11.720 7.990 11.860 8.390 ;
        RECT 13.590 7.990 14.950 8.300 ;
        RECT 16.680 7.990 16.820 8.390 ;
        RECT 21.640 7.990 21.780 8.390 ;
        RECT 35.230 8.320 35.950 91.910 ;
        RECT 30.930 8.310 35.950 8.320 ;
        RECT 23.510 8.260 35.950 8.310 ;
        RECT 23.510 7.990 36.110 8.260 ;
        RECT -293.030 7.860 36.110 7.990 ;
        RECT -293.030 7.850 32.250 7.860 ;
        RECT -290.840 7.450 -290.700 7.850 ;
        RECT -288.970 7.540 -287.610 7.850 ;
        RECT -285.880 7.450 -285.740 7.850 ;
        RECT -280.920 7.450 -280.780 7.850 ;
        RECT -279.050 7.540 -277.690 7.850 ;
        RECT -275.960 7.450 -275.820 7.850 ;
        RECT -271.000 7.450 -270.860 7.850 ;
        RECT -269.130 7.540 -267.770 7.850 ;
        RECT -266.040 7.450 -265.900 7.850 ;
        RECT -261.080 7.450 -260.940 7.850 ;
        RECT -259.210 7.540 -257.850 7.850 ;
        RECT -256.120 7.450 -255.980 7.850 ;
        RECT -251.160 7.450 -251.020 7.850 ;
        RECT -249.290 7.540 -247.930 7.850 ;
        RECT -246.200 7.450 -246.060 7.850 ;
        RECT -241.240 7.450 -241.100 7.850 ;
        RECT -239.370 7.540 -238.010 7.850 ;
        RECT -236.280 7.450 -236.140 7.850 ;
        RECT -231.320 7.450 -231.180 7.850 ;
        RECT -229.450 7.540 -228.090 7.850 ;
        RECT -226.360 7.450 -226.220 7.850 ;
        RECT -221.400 7.450 -221.260 7.850 ;
        RECT -219.530 7.540 -218.170 7.850 ;
        RECT -216.440 7.450 -216.300 7.850 ;
        RECT -211.480 7.450 -211.340 7.850 ;
        RECT -209.610 7.540 -208.250 7.850 ;
        RECT -206.520 7.450 -206.380 7.850 ;
        RECT -201.560 7.450 -201.420 7.850 ;
        RECT -199.690 7.540 -198.330 7.850 ;
        RECT -196.600 7.450 -196.460 7.850 ;
        RECT -191.640 7.450 -191.500 7.850 ;
        RECT -189.770 7.540 -188.410 7.850 ;
        RECT -186.680 7.450 -186.540 7.850 ;
        RECT -181.720 7.450 -181.580 7.850 ;
        RECT -179.850 7.540 -178.490 7.850 ;
        RECT -176.760 7.450 -176.620 7.850 ;
        RECT -171.800 7.450 -171.660 7.850 ;
        RECT -169.930 7.540 -168.570 7.850 ;
        RECT -166.840 7.450 -166.700 7.850 ;
        RECT -161.880 7.450 -161.740 7.850 ;
        RECT -160.010 7.540 -158.650 7.850 ;
        RECT -156.920 7.450 -156.780 7.850 ;
        RECT -151.960 7.450 -151.820 7.850 ;
        RECT -150.090 7.540 -148.730 7.850 ;
        RECT -147.000 7.450 -146.860 7.850 ;
        RECT -142.040 7.450 -141.900 7.850 ;
        RECT -140.170 7.540 -138.810 7.850 ;
        RECT -137.080 7.450 -136.940 7.850 ;
        RECT -132.120 7.450 -131.980 7.850 ;
        RECT -130.250 7.540 -128.890 7.850 ;
        RECT -127.160 7.450 -127.020 7.850 ;
        RECT -122.200 7.450 -122.060 7.850 ;
        RECT -120.330 7.540 -118.970 7.850 ;
        RECT -117.240 7.450 -117.100 7.850 ;
        RECT -112.280 7.450 -112.140 7.850 ;
        RECT -110.410 7.540 -109.050 7.850 ;
        RECT -107.320 7.450 -107.180 7.850 ;
        RECT -102.360 7.450 -102.220 7.850 ;
        RECT -100.490 7.540 -99.130 7.850 ;
        RECT -97.400 7.450 -97.260 7.850 ;
        RECT -92.440 7.450 -92.300 7.850 ;
        RECT -90.570 7.540 -89.210 7.850 ;
        RECT -87.480 7.450 -87.340 7.850 ;
        RECT -82.520 7.450 -82.380 7.850 ;
        RECT -80.650 7.540 -79.290 7.850 ;
        RECT -77.560 7.450 -77.420 7.850 ;
        RECT -72.600 7.450 -72.460 7.850 ;
        RECT -70.730 7.540 -69.370 7.850 ;
        RECT -67.640 7.450 -67.500 7.850 ;
        RECT -62.680 7.450 -62.540 7.850 ;
        RECT -60.810 7.540 -59.450 7.850 ;
        RECT -57.720 7.450 -57.580 7.850 ;
        RECT -52.760 7.450 -52.620 7.850 ;
        RECT -50.890 7.540 -49.530 7.850 ;
        RECT -47.800 7.450 -47.660 7.850 ;
        RECT -42.840 7.450 -42.700 7.850 ;
        RECT -40.970 7.540 -39.610 7.850 ;
        RECT -37.880 7.450 -37.740 7.850 ;
        RECT -32.920 7.450 -32.780 7.850 ;
        RECT -31.050 7.540 -29.690 7.850 ;
        RECT -27.960 7.450 -27.820 7.850 ;
        RECT -23.000 7.450 -22.860 7.850 ;
        RECT -21.130 7.540 -19.770 7.850 ;
        RECT -18.040 7.450 -17.900 7.850 ;
        RECT -13.080 7.450 -12.940 7.850 ;
        RECT -11.210 7.540 -9.850 7.850 ;
        RECT -8.120 7.450 -7.980 7.850 ;
        RECT -3.160 7.450 -3.020 7.850 ;
        RECT -1.290 7.540 0.070 7.850 ;
        RECT 1.800 7.450 1.940 7.850 ;
        RECT 6.760 7.450 6.900 7.850 ;
        RECT 8.630 7.540 9.990 7.850 ;
        RECT 11.720 7.450 11.860 7.850 ;
        RECT 16.680 7.450 16.820 7.850 ;
        RECT 18.550 7.540 19.910 7.850 ;
        RECT 21.640 7.450 21.780 7.850 ;
        RECT 35.220 5.070 36.110 7.860 ;
        RECT 35.220 4.870 36.200 5.070 ;
        RECT 35.210 4.380 36.200 4.870 ;
        RECT 35.220 4.100 36.200 4.380 ;
        RECT 35.480 -80.080 36.200 4.100 ;
        RECT -292.670 -80.960 -292.210 -80.650 ;
        RECT -290.480 -80.960 -290.340 -80.560 ;
        RECT -285.520 -80.960 -285.380 -80.560 ;
        RECT -283.650 -80.960 -282.290 -80.650 ;
        RECT -280.560 -80.960 -280.420 -80.560 ;
        RECT -275.600 -80.960 -275.460 -80.560 ;
        RECT -273.730 -80.960 -272.370 -80.650 ;
        RECT -270.640 -80.960 -270.500 -80.560 ;
        RECT -265.680 -80.960 -265.540 -80.560 ;
        RECT -263.810 -80.960 -262.450 -80.650 ;
        RECT -260.720 -80.960 -260.580 -80.560 ;
        RECT -255.760 -80.960 -255.620 -80.560 ;
        RECT -253.890 -80.960 -252.530 -80.650 ;
        RECT -250.800 -80.960 -250.660 -80.560 ;
        RECT -245.840 -80.960 -245.700 -80.560 ;
        RECT -243.970 -80.960 -242.610 -80.650 ;
        RECT -240.880 -80.960 -240.740 -80.560 ;
        RECT -235.920 -80.960 -235.780 -80.560 ;
        RECT -234.050 -80.960 -232.690 -80.650 ;
        RECT -230.960 -80.960 -230.820 -80.560 ;
        RECT -226.000 -80.960 -225.860 -80.560 ;
        RECT -224.130 -80.960 -222.770 -80.650 ;
        RECT -221.040 -80.960 -220.900 -80.560 ;
        RECT -216.080 -80.960 -215.940 -80.560 ;
        RECT -214.210 -80.960 -212.850 -80.650 ;
        RECT -211.120 -80.960 -210.980 -80.560 ;
        RECT -206.160 -80.960 -206.020 -80.560 ;
        RECT -204.290 -80.960 -202.930 -80.650 ;
        RECT -201.200 -80.960 -201.060 -80.560 ;
        RECT -196.240 -80.960 -196.100 -80.560 ;
        RECT -194.370 -80.960 -193.010 -80.650 ;
        RECT -191.280 -80.960 -191.140 -80.560 ;
        RECT -186.320 -80.960 -186.180 -80.560 ;
        RECT -184.450 -80.960 -183.090 -80.650 ;
        RECT -181.360 -80.960 -181.220 -80.560 ;
        RECT -176.400 -80.960 -176.260 -80.560 ;
        RECT -174.530 -80.960 -173.170 -80.650 ;
        RECT -171.440 -80.960 -171.300 -80.560 ;
        RECT -166.480 -80.960 -166.340 -80.560 ;
        RECT -164.610 -80.960 -163.250 -80.650 ;
        RECT -161.520 -80.960 -161.380 -80.560 ;
        RECT -156.560 -80.960 -156.420 -80.560 ;
        RECT -154.690 -80.960 -153.330 -80.650 ;
        RECT -151.600 -80.960 -151.460 -80.560 ;
        RECT -146.640 -80.960 -146.500 -80.560 ;
        RECT -144.770 -80.960 -143.410 -80.650 ;
        RECT -141.680 -80.960 -141.540 -80.560 ;
        RECT -136.720 -80.960 -136.580 -80.560 ;
        RECT -134.850 -80.960 -133.490 -80.650 ;
        RECT -131.760 -80.960 -131.620 -80.560 ;
        RECT -126.800 -80.960 -126.660 -80.560 ;
        RECT -124.930 -80.960 -123.570 -80.650 ;
        RECT -121.840 -80.960 -121.700 -80.560 ;
        RECT -116.880 -80.960 -116.740 -80.560 ;
        RECT -115.010 -80.960 -113.650 -80.650 ;
        RECT -111.920 -80.960 -111.780 -80.560 ;
        RECT -106.960 -80.960 -106.820 -80.560 ;
        RECT -105.090 -80.960 -103.730 -80.650 ;
        RECT -102.000 -80.960 -101.860 -80.560 ;
        RECT -97.040 -80.960 -96.900 -80.560 ;
        RECT -95.170 -80.960 -93.810 -80.650 ;
        RECT -92.080 -80.960 -91.940 -80.560 ;
        RECT -87.120 -80.960 -86.980 -80.560 ;
        RECT -85.250 -80.960 -83.890 -80.650 ;
        RECT -82.160 -80.960 -82.020 -80.560 ;
        RECT -77.200 -80.960 -77.060 -80.560 ;
        RECT -75.330 -80.960 -73.970 -80.650 ;
        RECT -72.240 -80.960 -72.100 -80.560 ;
        RECT -67.280 -80.960 -67.140 -80.560 ;
        RECT -65.410 -80.960 -64.050 -80.650 ;
        RECT -62.320 -80.960 -62.180 -80.560 ;
        RECT -57.360 -80.960 -57.220 -80.560 ;
        RECT -55.490 -80.960 -54.130 -80.650 ;
        RECT -52.400 -80.960 -52.260 -80.560 ;
        RECT -47.440 -80.960 -47.300 -80.560 ;
        RECT -45.570 -80.960 -44.210 -80.650 ;
        RECT -42.480 -80.960 -42.340 -80.560 ;
        RECT -37.520 -80.960 -37.380 -80.560 ;
        RECT -35.650 -80.960 -34.290 -80.650 ;
        RECT -32.560 -80.960 -32.420 -80.560 ;
        RECT -27.600 -80.960 -27.460 -80.560 ;
        RECT -25.730 -80.960 -24.370 -80.650 ;
        RECT -22.640 -80.960 -22.500 -80.560 ;
        RECT -17.680 -80.960 -17.540 -80.560 ;
        RECT -15.810 -80.960 -14.450 -80.650 ;
        RECT -12.720 -80.960 -12.580 -80.560 ;
        RECT -7.760 -80.960 -7.620 -80.560 ;
        RECT -5.890 -80.960 -4.530 -80.650 ;
        RECT -2.800 -80.960 -2.660 -80.560 ;
        RECT 2.160 -80.960 2.300 -80.560 ;
        RECT 4.030 -80.960 5.390 -80.650 ;
        RECT 7.120 -80.960 7.260 -80.560 ;
        RECT 12.080 -80.960 12.220 -80.560 ;
        RECT 13.950 -80.960 15.310 -80.650 ;
        RECT 17.040 -80.960 17.180 -80.560 ;
        RECT 22.000 -80.960 22.140 -80.560 ;
        RECT 35.600 -80.630 36.060 -80.080 ;
        RECT 31.290 -80.640 36.060 -80.630 ;
        RECT 23.870 -80.960 36.060 -80.640 ;
        RECT -292.670 -81.090 36.060 -80.960 ;
        RECT -292.670 -81.100 32.610 -81.090 ;
        RECT -290.480 -81.500 -290.340 -81.100 ;
        RECT -288.610 -81.410 -287.250 -81.100 ;
        RECT -285.520 -81.500 -285.380 -81.100 ;
        RECT -280.560 -81.500 -280.420 -81.100 ;
        RECT -278.690 -81.410 -277.330 -81.100 ;
        RECT -275.600 -81.500 -275.460 -81.100 ;
        RECT -270.640 -81.500 -270.500 -81.100 ;
        RECT -268.770 -81.410 -267.410 -81.100 ;
        RECT -265.680 -81.500 -265.540 -81.100 ;
        RECT -260.720 -81.500 -260.580 -81.100 ;
        RECT -258.850 -81.410 -257.490 -81.100 ;
        RECT -255.760 -81.500 -255.620 -81.100 ;
        RECT -250.800 -81.500 -250.660 -81.100 ;
        RECT -248.930 -81.410 -247.570 -81.100 ;
        RECT -245.840 -81.500 -245.700 -81.100 ;
        RECT -240.880 -81.500 -240.740 -81.100 ;
        RECT -239.010 -81.410 -237.650 -81.100 ;
        RECT -235.920 -81.500 -235.780 -81.100 ;
        RECT -230.960 -81.500 -230.820 -81.100 ;
        RECT -229.090 -81.410 -227.730 -81.100 ;
        RECT -226.000 -81.500 -225.860 -81.100 ;
        RECT -221.040 -81.500 -220.900 -81.100 ;
        RECT -219.170 -81.410 -217.810 -81.100 ;
        RECT -216.080 -81.500 -215.940 -81.100 ;
        RECT -211.120 -81.500 -210.980 -81.100 ;
        RECT -209.250 -81.410 -207.890 -81.100 ;
        RECT -206.160 -81.500 -206.020 -81.100 ;
        RECT -201.200 -81.500 -201.060 -81.100 ;
        RECT -199.330 -81.410 -197.970 -81.100 ;
        RECT -196.240 -81.500 -196.100 -81.100 ;
        RECT -191.280 -81.500 -191.140 -81.100 ;
        RECT -189.410 -81.410 -188.050 -81.100 ;
        RECT -186.320 -81.500 -186.180 -81.100 ;
        RECT -181.360 -81.500 -181.220 -81.100 ;
        RECT -179.490 -81.410 -178.130 -81.100 ;
        RECT -176.400 -81.500 -176.260 -81.100 ;
        RECT -171.440 -81.500 -171.300 -81.100 ;
        RECT -169.570 -81.410 -168.210 -81.100 ;
        RECT -166.480 -81.500 -166.340 -81.100 ;
        RECT -161.520 -81.500 -161.380 -81.100 ;
        RECT -159.650 -81.410 -158.290 -81.100 ;
        RECT -156.560 -81.500 -156.420 -81.100 ;
        RECT -151.600 -81.500 -151.460 -81.100 ;
        RECT -149.730 -81.410 -148.370 -81.100 ;
        RECT -146.640 -81.500 -146.500 -81.100 ;
        RECT -141.680 -81.500 -141.540 -81.100 ;
        RECT -139.810 -81.410 -138.450 -81.100 ;
        RECT -136.720 -81.500 -136.580 -81.100 ;
        RECT -131.760 -81.500 -131.620 -81.100 ;
        RECT -129.890 -81.410 -128.530 -81.100 ;
        RECT -126.800 -81.500 -126.660 -81.100 ;
        RECT -121.840 -81.500 -121.700 -81.100 ;
        RECT -119.970 -81.410 -118.610 -81.100 ;
        RECT -116.880 -81.500 -116.740 -81.100 ;
        RECT -111.920 -81.500 -111.780 -81.100 ;
        RECT -110.050 -81.410 -108.690 -81.100 ;
        RECT -106.960 -81.500 -106.820 -81.100 ;
        RECT -102.000 -81.500 -101.860 -81.100 ;
        RECT -100.130 -81.410 -98.770 -81.100 ;
        RECT -97.040 -81.500 -96.900 -81.100 ;
        RECT -92.080 -81.500 -91.940 -81.100 ;
        RECT -90.210 -81.410 -88.850 -81.100 ;
        RECT -87.120 -81.500 -86.980 -81.100 ;
        RECT -82.160 -81.500 -82.020 -81.100 ;
        RECT -80.290 -81.410 -78.930 -81.100 ;
        RECT -77.200 -81.500 -77.060 -81.100 ;
        RECT -72.240 -81.500 -72.100 -81.100 ;
        RECT -70.370 -81.410 -69.010 -81.100 ;
        RECT -67.280 -81.500 -67.140 -81.100 ;
        RECT -62.320 -81.500 -62.180 -81.100 ;
        RECT -60.450 -81.410 -59.090 -81.100 ;
        RECT -57.360 -81.500 -57.220 -81.100 ;
        RECT -52.400 -81.500 -52.260 -81.100 ;
        RECT -50.530 -81.410 -49.170 -81.100 ;
        RECT -47.440 -81.500 -47.300 -81.100 ;
        RECT -42.480 -81.500 -42.340 -81.100 ;
        RECT -40.610 -81.410 -39.250 -81.100 ;
        RECT -37.520 -81.500 -37.380 -81.100 ;
        RECT -32.560 -81.500 -32.420 -81.100 ;
        RECT -30.690 -81.410 -29.330 -81.100 ;
        RECT -27.600 -81.500 -27.460 -81.100 ;
        RECT -22.640 -81.500 -22.500 -81.100 ;
        RECT -20.770 -81.410 -19.410 -81.100 ;
        RECT -17.680 -81.500 -17.540 -81.100 ;
        RECT -12.720 -81.500 -12.580 -81.100 ;
        RECT -10.850 -81.410 -9.490 -81.100 ;
        RECT -7.760 -81.500 -7.620 -81.100 ;
        RECT -2.800 -81.500 -2.660 -81.100 ;
        RECT -0.930 -81.410 0.430 -81.100 ;
        RECT 2.160 -81.500 2.300 -81.100 ;
        RECT 7.120 -81.500 7.260 -81.100 ;
        RECT 8.990 -81.410 10.350 -81.100 ;
        RECT 12.080 -81.500 12.220 -81.100 ;
        RECT 17.040 -81.500 17.180 -81.100 ;
        RECT 18.910 -81.410 20.270 -81.100 ;
        RECT 22.000 -81.500 22.140 -81.100 ;
        RECT -294.430 -175.540 -293.970 -175.230 ;
        RECT -292.240 -175.540 -292.100 -175.140 ;
        RECT -287.280 -175.540 -287.140 -175.140 ;
        RECT -285.410 -175.540 -284.050 -175.230 ;
        RECT -282.320 -175.540 -282.180 -175.140 ;
        RECT -277.360 -175.540 -277.220 -175.140 ;
        RECT -275.490 -175.540 -274.130 -175.230 ;
        RECT -272.400 -175.540 -272.260 -175.140 ;
        RECT -267.440 -175.540 -267.300 -175.140 ;
        RECT -265.570 -175.540 -264.210 -175.230 ;
        RECT -262.480 -175.540 -262.340 -175.140 ;
        RECT -257.520 -175.540 -257.380 -175.140 ;
        RECT -255.650 -175.540 -254.290 -175.230 ;
        RECT -252.560 -175.540 -252.420 -175.140 ;
        RECT -247.600 -175.540 -247.460 -175.140 ;
        RECT -245.730 -175.540 -244.370 -175.230 ;
        RECT -242.640 -175.540 -242.500 -175.140 ;
        RECT -237.680 -175.540 -237.540 -175.140 ;
        RECT -235.810 -175.540 -234.450 -175.230 ;
        RECT -232.720 -175.540 -232.580 -175.140 ;
        RECT -227.760 -175.540 -227.620 -175.140 ;
        RECT -225.890 -175.540 -224.530 -175.230 ;
        RECT -222.800 -175.540 -222.660 -175.140 ;
        RECT -217.840 -175.540 -217.700 -175.140 ;
        RECT -215.970 -175.540 -214.610 -175.230 ;
        RECT -212.880 -175.540 -212.740 -175.140 ;
        RECT -207.920 -175.540 -207.780 -175.140 ;
        RECT -206.050 -175.540 -204.690 -175.230 ;
        RECT -202.960 -175.540 -202.820 -175.140 ;
        RECT -198.000 -175.540 -197.860 -175.140 ;
        RECT -196.130 -175.540 -194.770 -175.230 ;
        RECT -193.040 -175.540 -192.900 -175.140 ;
        RECT -188.080 -175.540 -187.940 -175.140 ;
        RECT -186.210 -175.540 -184.850 -175.230 ;
        RECT -183.120 -175.540 -182.980 -175.140 ;
        RECT -178.160 -175.540 -178.020 -175.140 ;
        RECT -176.290 -175.540 -174.930 -175.230 ;
        RECT -173.200 -175.540 -173.060 -175.140 ;
        RECT -168.240 -175.540 -168.100 -175.140 ;
        RECT -166.370 -175.540 -165.010 -175.230 ;
        RECT -163.280 -175.540 -163.140 -175.140 ;
        RECT -158.320 -175.540 -158.180 -175.140 ;
        RECT -156.450 -175.540 -155.090 -175.230 ;
        RECT -153.360 -175.540 -153.220 -175.140 ;
        RECT -148.400 -175.540 -148.260 -175.140 ;
        RECT -146.530 -175.540 -145.170 -175.230 ;
        RECT -143.440 -175.540 -143.300 -175.140 ;
        RECT -138.480 -175.540 -138.340 -175.140 ;
        RECT -136.610 -175.540 -135.250 -175.230 ;
        RECT -133.520 -175.540 -133.380 -175.140 ;
        RECT -128.560 -175.540 -128.420 -175.140 ;
        RECT -126.690 -175.540 -125.330 -175.230 ;
        RECT -123.600 -175.540 -123.460 -175.140 ;
        RECT -118.640 -175.540 -118.500 -175.140 ;
        RECT -116.770 -175.540 -115.410 -175.230 ;
        RECT -113.680 -175.540 -113.540 -175.140 ;
        RECT -108.720 -175.540 -108.580 -175.140 ;
        RECT -106.850 -175.540 -105.490 -175.230 ;
        RECT -103.760 -175.540 -103.620 -175.140 ;
        RECT -98.800 -175.540 -98.660 -175.140 ;
        RECT -96.930 -175.540 -95.570 -175.230 ;
        RECT -93.840 -175.540 -93.700 -175.140 ;
        RECT -88.880 -175.540 -88.740 -175.140 ;
        RECT -87.010 -175.540 -85.650 -175.230 ;
        RECT -83.920 -175.540 -83.780 -175.140 ;
        RECT -78.960 -175.540 -78.820 -175.140 ;
        RECT -77.090 -175.540 -75.730 -175.230 ;
        RECT -74.000 -175.540 -73.860 -175.140 ;
        RECT -69.040 -175.540 -68.900 -175.140 ;
        RECT -67.170 -175.540 -65.810 -175.230 ;
        RECT -64.080 -175.540 -63.940 -175.140 ;
        RECT -59.120 -175.540 -58.980 -175.140 ;
        RECT -57.250 -175.540 -55.890 -175.230 ;
        RECT -54.160 -175.540 -54.020 -175.140 ;
        RECT -49.200 -175.540 -49.060 -175.140 ;
        RECT -47.330 -175.540 -45.970 -175.230 ;
        RECT -44.240 -175.540 -44.100 -175.140 ;
        RECT -39.280 -175.540 -39.140 -175.140 ;
        RECT -37.410 -175.540 -36.050 -175.230 ;
        RECT -34.320 -175.540 -34.180 -175.140 ;
        RECT -29.360 -175.540 -29.220 -175.140 ;
        RECT -27.490 -175.540 -26.130 -175.230 ;
        RECT -24.400 -175.540 -24.260 -175.140 ;
        RECT -19.440 -175.540 -19.300 -175.140 ;
        RECT -17.570 -175.540 -16.210 -175.230 ;
        RECT -14.480 -175.540 -14.340 -175.140 ;
        RECT -9.520 -175.540 -9.380 -175.140 ;
        RECT -7.650 -175.540 -6.290 -175.230 ;
        RECT -4.560 -175.540 -4.420 -175.140 ;
        RECT 0.400 -175.540 0.540 -175.140 ;
        RECT 2.270 -175.540 3.630 -175.230 ;
        RECT 5.360 -175.540 5.500 -175.140 ;
        RECT 10.320 -175.540 10.460 -175.140 ;
        RECT 12.190 -175.540 13.550 -175.230 ;
        RECT 15.280 -175.540 15.420 -175.140 ;
        RECT 20.240 -175.540 20.380 -175.140 ;
        RECT 33.770 -175.210 34.510 -81.090 ;
        RECT 29.530 -175.220 34.510 -175.210 ;
        RECT 22.110 -175.540 34.510 -175.220 ;
        RECT -294.430 -175.670 34.510 -175.540 ;
        RECT -294.430 -175.680 30.850 -175.670 ;
        RECT -292.240 -176.080 -292.100 -175.680 ;
        RECT -290.370 -175.990 -289.010 -175.680 ;
        RECT -287.280 -176.080 -287.140 -175.680 ;
        RECT -282.320 -176.080 -282.180 -175.680 ;
        RECT -280.450 -175.990 -279.090 -175.680 ;
        RECT -277.360 -176.080 -277.220 -175.680 ;
        RECT -272.400 -176.080 -272.260 -175.680 ;
        RECT -270.530 -175.990 -269.170 -175.680 ;
        RECT -267.440 -176.080 -267.300 -175.680 ;
        RECT -262.480 -176.080 -262.340 -175.680 ;
        RECT -260.610 -175.990 -259.250 -175.680 ;
        RECT -257.520 -176.080 -257.380 -175.680 ;
        RECT -252.560 -176.080 -252.420 -175.680 ;
        RECT -250.690 -175.990 -249.330 -175.680 ;
        RECT -247.600 -176.080 -247.460 -175.680 ;
        RECT -242.640 -176.080 -242.500 -175.680 ;
        RECT -240.770 -175.990 -239.410 -175.680 ;
        RECT -237.680 -176.080 -237.540 -175.680 ;
        RECT -232.720 -176.080 -232.580 -175.680 ;
        RECT -230.850 -175.990 -229.490 -175.680 ;
        RECT -227.760 -176.080 -227.620 -175.680 ;
        RECT -222.800 -176.080 -222.660 -175.680 ;
        RECT -220.930 -175.990 -219.570 -175.680 ;
        RECT -217.840 -176.080 -217.700 -175.680 ;
        RECT -212.880 -176.080 -212.740 -175.680 ;
        RECT -211.010 -175.990 -209.650 -175.680 ;
        RECT -207.920 -176.080 -207.780 -175.680 ;
        RECT -202.960 -176.080 -202.820 -175.680 ;
        RECT -201.090 -175.990 -199.730 -175.680 ;
        RECT -198.000 -176.080 -197.860 -175.680 ;
        RECT -193.040 -176.080 -192.900 -175.680 ;
        RECT -191.170 -175.990 -189.810 -175.680 ;
        RECT -188.080 -176.080 -187.940 -175.680 ;
        RECT -183.120 -176.080 -182.980 -175.680 ;
        RECT -181.250 -175.990 -179.890 -175.680 ;
        RECT -178.160 -176.080 -178.020 -175.680 ;
        RECT -173.200 -176.080 -173.060 -175.680 ;
        RECT -171.330 -175.990 -169.970 -175.680 ;
        RECT -168.240 -176.080 -168.100 -175.680 ;
        RECT -163.280 -176.080 -163.140 -175.680 ;
        RECT -161.410 -175.990 -160.050 -175.680 ;
        RECT -158.320 -176.080 -158.180 -175.680 ;
        RECT -153.360 -176.080 -153.220 -175.680 ;
        RECT -151.490 -175.990 -150.130 -175.680 ;
        RECT -148.400 -176.080 -148.260 -175.680 ;
        RECT -143.440 -176.080 -143.300 -175.680 ;
        RECT -141.570 -175.990 -140.210 -175.680 ;
        RECT -138.480 -176.080 -138.340 -175.680 ;
        RECT -133.520 -176.080 -133.380 -175.680 ;
        RECT -131.650 -175.990 -130.290 -175.680 ;
        RECT -128.560 -176.080 -128.420 -175.680 ;
        RECT -123.600 -176.080 -123.460 -175.680 ;
        RECT -121.730 -175.990 -120.370 -175.680 ;
        RECT -118.640 -176.080 -118.500 -175.680 ;
        RECT -113.680 -176.080 -113.540 -175.680 ;
        RECT -111.810 -175.990 -110.450 -175.680 ;
        RECT -108.720 -176.080 -108.580 -175.680 ;
        RECT -103.760 -176.080 -103.620 -175.680 ;
        RECT -101.890 -175.990 -100.530 -175.680 ;
        RECT -98.800 -176.080 -98.660 -175.680 ;
        RECT -93.840 -176.080 -93.700 -175.680 ;
        RECT -91.970 -175.990 -90.610 -175.680 ;
        RECT -88.880 -176.080 -88.740 -175.680 ;
        RECT -83.920 -176.080 -83.780 -175.680 ;
        RECT -82.050 -175.990 -80.690 -175.680 ;
        RECT -78.960 -176.080 -78.820 -175.680 ;
        RECT -74.000 -176.080 -73.860 -175.680 ;
        RECT -72.130 -175.990 -70.770 -175.680 ;
        RECT -69.040 -176.080 -68.900 -175.680 ;
        RECT -64.080 -176.080 -63.940 -175.680 ;
        RECT -62.210 -175.990 -60.850 -175.680 ;
        RECT -59.120 -176.080 -58.980 -175.680 ;
        RECT -54.160 -176.080 -54.020 -175.680 ;
        RECT -52.290 -175.990 -50.930 -175.680 ;
        RECT -49.200 -176.080 -49.060 -175.680 ;
        RECT -44.240 -176.080 -44.100 -175.680 ;
        RECT -42.370 -175.990 -41.010 -175.680 ;
        RECT -39.280 -176.080 -39.140 -175.680 ;
        RECT -34.320 -176.080 -34.180 -175.680 ;
        RECT -32.450 -175.990 -31.090 -175.680 ;
        RECT -29.360 -176.080 -29.220 -175.680 ;
        RECT -24.400 -176.080 -24.260 -175.680 ;
        RECT -22.530 -175.990 -21.170 -175.680 ;
        RECT -19.440 -176.080 -19.300 -175.680 ;
        RECT -14.480 -176.080 -14.340 -175.680 ;
        RECT -12.610 -175.990 -11.250 -175.680 ;
        RECT -9.520 -176.080 -9.380 -175.680 ;
        RECT -4.560 -176.080 -4.420 -175.680 ;
        RECT -2.690 -175.990 -1.330 -175.680 ;
        RECT 0.400 -176.080 0.540 -175.680 ;
        RECT 5.360 -176.080 5.500 -175.680 ;
        RECT 7.230 -175.990 8.590 -175.680 ;
        RECT 10.320 -176.080 10.460 -175.680 ;
        RECT 15.280 -176.080 15.420 -175.680 ;
        RECT 17.150 -175.990 18.510 -175.680 ;
        RECT 20.240 -176.080 20.380 -175.680 ;
    END
  END i_srclk
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -288.220 95.135 -284.260 95.140 ;
        RECT -278.300 95.135 -274.340 95.140 ;
        RECT -268.380 95.135 -264.420 95.140 ;
        RECT -258.460 95.135 -254.500 95.140 ;
        RECT -248.540 95.135 -244.580 95.140 ;
        RECT -238.620 95.135 -234.660 95.140 ;
        RECT -228.700 95.135 -224.740 95.140 ;
        RECT -218.780 95.135 -214.820 95.140 ;
        RECT -208.860 95.135 -204.900 95.140 ;
        RECT -198.940 95.135 -194.980 95.140 ;
        RECT -189.020 95.135 -185.060 95.140 ;
        RECT -179.100 95.135 -175.140 95.140 ;
        RECT -169.180 95.135 -165.220 95.140 ;
        RECT -159.260 95.135 -155.300 95.140 ;
        RECT -149.340 95.135 -145.380 95.140 ;
        RECT -139.420 95.135 -135.460 95.140 ;
        RECT -129.500 95.135 -125.540 95.140 ;
        RECT -119.580 95.135 -115.620 95.140 ;
        RECT -109.660 95.135 -105.700 95.140 ;
        RECT -99.740 95.135 -95.780 95.140 ;
        RECT -89.820 95.135 -85.860 95.140 ;
        RECT -79.900 95.135 -75.940 95.140 ;
        RECT -69.980 95.135 -66.020 95.140 ;
        RECT -60.060 95.135 -56.100 95.140 ;
        RECT -50.140 95.135 -46.180 95.140 ;
        RECT -40.220 95.135 -36.260 95.140 ;
        RECT -30.300 95.135 -26.340 95.140 ;
        RECT -20.380 95.135 -16.420 95.140 ;
        RECT -10.460 95.135 -6.500 95.140 ;
        RECT -0.540 95.135 3.420 95.140 ;
        RECT 9.380 95.135 13.340 95.140 ;
        RECT 19.300 95.135 23.260 95.140 ;
        RECT -288.925 93.765 -283.615 95.135 ;
        RECT -279.005 93.765 -273.695 95.135 ;
        RECT -269.085 93.765 -263.775 95.135 ;
        RECT -259.165 93.765 -253.855 95.135 ;
        RECT -249.245 93.765 -243.935 95.135 ;
        RECT -239.325 93.765 -234.015 95.135 ;
        RECT -229.405 93.765 -224.095 95.135 ;
        RECT -219.485 93.765 -214.175 95.135 ;
        RECT -209.565 93.765 -204.255 95.135 ;
        RECT -199.645 93.765 -194.335 95.135 ;
        RECT -189.725 93.765 -184.415 95.135 ;
        RECT -179.805 93.765 -174.495 95.135 ;
        RECT -169.885 93.765 -164.575 95.135 ;
        RECT -159.965 93.765 -154.655 95.135 ;
        RECT -150.045 93.765 -144.735 95.135 ;
        RECT -140.125 93.765 -134.815 95.135 ;
        RECT -130.205 93.765 -124.895 95.135 ;
        RECT -120.285 93.765 -114.975 95.135 ;
        RECT -110.365 93.765 -105.055 95.135 ;
        RECT -100.445 93.765 -95.135 95.135 ;
        RECT -90.525 93.765 -85.215 95.135 ;
        RECT -80.605 93.765 -75.295 95.135 ;
        RECT -70.685 93.765 -65.375 95.135 ;
        RECT -60.765 93.765 -55.455 95.135 ;
        RECT -50.845 93.765 -45.535 95.135 ;
        RECT -40.925 93.765 -35.615 95.135 ;
        RECT -31.005 93.765 -25.695 95.135 ;
        RECT -21.085 93.765 -15.775 95.135 ;
        RECT -11.165 93.765 -5.855 95.135 ;
        RECT -1.245 93.765 4.065 95.135 ;
        RECT 8.675 93.765 13.985 95.135 ;
        RECT 18.595 93.765 23.905 95.135 ;
        RECT -288.220 93.760 -284.260 93.765 ;
        RECT -278.300 93.760 -274.340 93.765 ;
        RECT -268.380 93.760 -264.420 93.765 ;
        RECT -258.460 93.760 -254.500 93.765 ;
        RECT -248.540 93.760 -244.580 93.765 ;
        RECT -238.620 93.760 -234.660 93.765 ;
        RECT -228.700 93.760 -224.740 93.765 ;
        RECT -218.780 93.760 -214.820 93.765 ;
        RECT -208.860 93.760 -204.900 93.765 ;
        RECT -198.940 93.760 -194.980 93.765 ;
        RECT -189.020 93.760 -185.060 93.765 ;
        RECT -179.100 93.760 -175.140 93.765 ;
        RECT -169.180 93.760 -165.220 93.765 ;
        RECT -159.260 93.760 -155.300 93.765 ;
        RECT -149.340 93.760 -145.380 93.765 ;
        RECT -139.420 93.760 -135.460 93.765 ;
        RECT -129.500 93.760 -125.540 93.765 ;
        RECT -119.580 93.760 -115.620 93.765 ;
        RECT -109.660 93.760 -105.700 93.765 ;
        RECT -99.740 93.760 -95.780 93.765 ;
        RECT -89.820 93.760 -85.860 93.765 ;
        RECT -79.900 93.760 -75.940 93.765 ;
        RECT -69.980 93.760 -66.020 93.765 ;
        RECT -60.060 93.760 -56.100 93.765 ;
        RECT -50.140 93.760 -46.180 93.765 ;
        RECT -40.220 93.760 -36.260 93.765 ;
        RECT -30.300 93.760 -26.340 93.765 ;
        RECT -20.380 93.760 -16.420 93.765 ;
        RECT -10.460 93.760 -6.500 93.765 ;
        RECT -0.540 93.760 3.420 93.765 ;
        RECT 9.380 93.760 13.340 93.765 ;
        RECT 19.300 93.760 23.260 93.765 ;
        RECT -281.850 93.225 -281.680 93.415 ;
        RECT -280.940 93.225 -280.770 93.415 ;
        RECT -271.930 93.225 -271.760 93.415 ;
        RECT -271.020 93.225 -270.850 93.415 ;
        RECT -262.010 93.225 -261.840 93.415 ;
        RECT -261.100 93.225 -260.930 93.415 ;
        RECT -252.090 93.225 -251.920 93.415 ;
        RECT -251.180 93.225 -251.010 93.415 ;
        RECT -242.170 93.225 -242.000 93.415 ;
        RECT -241.260 93.225 -241.090 93.415 ;
        RECT -232.250 93.225 -232.080 93.415 ;
        RECT -231.340 93.225 -231.170 93.415 ;
        RECT -222.330 93.225 -222.160 93.415 ;
        RECT -221.420 93.225 -221.250 93.415 ;
        RECT -212.410 93.225 -212.240 93.415 ;
        RECT -211.500 93.225 -211.330 93.415 ;
        RECT -202.490 93.225 -202.320 93.415 ;
        RECT -201.580 93.225 -201.410 93.415 ;
        RECT -192.570 93.225 -192.400 93.415 ;
        RECT -191.660 93.225 -191.490 93.415 ;
        RECT -182.650 93.225 -182.480 93.415 ;
        RECT -181.740 93.225 -181.570 93.415 ;
        RECT -172.730 93.225 -172.560 93.415 ;
        RECT -171.820 93.225 -171.650 93.415 ;
        RECT -162.810 93.225 -162.640 93.415 ;
        RECT -161.900 93.225 -161.730 93.415 ;
        RECT -152.890 93.225 -152.720 93.415 ;
        RECT -151.980 93.225 -151.810 93.415 ;
        RECT -142.970 93.225 -142.800 93.415 ;
        RECT -142.060 93.225 -141.890 93.415 ;
        RECT -133.050 93.225 -132.880 93.415 ;
        RECT -132.140 93.225 -131.970 93.415 ;
        RECT -123.130 93.225 -122.960 93.415 ;
        RECT -122.220 93.225 -122.050 93.415 ;
        RECT -113.210 93.225 -113.040 93.415 ;
        RECT -112.300 93.225 -112.130 93.415 ;
        RECT -103.290 93.225 -103.120 93.415 ;
        RECT -102.380 93.225 -102.210 93.415 ;
        RECT -93.370 93.225 -93.200 93.415 ;
        RECT -92.460 93.225 -92.290 93.415 ;
        RECT -83.450 93.225 -83.280 93.415 ;
        RECT -82.540 93.225 -82.370 93.415 ;
        RECT -73.530 93.225 -73.360 93.415 ;
        RECT -72.620 93.225 -72.450 93.415 ;
        RECT -63.610 93.225 -63.440 93.415 ;
        RECT -62.700 93.225 -62.530 93.415 ;
        RECT -53.690 93.225 -53.520 93.415 ;
        RECT -52.780 93.225 -52.610 93.415 ;
        RECT -43.770 93.225 -43.600 93.415 ;
        RECT -42.860 93.225 -42.690 93.415 ;
        RECT -33.850 93.225 -33.680 93.415 ;
        RECT -32.940 93.225 -32.770 93.415 ;
        RECT -23.930 93.225 -23.760 93.415 ;
        RECT -23.020 93.225 -22.850 93.415 ;
        RECT -14.010 93.225 -13.840 93.415 ;
        RECT -13.100 93.225 -12.930 93.415 ;
        RECT -4.090 93.225 -3.920 93.415 ;
        RECT -3.180 93.225 -3.010 93.415 ;
        RECT 5.830 93.225 6.000 93.415 ;
        RECT 6.740 93.225 6.910 93.415 ;
        RECT 15.750 93.225 15.920 93.415 ;
        RECT 16.660 93.225 16.830 93.415 ;
        RECT -282.915 93.220 -281.565 93.225 ;
        RECT -281.055 93.220 -279.705 93.225 ;
        RECT -282.915 92.320 -279.705 93.220 ;
        RECT -282.915 92.315 -281.565 92.320 ;
        RECT -281.055 92.315 -279.705 92.320 ;
        RECT -272.995 93.220 -271.645 93.225 ;
        RECT -271.135 93.220 -269.785 93.225 ;
        RECT -272.995 92.320 -269.785 93.220 ;
        RECT -272.995 92.315 -271.645 92.320 ;
        RECT -271.135 92.315 -269.785 92.320 ;
        RECT -263.075 93.220 -261.725 93.225 ;
        RECT -261.215 93.220 -259.865 93.225 ;
        RECT -263.075 92.320 -259.865 93.220 ;
        RECT -263.075 92.315 -261.725 92.320 ;
        RECT -261.215 92.315 -259.865 92.320 ;
        RECT -253.155 93.220 -251.805 93.225 ;
        RECT -251.295 93.220 -249.945 93.225 ;
        RECT -253.155 92.320 -249.945 93.220 ;
        RECT -253.155 92.315 -251.805 92.320 ;
        RECT -251.295 92.315 -249.945 92.320 ;
        RECT -243.235 93.220 -241.885 93.225 ;
        RECT -241.375 93.220 -240.025 93.225 ;
        RECT -243.235 92.320 -240.025 93.220 ;
        RECT -243.235 92.315 -241.885 92.320 ;
        RECT -241.375 92.315 -240.025 92.320 ;
        RECT -233.315 93.220 -231.965 93.225 ;
        RECT -231.455 93.220 -230.105 93.225 ;
        RECT -233.315 92.320 -230.105 93.220 ;
        RECT -233.315 92.315 -231.965 92.320 ;
        RECT -231.455 92.315 -230.105 92.320 ;
        RECT -223.395 93.220 -222.045 93.225 ;
        RECT -221.535 93.220 -220.185 93.225 ;
        RECT -223.395 92.320 -220.185 93.220 ;
        RECT -223.395 92.315 -222.045 92.320 ;
        RECT -221.535 92.315 -220.185 92.320 ;
        RECT -213.475 93.220 -212.125 93.225 ;
        RECT -211.615 93.220 -210.265 93.225 ;
        RECT -213.475 92.320 -210.265 93.220 ;
        RECT -213.475 92.315 -212.125 92.320 ;
        RECT -211.615 92.315 -210.265 92.320 ;
        RECT -203.555 93.220 -202.205 93.225 ;
        RECT -201.695 93.220 -200.345 93.225 ;
        RECT -203.555 92.320 -200.345 93.220 ;
        RECT -203.555 92.315 -202.205 92.320 ;
        RECT -201.695 92.315 -200.345 92.320 ;
        RECT -193.635 93.220 -192.285 93.225 ;
        RECT -191.775 93.220 -190.425 93.225 ;
        RECT -193.635 92.320 -190.425 93.220 ;
        RECT -193.635 92.315 -192.285 92.320 ;
        RECT -191.775 92.315 -190.425 92.320 ;
        RECT -183.715 93.220 -182.365 93.225 ;
        RECT -181.855 93.220 -180.505 93.225 ;
        RECT -183.715 92.320 -180.505 93.220 ;
        RECT -183.715 92.315 -182.365 92.320 ;
        RECT -181.855 92.315 -180.505 92.320 ;
        RECT -173.795 93.220 -172.445 93.225 ;
        RECT -171.935 93.220 -170.585 93.225 ;
        RECT -173.795 92.320 -170.585 93.220 ;
        RECT -173.795 92.315 -172.445 92.320 ;
        RECT -171.935 92.315 -170.585 92.320 ;
        RECT -163.875 93.220 -162.525 93.225 ;
        RECT -162.015 93.220 -160.665 93.225 ;
        RECT -163.875 92.320 -160.665 93.220 ;
        RECT -163.875 92.315 -162.525 92.320 ;
        RECT -162.015 92.315 -160.665 92.320 ;
        RECT -153.955 93.220 -152.605 93.225 ;
        RECT -152.095 93.220 -150.745 93.225 ;
        RECT -153.955 92.320 -150.745 93.220 ;
        RECT -153.955 92.315 -152.605 92.320 ;
        RECT -152.095 92.315 -150.745 92.320 ;
        RECT -144.035 93.220 -142.685 93.225 ;
        RECT -142.175 93.220 -140.825 93.225 ;
        RECT -144.035 92.320 -140.825 93.220 ;
        RECT -144.035 92.315 -142.685 92.320 ;
        RECT -142.175 92.315 -140.825 92.320 ;
        RECT -134.115 93.220 -132.765 93.225 ;
        RECT -132.255 93.220 -130.905 93.225 ;
        RECT -134.115 92.320 -130.905 93.220 ;
        RECT -134.115 92.315 -132.765 92.320 ;
        RECT -132.255 92.315 -130.905 92.320 ;
        RECT -124.195 93.220 -122.845 93.225 ;
        RECT -122.335 93.220 -120.985 93.225 ;
        RECT -124.195 92.320 -120.985 93.220 ;
        RECT -124.195 92.315 -122.845 92.320 ;
        RECT -122.335 92.315 -120.985 92.320 ;
        RECT -114.275 93.220 -112.925 93.225 ;
        RECT -112.415 93.220 -111.065 93.225 ;
        RECT -114.275 92.320 -111.065 93.220 ;
        RECT -114.275 92.315 -112.925 92.320 ;
        RECT -112.415 92.315 -111.065 92.320 ;
        RECT -104.355 93.220 -103.005 93.225 ;
        RECT -102.495 93.220 -101.145 93.225 ;
        RECT -104.355 92.320 -101.145 93.220 ;
        RECT -104.355 92.315 -103.005 92.320 ;
        RECT -102.495 92.315 -101.145 92.320 ;
        RECT -94.435 93.220 -93.085 93.225 ;
        RECT -92.575 93.220 -91.225 93.225 ;
        RECT -94.435 92.320 -91.225 93.220 ;
        RECT -94.435 92.315 -93.085 92.320 ;
        RECT -92.575 92.315 -91.225 92.320 ;
        RECT -84.515 93.220 -83.165 93.225 ;
        RECT -82.655 93.220 -81.305 93.225 ;
        RECT -84.515 92.320 -81.305 93.220 ;
        RECT -84.515 92.315 -83.165 92.320 ;
        RECT -82.655 92.315 -81.305 92.320 ;
        RECT -74.595 93.220 -73.245 93.225 ;
        RECT -72.735 93.220 -71.385 93.225 ;
        RECT -74.595 92.320 -71.385 93.220 ;
        RECT -74.595 92.315 -73.245 92.320 ;
        RECT -72.735 92.315 -71.385 92.320 ;
        RECT -64.675 93.220 -63.325 93.225 ;
        RECT -62.815 93.220 -61.465 93.225 ;
        RECT -64.675 92.320 -61.465 93.220 ;
        RECT -64.675 92.315 -63.325 92.320 ;
        RECT -62.815 92.315 -61.465 92.320 ;
        RECT -54.755 93.220 -53.405 93.225 ;
        RECT -52.895 93.220 -51.545 93.225 ;
        RECT -54.755 92.320 -51.545 93.220 ;
        RECT -54.755 92.315 -53.405 92.320 ;
        RECT -52.895 92.315 -51.545 92.320 ;
        RECT -44.835 93.220 -43.485 93.225 ;
        RECT -42.975 93.220 -41.625 93.225 ;
        RECT -44.835 92.320 -41.625 93.220 ;
        RECT -44.835 92.315 -43.485 92.320 ;
        RECT -42.975 92.315 -41.625 92.320 ;
        RECT -34.915 93.220 -33.565 93.225 ;
        RECT -33.055 93.220 -31.705 93.225 ;
        RECT -34.915 92.320 -31.705 93.220 ;
        RECT -34.915 92.315 -33.565 92.320 ;
        RECT -33.055 92.315 -31.705 92.320 ;
        RECT -24.995 93.220 -23.645 93.225 ;
        RECT -23.135 93.220 -21.785 93.225 ;
        RECT -24.995 92.320 -21.785 93.220 ;
        RECT -24.995 92.315 -23.645 92.320 ;
        RECT -23.135 92.315 -21.785 92.320 ;
        RECT -15.075 93.220 -13.725 93.225 ;
        RECT -13.215 93.220 -11.865 93.225 ;
        RECT -15.075 92.320 -11.865 93.220 ;
        RECT -15.075 92.315 -13.725 92.320 ;
        RECT -13.215 92.315 -11.865 92.320 ;
        RECT -5.155 93.220 -3.805 93.225 ;
        RECT -3.295 93.220 -1.945 93.225 ;
        RECT -5.155 92.320 -1.945 93.220 ;
        RECT -5.155 92.315 -3.805 92.320 ;
        RECT -3.295 92.315 -1.945 92.320 ;
        RECT 4.765 93.220 6.115 93.225 ;
        RECT 6.625 93.220 7.975 93.225 ;
        RECT 4.765 92.320 7.975 93.220 ;
        RECT 4.765 92.315 6.115 92.320 ;
        RECT 6.625 92.315 7.975 92.320 ;
        RECT 14.685 93.220 16.035 93.225 ;
        RECT 16.545 93.220 17.895 93.225 ;
        RECT 14.685 92.320 17.895 93.220 ;
        RECT 14.685 92.315 16.035 92.320 ;
        RECT 16.545 92.315 17.895 92.320 ;
        RECT -287.875 91.620 -286.525 91.625 ;
        RECT -286.015 91.620 -284.665 91.625 ;
        RECT -287.875 90.720 -284.665 91.620 ;
        RECT -287.875 90.715 -286.525 90.720 ;
        RECT -286.015 90.715 -284.665 90.720 ;
        RECT -277.955 91.620 -276.605 91.625 ;
        RECT -276.095 91.620 -274.745 91.625 ;
        RECT -277.955 90.720 -274.745 91.620 ;
        RECT -277.955 90.715 -276.605 90.720 ;
        RECT -276.095 90.715 -274.745 90.720 ;
        RECT -268.035 91.620 -266.685 91.625 ;
        RECT -266.175 91.620 -264.825 91.625 ;
        RECT -268.035 90.720 -264.825 91.620 ;
        RECT -268.035 90.715 -266.685 90.720 ;
        RECT -266.175 90.715 -264.825 90.720 ;
        RECT -258.115 91.620 -256.765 91.625 ;
        RECT -256.255 91.620 -254.905 91.625 ;
        RECT -258.115 90.720 -254.905 91.620 ;
        RECT -258.115 90.715 -256.765 90.720 ;
        RECT -256.255 90.715 -254.905 90.720 ;
        RECT -248.195 91.620 -246.845 91.625 ;
        RECT -246.335 91.620 -244.985 91.625 ;
        RECT -248.195 90.720 -244.985 91.620 ;
        RECT -248.195 90.715 -246.845 90.720 ;
        RECT -246.335 90.715 -244.985 90.720 ;
        RECT -238.275 91.620 -236.925 91.625 ;
        RECT -236.415 91.620 -235.065 91.625 ;
        RECT -238.275 90.720 -235.065 91.620 ;
        RECT -238.275 90.715 -236.925 90.720 ;
        RECT -236.415 90.715 -235.065 90.720 ;
        RECT -228.355 91.620 -227.005 91.625 ;
        RECT -226.495 91.620 -225.145 91.625 ;
        RECT -228.355 90.720 -225.145 91.620 ;
        RECT -228.355 90.715 -227.005 90.720 ;
        RECT -226.495 90.715 -225.145 90.720 ;
        RECT -218.435 91.620 -217.085 91.625 ;
        RECT -216.575 91.620 -215.225 91.625 ;
        RECT -218.435 90.720 -215.225 91.620 ;
        RECT -218.435 90.715 -217.085 90.720 ;
        RECT -216.575 90.715 -215.225 90.720 ;
        RECT -208.515 91.620 -207.165 91.625 ;
        RECT -206.655 91.620 -205.305 91.625 ;
        RECT -208.515 90.720 -205.305 91.620 ;
        RECT -208.515 90.715 -207.165 90.720 ;
        RECT -206.655 90.715 -205.305 90.720 ;
        RECT -198.595 91.620 -197.245 91.625 ;
        RECT -196.735 91.620 -195.385 91.625 ;
        RECT -198.595 90.720 -195.385 91.620 ;
        RECT -198.595 90.715 -197.245 90.720 ;
        RECT -196.735 90.715 -195.385 90.720 ;
        RECT -188.675 91.620 -187.325 91.625 ;
        RECT -186.815 91.620 -185.465 91.625 ;
        RECT -188.675 90.720 -185.465 91.620 ;
        RECT -188.675 90.715 -187.325 90.720 ;
        RECT -186.815 90.715 -185.465 90.720 ;
        RECT -178.755 91.620 -177.405 91.625 ;
        RECT -176.895 91.620 -175.545 91.625 ;
        RECT -178.755 90.720 -175.545 91.620 ;
        RECT -178.755 90.715 -177.405 90.720 ;
        RECT -176.895 90.715 -175.545 90.720 ;
        RECT -168.835 91.620 -167.485 91.625 ;
        RECT -166.975 91.620 -165.625 91.625 ;
        RECT -168.835 90.720 -165.625 91.620 ;
        RECT -168.835 90.715 -167.485 90.720 ;
        RECT -166.975 90.715 -165.625 90.720 ;
        RECT -158.915 91.620 -157.565 91.625 ;
        RECT -157.055 91.620 -155.705 91.625 ;
        RECT -158.915 90.720 -155.705 91.620 ;
        RECT -158.915 90.715 -157.565 90.720 ;
        RECT -157.055 90.715 -155.705 90.720 ;
        RECT -148.995 91.620 -147.645 91.625 ;
        RECT -147.135 91.620 -145.785 91.625 ;
        RECT -148.995 90.720 -145.785 91.620 ;
        RECT -148.995 90.715 -147.645 90.720 ;
        RECT -147.135 90.715 -145.785 90.720 ;
        RECT -139.075 91.620 -137.725 91.625 ;
        RECT -137.215 91.620 -135.865 91.625 ;
        RECT -139.075 90.720 -135.865 91.620 ;
        RECT -139.075 90.715 -137.725 90.720 ;
        RECT -137.215 90.715 -135.865 90.720 ;
        RECT -129.155 91.620 -127.805 91.625 ;
        RECT -127.295 91.620 -125.945 91.625 ;
        RECT -129.155 90.720 -125.945 91.620 ;
        RECT -129.155 90.715 -127.805 90.720 ;
        RECT -127.295 90.715 -125.945 90.720 ;
        RECT -119.235 91.620 -117.885 91.625 ;
        RECT -117.375 91.620 -116.025 91.625 ;
        RECT -119.235 90.720 -116.025 91.620 ;
        RECT -119.235 90.715 -117.885 90.720 ;
        RECT -117.375 90.715 -116.025 90.720 ;
        RECT -109.315 91.620 -107.965 91.625 ;
        RECT -107.455 91.620 -106.105 91.625 ;
        RECT -109.315 90.720 -106.105 91.620 ;
        RECT -109.315 90.715 -107.965 90.720 ;
        RECT -107.455 90.715 -106.105 90.720 ;
        RECT -99.395 91.620 -98.045 91.625 ;
        RECT -97.535 91.620 -96.185 91.625 ;
        RECT -99.395 90.720 -96.185 91.620 ;
        RECT -99.395 90.715 -98.045 90.720 ;
        RECT -97.535 90.715 -96.185 90.720 ;
        RECT -89.475 91.620 -88.125 91.625 ;
        RECT -87.615 91.620 -86.265 91.625 ;
        RECT -89.475 90.720 -86.265 91.620 ;
        RECT -89.475 90.715 -88.125 90.720 ;
        RECT -87.615 90.715 -86.265 90.720 ;
        RECT -79.555 91.620 -78.205 91.625 ;
        RECT -77.695 91.620 -76.345 91.625 ;
        RECT -79.555 90.720 -76.345 91.620 ;
        RECT -79.555 90.715 -78.205 90.720 ;
        RECT -77.695 90.715 -76.345 90.720 ;
        RECT -69.635 91.620 -68.285 91.625 ;
        RECT -67.775 91.620 -66.425 91.625 ;
        RECT -69.635 90.720 -66.425 91.620 ;
        RECT -69.635 90.715 -68.285 90.720 ;
        RECT -67.775 90.715 -66.425 90.720 ;
        RECT -59.715 91.620 -58.365 91.625 ;
        RECT -57.855 91.620 -56.505 91.625 ;
        RECT -59.715 90.720 -56.505 91.620 ;
        RECT -59.715 90.715 -58.365 90.720 ;
        RECT -57.855 90.715 -56.505 90.720 ;
        RECT -49.795 91.620 -48.445 91.625 ;
        RECT -47.935 91.620 -46.585 91.625 ;
        RECT -49.795 90.720 -46.585 91.620 ;
        RECT -49.795 90.715 -48.445 90.720 ;
        RECT -47.935 90.715 -46.585 90.720 ;
        RECT -39.875 91.620 -38.525 91.625 ;
        RECT -38.015 91.620 -36.665 91.625 ;
        RECT -39.875 90.720 -36.665 91.620 ;
        RECT -39.875 90.715 -38.525 90.720 ;
        RECT -38.015 90.715 -36.665 90.720 ;
        RECT -29.955 91.620 -28.605 91.625 ;
        RECT -28.095 91.620 -26.745 91.625 ;
        RECT -29.955 90.720 -26.745 91.620 ;
        RECT -29.955 90.715 -28.605 90.720 ;
        RECT -28.095 90.715 -26.745 90.720 ;
        RECT -20.035 91.620 -18.685 91.625 ;
        RECT -18.175 91.620 -16.825 91.625 ;
        RECT -20.035 90.720 -16.825 91.620 ;
        RECT -20.035 90.715 -18.685 90.720 ;
        RECT -18.175 90.715 -16.825 90.720 ;
        RECT -10.115 91.620 -8.765 91.625 ;
        RECT -8.255 91.620 -6.905 91.625 ;
        RECT -10.115 90.720 -6.905 91.620 ;
        RECT -10.115 90.715 -8.765 90.720 ;
        RECT -8.255 90.715 -6.905 90.720 ;
        RECT -0.195 91.620 1.155 91.625 ;
        RECT 1.665 91.620 3.015 91.625 ;
        RECT -0.195 90.720 3.015 91.620 ;
        RECT -0.195 90.715 1.155 90.720 ;
        RECT 1.665 90.715 3.015 90.720 ;
        RECT 9.725 91.620 11.075 91.625 ;
        RECT 11.585 91.620 12.935 91.625 ;
        RECT 9.725 90.720 12.935 91.620 ;
        RECT 9.725 90.715 11.075 90.720 ;
        RECT 11.585 90.715 12.935 90.720 ;
        RECT 19.645 91.620 20.995 91.625 ;
        RECT 21.505 91.620 22.855 91.625 ;
        RECT 19.645 90.720 22.855 91.620 ;
        RECT 19.645 90.715 20.995 90.720 ;
        RECT 21.505 90.715 22.855 90.720 ;
        RECT -286.810 90.525 -286.640 90.715 ;
        RECT -285.900 90.525 -285.730 90.715 ;
        RECT -276.890 90.525 -276.720 90.715 ;
        RECT -275.980 90.525 -275.810 90.715 ;
        RECT -266.970 90.525 -266.800 90.715 ;
        RECT -266.060 90.525 -265.890 90.715 ;
        RECT -257.050 90.525 -256.880 90.715 ;
        RECT -256.140 90.525 -255.970 90.715 ;
        RECT -247.130 90.525 -246.960 90.715 ;
        RECT -246.220 90.525 -246.050 90.715 ;
        RECT -237.210 90.525 -237.040 90.715 ;
        RECT -236.300 90.525 -236.130 90.715 ;
        RECT -227.290 90.525 -227.120 90.715 ;
        RECT -226.380 90.525 -226.210 90.715 ;
        RECT -217.370 90.525 -217.200 90.715 ;
        RECT -216.460 90.525 -216.290 90.715 ;
        RECT -207.450 90.525 -207.280 90.715 ;
        RECT -206.540 90.525 -206.370 90.715 ;
        RECT -197.530 90.525 -197.360 90.715 ;
        RECT -196.620 90.525 -196.450 90.715 ;
        RECT -187.610 90.525 -187.440 90.715 ;
        RECT -186.700 90.525 -186.530 90.715 ;
        RECT -177.690 90.525 -177.520 90.715 ;
        RECT -176.780 90.525 -176.610 90.715 ;
        RECT -167.770 90.525 -167.600 90.715 ;
        RECT -166.860 90.525 -166.690 90.715 ;
        RECT -157.850 90.525 -157.680 90.715 ;
        RECT -156.940 90.525 -156.770 90.715 ;
        RECT -147.930 90.525 -147.760 90.715 ;
        RECT -147.020 90.525 -146.850 90.715 ;
        RECT -138.010 90.525 -137.840 90.715 ;
        RECT -137.100 90.525 -136.930 90.715 ;
        RECT -128.090 90.525 -127.920 90.715 ;
        RECT -127.180 90.525 -127.010 90.715 ;
        RECT -118.170 90.525 -118.000 90.715 ;
        RECT -117.260 90.525 -117.090 90.715 ;
        RECT -108.250 90.525 -108.080 90.715 ;
        RECT -107.340 90.525 -107.170 90.715 ;
        RECT -98.330 90.525 -98.160 90.715 ;
        RECT -97.420 90.525 -97.250 90.715 ;
        RECT -88.410 90.525 -88.240 90.715 ;
        RECT -87.500 90.525 -87.330 90.715 ;
        RECT -78.490 90.525 -78.320 90.715 ;
        RECT -77.580 90.525 -77.410 90.715 ;
        RECT -68.570 90.525 -68.400 90.715 ;
        RECT -67.660 90.525 -67.490 90.715 ;
        RECT -58.650 90.525 -58.480 90.715 ;
        RECT -57.740 90.525 -57.570 90.715 ;
        RECT -48.730 90.525 -48.560 90.715 ;
        RECT -47.820 90.525 -47.650 90.715 ;
        RECT -38.810 90.525 -38.640 90.715 ;
        RECT -37.900 90.525 -37.730 90.715 ;
        RECT -28.890 90.525 -28.720 90.715 ;
        RECT -27.980 90.525 -27.810 90.715 ;
        RECT -18.970 90.525 -18.800 90.715 ;
        RECT -18.060 90.525 -17.890 90.715 ;
        RECT -9.050 90.525 -8.880 90.715 ;
        RECT -8.140 90.525 -7.970 90.715 ;
        RECT 0.870 90.525 1.040 90.715 ;
        RECT 1.780 90.525 1.950 90.715 ;
        RECT 10.790 90.525 10.960 90.715 ;
        RECT 11.700 90.525 11.870 90.715 ;
        RECT 20.710 90.525 20.880 90.715 ;
        RECT 21.620 90.525 21.790 90.715 ;
        RECT -281.525 90.180 -281.095 90.195 ;
        RECT -271.605 90.180 -271.175 90.195 ;
        RECT -261.685 90.180 -261.255 90.195 ;
        RECT -251.765 90.180 -251.335 90.195 ;
        RECT -241.845 90.180 -241.415 90.195 ;
        RECT -231.925 90.180 -231.495 90.195 ;
        RECT -222.005 90.180 -221.575 90.195 ;
        RECT -212.085 90.180 -211.655 90.195 ;
        RECT -202.165 90.180 -201.735 90.195 ;
        RECT -192.245 90.180 -191.815 90.195 ;
        RECT -182.325 90.180 -181.895 90.195 ;
        RECT -172.405 90.180 -171.975 90.195 ;
        RECT -162.485 90.180 -162.055 90.195 ;
        RECT -152.565 90.180 -152.135 90.195 ;
        RECT -142.645 90.180 -142.215 90.195 ;
        RECT -132.725 90.180 -132.295 90.195 ;
        RECT -122.805 90.180 -122.375 90.195 ;
        RECT -112.885 90.180 -112.455 90.195 ;
        RECT -102.965 90.180 -102.535 90.195 ;
        RECT -93.045 90.180 -92.615 90.195 ;
        RECT -83.125 90.180 -82.695 90.195 ;
        RECT -73.205 90.180 -72.775 90.195 ;
        RECT -63.285 90.180 -62.855 90.195 ;
        RECT -53.365 90.180 -52.935 90.195 ;
        RECT -43.445 90.180 -43.015 90.195 ;
        RECT -33.525 90.180 -33.095 90.195 ;
        RECT -23.605 90.180 -23.175 90.195 ;
        RECT -13.685 90.180 -13.255 90.195 ;
        RECT -3.765 90.180 -3.335 90.195 ;
        RECT 6.155 90.180 6.585 90.195 ;
        RECT 16.075 90.180 16.505 90.195 ;
        RECT -283.360 90.175 -279.420 90.180 ;
        RECT -273.400 90.175 -269.380 90.180 ;
        RECT -263.520 90.175 -259.580 90.180 ;
        RECT -283.965 88.820 -278.655 90.175 ;
        RECT -283.965 88.805 -283.185 88.820 ;
        RECT -279.435 88.805 -278.655 88.820 ;
        RECT -274.045 88.805 -268.735 90.175 ;
        RECT -264.125 88.820 -258.815 90.175 ;
        RECT -264.125 88.805 -263.345 88.820 ;
        RECT -259.595 88.805 -258.815 88.820 ;
        RECT -254.205 90.170 -253.425 90.175 ;
        RECT -253.360 90.170 -249.910 90.180 ;
        RECT -243.680 90.175 -239.740 90.180 ;
        RECT -233.720 90.175 -229.700 90.180 ;
        RECT -223.840 90.175 -219.900 90.180 ;
        RECT -213.840 90.175 -209.770 90.180 ;
        RECT -204.000 90.175 -200.060 90.180 ;
        RECT -194.040 90.175 -190.020 90.180 ;
        RECT -184.160 90.175 -180.220 90.180 ;
        RECT -249.675 90.170 -248.895 90.175 ;
        RECT -254.205 88.805 -248.895 90.170 ;
        RECT -244.285 88.820 -238.975 90.175 ;
        RECT -244.285 88.805 -243.505 88.820 ;
        RECT -239.755 88.805 -238.975 88.820 ;
        RECT -234.365 88.805 -229.055 90.175 ;
        RECT -224.445 88.820 -219.135 90.175 ;
        RECT -224.445 88.805 -223.665 88.820 ;
        RECT -219.915 88.805 -219.135 88.820 ;
        RECT -214.525 88.810 -209.215 90.175 ;
        RECT -214.525 88.805 -213.745 88.810 ;
        RECT -209.995 88.805 -209.215 88.810 ;
        RECT -204.605 88.820 -199.295 90.175 ;
        RECT -204.605 88.805 -203.825 88.820 ;
        RECT -200.075 88.805 -199.295 88.820 ;
        RECT -194.685 88.805 -189.375 90.175 ;
        RECT -184.765 88.820 -179.455 90.175 ;
        RECT -184.765 88.805 -183.985 88.820 ;
        RECT -180.235 88.805 -179.455 88.820 ;
        RECT -174.845 90.170 -174.065 90.175 ;
        RECT -174.000 90.170 -170.550 90.180 ;
        RECT -164.320 90.175 -160.380 90.180 ;
        RECT -154.360 90.175 -150.340 90.180 ;
        RECT -144.480 90.175 -140.540 90.180 ;
        RECT -134.440 90.175 -130.500 90.180 ;
        RECT -124.640 90.175 -120.700 90.180 ;
        RECT -114.680 90.175 -110.660 90.180 ;
        RECT -104.800 90.175 -100.860 90.180 ;
        RECT -170.315 90.170 -169.535 90.175 ;
        RECT -174.845 88.805 -169.535 90.170 ;
        RECT -164.925 88.820 -159.615 90.175 ;
        RECT -164.925 88.805 -164.145 88.820 ;
        RECT -160.395 88.805 -159.615 88.820 ;
        RECT -155.005 88.805 -149.695 90.175 ;
        RECT -145.085 88.820 -139.775 90.175 ;
        RECT -145.085 88.805 -144.305 88.820 ;
        RECT -140.555 88.805 -139.775 88.820 ;
        RECT -135.165 88.820 -129.855 90.175 ;
        RECT -135.165 88.805 -134.385 88.820 ;
        RECT -130.635 88.805 -129.855 88.820 ;
        RECT -125.245 88.820 -119.935 90.175 ;
        RECT -125.245 88.805 -124.465 88.820 ;
        RECT -120.715 88.805 -119.935 88.820 ;
        RECT -115.325 88.805 -110.015 90.175 ;
        RECT -105.405 88.820 -100.095 90.175 ;
        RECT -105.405 88.805 -104.625 88.820 ;
        RECT -100.875 88.805 -100.095 88.820 ;
        RECT -95.485 90.170 -94.705 90.175 ;
        RECT -94.640 90.170 -91.190 90.180 ;
        RECT -84.960 90.175 -81.020 90.180 ;
        RECT -75.000 90.175 -70.980 90.180 ;
        RECT -65.120 90.175 -61.180 90.180 ;
        RECT -55.120 90.175 -51.050 90.180 ;
        RECT -45.280 90.175 -41.340 90.180 ;
        RECT -35.320 90.175 -31.300 90.180 ;
        RECT -25.440 90.175 -21.500 90.180 ;
        RECT -90.955 90.170 -90.175 90.175 ;
        RECT -95.485 88.805 -90.175 90.170 ;
        RECT -85.565 88.820 -80.255 90.175 ;
        RECT -85.565 88.805 -84.785 88.820 ;
        RECT -81.035 88.805 -80.255 88.820 ;
        RECT -75.645 88.805 -70.335 90.175 ;
        RECT -65.725 88.820 -60.415 90.175 ;
        RECT -65.725 88.805 -64.945 88.820 ;
        RECT -61.195 88.805 -60.415 88.820 ;
        RECT -55.805 88.810 -50.495 90.175 ;
        RECT -55.805 88.805 -55.025 88.810 ;
        RECT -51.275 88.805 -50.495 88.810 ;
        RECT -45.885 88.820 -40.575 90.175 ;
        RECT -45.885 88.805 -45.105 88.820 ;
        RECT -41.355 88.805 -40.575 88.820 ;
        RECT -35.965 88.805 -30.655 90.175 ;
        RECT -26.045 88.820 -20.735 90.175 ;
        RECT -26.045 88.805 -25.265 88.820 ;
        RECT -21.515 88.805 -20.735 88.820 ;
        RECT -16.125 90.170 -15.345 90.175 ;
        RECT -15.280 90.170 -11.830 90.180 ;
        RECT -5.600 90.175 -1.660 90.180 ;
        RECT 4.360 90.175 8.380 90.180 ;
        RECT 14.240 90.175 18.180 90.180 ;
        RECT -11.595 90.170 -10.815 90.175 ;
        RECT -16.125 88.805 -10.815 90.170 ;
        RECT -6.205 88.820 -0.895 90.175 ;
        RECT -6.205 88.805 -5.425 88.820 ;
        RECT -1.675 88.805 -0.895 88.820 ;
        RECT 3.715 88.805 9.025 90.175 ;
        RECT 13.635 88.820 18.945 90.175 ;
        RECT 13.635 88.805 14.415 88.820 ;
        RECT 18.165 88.805 18.945 88.820 ;
        RECT -273.400 88.800 -269.380 88.805 ;
        RECT -253.480 88.800 -249.640 88.805 ;
        RECT -233.720 88.800 -229.700 88.805 ;
        RECT -194.040 88.800 -190.020 88.805 ;
        RECT -174.120 88.800 -170.280 88.805 ;
        RECT -154.360 88.800 -150.340 88.805 ;
        RECT -114.680 88.800 -110.660 88.805 ;
        RECT -94.760 88.800 -90.920 88.805 ;
        RECT -75.000 88.800 -70.980 88.805 ;
        RECT -35.320 88.800 -31.300 88.805 ;
        RECT -15.400 88.800 -11.560 88.805 ;
        RECT 4.360 88.800 8.380 88.805 ;
        RECT -290.240 11.085 -286.280 11.090 ;
        RECT -280.320 11.085 -276.360 11.090 ;
        RECT -270.400 11.085 -266.440 11.090 ;
        RECT -260.480 11.085 -256.520 11.090 ;
        RECT -250.560 11.085 -246.600 11.090 ;
        RECT -240.640 11.085 -236.680 11.090 ;
        RECT -230.720 11.085 -226.760 11.090 ;
        RECT -220.800 11.085 -216.840 11.090 ;
        RECT -210.880 11.085 -206.920 11.090 ;
        RECT -200.960 11.085 -197.000 11.090 ;
        RECT -191.040 11.085 -187.080 11.090 ;
        RECT -181.120 11.085 -177.160 11.090 ;
        RECT -171.200 11.085 -167.240 11.090 ;
        RECT -161.280 11.085 -157.320 11.090 ;
        RECT -151.360 11.085 -147.400 11.090 ;
        RECT -141.440 11.085 -137.480 11.090 ;
        RECT -131.520 11.085 -127.560 11.090 ;
        RECT -121.600 11.085 -117.640 11.090 ;
        RECT -111.680 11.085 -107.720 11.090 ;
        RECT -101.760 11.085 -97.800 11.090 ;
        RECT -91.840 11.085 -87.880 11.090 ;
        RECT -81.920 11.085 -77.960 11.090 ;
        RECT -72.000 11.085 -68.040 11.090 ;
        RECT -62.080 11.085 -58.120 11.090 ;
        RECT -52.160 11.085 -48.200 11.090 ;
        RECT -42.240 11.085 -38.280 11.090 ;
        RECT -32.320 11.085 -28.360 11.090 ;
        RECT -22.400 11.085 -18.440 11.090 ;
        RECT -12.480 11.085 -8.520 11.090 ;
        RECT -2.560 11.085 1.400 11.090 ;
        RECT 7.360 11.085 11.320 11.090 ;
        RECT 17.280 11.085 21.240 11.090 ;
        RECT -290.945 9.715 -285.635 11.085 ;
        RECT -281.025 9.715 -275.715 11.085 ;
        RECT -271.105 9.715 -265.795 11.085 ;
        RECT -261.185 9.715 -255.875 11.085 ;
        RECT -251.265 9.715 -245.955 11.085 ;
        RECT -241.345 9.715 -236.035 11.085 ;
        RECT -231.425 9.715 -226.115 11.085 ;
        RECT -221.505 9.715 -216.195 11.085 ;
        RECT -211.585 9.715 -206.275 11.085 ;
        RECT -201.665 9.715 -196.355 11.085 ;
        RECT -191.745 9.715 -186.435 11.085 ;
        RECT -181.825 9.715 -176.515 11.085 ;
        RECT -171.905 9.715 -166.595 11.085 ;
        RECT -161.985 9.715 -156.675 11.085 ;
        RECT -152.065 9.715 -146.755 11.085 ;
        RECT -142.145 9.715 -136.835 11.085 ;
        RECT -132.225 9.715 -126.915 11.085 ;
        RECT -122.305 9.715 -116.995 11.085 ;
        RECT -112.385 9.715 -107.075 11.085 ;
        RECT -102.465 9.715 -97.155 11.085 ;
        RECT -92.545 9.715 -87.235 11.085 ;
        RECT -82.625 9.715 -77.315 11.085 ;
        RECT -72.705 9.715 -67.395 11.085 ;
        RECT -62.785 9.715 -57.475 11.085 ;
        RECT -52.865 9.715 -47.555 11.085 ;
        RECT -42.945 9.715 -37.635 11.085 ;
        RECT -33.025 9.715 -27.715 11.085 ;
        RECT -23.105 9.715 -17.795 11.085 ;
        RECT -13.185 9.715 -7.875 11.085 ;
        RECT -3.265 9.715 2.045 11.085 ;
        RECT 6.655 9.715 11.965 11.085 ;
        RECT 16.575 9.715 21.885 11.085 ;
        RECT -290.240 9.710 -286.280 9.715 ;
        RECT -280.320 9.710 -276.360 9.715 ;
        RECT -270.400 9.710 -266.440 9.715 ;
        RECT -260.480 9.710 -256.520 9.715 ;
        RECT -250.560 9.710 -246.600 9.715 ;
        RECT -240.640 9.710 -236.680 9.715 ;
        RECT -230.720 9.710 -226.760 9.715 ;
        RECT -220.800 9.710 -216.840 9.715 ;
        RECT -210.880 9.710 -206.920 9.715 ;
        RECT -200.960 9.710 -197.000 9.715 ;
        RECT -191.040 9.710 -187.080 9.715 ;
        RECT -181.120 9.710 -177.160 9.715 ;
        RECT -171.200 9.710 -167.240 9.715 ;
        RECT -161.280 9.710 -157.320 9.715 ;
        RECT -151.360 9.710 -147.400 9.715 ;
        RECT -141.440 9.710 -137.480 9.715 ;
        RECT -131.520 9.710 -127.560 9.715 ;
        RECT -121.600 9.710 -117.640 9.715 ;
        RECT -111.680 9.710 -107.720 9.715 ;
        RECT -101.760 9.710 -97.800 9.715 ;
        RECT -91.840 9.710 -87.880 9.715 ;
        RECT -81.920 9.710 -77.960 9.715 ;
        RECT -72.000 9.710 -68.040 9.715 ;
        RECT -62.080 9.710 -58.120 9.715 ;
        RECT -52.160 9.710 -48.200 9.715 ;
        RECT -42.240 9.710 -38.280 9.715 ;
        RECT -32.320 9.710 -28.360 9.715 ;
        RECT -22.400 9.710 -18.440 9.715 ;
        RECT -12.480 9.710 -8.520 9.715 ;
        RECT -2.560 9.710 1.400 9.715 ;
        RECT 7.360 9.710 11.320 9.715 ;
        RECT 17.280 9.710 21.240 9.715 ;
        RECT -283.870 9.175 -283.700 9.365 ;
        RECT -282.960 9.175 -282.790 9.365 ;
        RECT -273.950 9.175 -273.780 9.365 ;
        RECT -273.040 9.175 -272.870 9.365 ;
        RECT -264.030 9.175 -263.860 9.365 ;
        RECT -263.120 9.175 -262.950 9.365 ;
        RECT -254.110 9.175 -253.940 9.365 ;
        RECT -253.200 9.175 -253.030 9.365 ;
        RECT -244.190 9.175 -244.020 9.365 ;
        RECT -243.280 9.175 -243.110 9.365 ;
        RECT -234.270 9.175 -234.100 9.365 ;
        RECT -233.360 9.175 -233.190 9.365 ;
        RECT -224.350 9.175 -224.180 9.365 ;
        RECT -223.440 9.175 -223.270 9.365 ;
        RECT -214.430 9.175 -214.260 9.365 ;
        RECT -213.520 9.175 -213.350 9.365 ;
        RECT -204.510 9.175 -204.340 9.365 ;
        RECT -203.600 9.175 -203.430 9.365 ;
        RECT -194.590 9.175 -194.420 9.365 ;
        RECT -193.680 9.175 -193.510 9.365 ;
        RECT -184.670 9.175 -184.500 9.365 ;
        RECT -183.760 9.175 -183.590 9.365 ;
        RECT -174.750 9.175 -174.580 9.365 ;
        RECT -173.840 9.175 -173.670 9.365 ;
        RECT -164.830 9.175 -164.660 9.365 ;
        RECT -163.920 9.175 -163.750 9.365 ;
        RECT -154.910 9.175 -154.740 9.365 ;
        RECT -154.000 9.175 -153.830 9.365 ;
        RECT -144.990 9.175 -144.820 9.365 ;
        RECT -144.080 9.175 -143.910 9.365 ;
        RECT -135.070 9.175 -134.900 9.365 ;
        RECT -134.160 9.175 -133.990 9.365 ;
        RECT -125.150 9.175 -124.980 9.365 ;
        RECT -124.240 9.175 -124.070 9.365 ;
        RECT -115.230 9.175 -115.060 9.365 ;
        RECT -114.320 9.175 -114.150 9.365 ;
        RECT -105.310 9.175 -105.140 9.365 ;
        RECT -104.400 9.175 -104.230 9.365 ;
        RECT -95.390 9.175 -95.220 9.365 ;
        RECT -94.480 9.175 -94.310 9.365 ;
        RECT -85.470 9.175 -85.300 9.365 ;
        RECT -84.560 9.175 -84.390 9.365 ;
        RECT -75.550 9.175 -75.380 9.365 ;
        RECT -74.640 9.175 -74.470 9.365 ;
        RECT -65.630 9.175 -65.460 9.365 ;
        RECT -64.720 9.175 -64.550 9.365 ;
        RECT -55.710 9.175 -55.540 9.365 ;
        RECT -54.800 9.175 -54.630 9.365 ;
        RECT -45.790 9.175 -45.620 9.365 ;
        RECT -44.880 9.175 -44.710 9.365 ;
        RECT -35.870 9.175 -35.700 9.365 ;
        RECT -34.960 9.175 -34.790 9.365 ;
        RECT -25.950 9.175 -25.780 9.365 ;
        RECT -25.040 9.175 -24.870 9.365 ;
        RECT -16.030 9.175 -15.860 9.365 ;
        RECT -15.120 9.175 -14.950 9.365 ;
        RECT -6.110 9.175 -5.940 9.365 ;
        RECT -5.200 9.175 -5.030 9.365 ;
        RECT 3.810 9.175 3.980 9.365 ;
        RECT 4.720 9.175 4.890 9.365 ;
        RECT 13.730 9.175 13.900 9.365 ;
        RECT 14.640 9.175 14.810 9.365 ;
        RECT -284.935 9.170 -283.585 9.175 ;
        RECT -283.075 9.170 -281.725 9.175 ;
        RECT -284.935 8.270 -281.725 9.170 ;
        RECT -284.935 8.265 -283.585 8.270 ;
        RECT -283.075 8.265 -281.725 8.270 ;
        RECT -275.015 9.170 -273.665 9.175 ;
        RECT -273.155 9.170 -271.805 9.175 ;
        RECT -275.015 8.270 -271.805 9.170 ;
        RECT -275.015 8.265 -273.665 8.270 ;
        RECT -273.155 8.265 -271.805 8.270 ;
        RECT -265.095 9.170 -263.745 9.175 ;
        RECT -263.235 9.170 -261.885 9.175 ;
        RECT -265.095 8.270 -261.885 9.170 ;
        RECT -265.095 8.265 -263.745 8.270 ;
        RECT -263.235 8.265 -261.885 8.270 ;
        RECT -255.175 9.170 -253.825 9.175 ;
        RECT -253.315 9.170 -251.965 9.175 ;
        RECT -255.175 8.270 -251.965 9.170 ;
        RECT -255.175 8.265 -253.825 8.270 ;
        RECT -253.315 8.265 -251.965 8.270 ;
        RECT -245.255 9.170 -243.905 9.175 ;
        RECT -243.395 9.170 -242.045 9.175 ;
        RECT -245.255 8.270 -242.045 9.170 ;
        RECT -245.255 8.265 -243.905 8.270 ;
        RECT -243.395 8.265 -242.045 8.270 ;
        RECT -235.335 9.170 -233.985 9.175 ;
        RECT -233.475 9.170 -232.125 9.175 ;
        RECT -235.335 8.270 -232.125 9.170 ;
        RECT -235.335 8.265 -233.985 8.270 ;
        RECT -233.475 8.265 -232.125 8.270 ;
        RECT -225.415 9.170 -224.065 9.175 ;
        RECT -223.555 9.170 -222.205 9.175 ;
        RECT -225.415 8.270 -222.205 9.170 ;
        RECT -225.415 8.265 -224.065 8.270 ;
        RECT -223.555 8.265 -222.205 8.270 ;
        RECT -215.495 9.170 -214.145 9.175 ;
        RECT -213.635 9.170 -212.285 9.175 ;
        RECT -215.495 8.270 -212.285 9.170 ;
        RECT -215.495 8.265 -214.145 8.270 ;
        RECT -213.635 8.265 -212.285 8.270 ;
        RECT -205.575 9.170 -204.225 9.175 ;
        RECT -203.715 9.170 -202.365 9.175 ;
        RECT -205.575 8.270 -202.365 9.170 ;
        RECT -205.575 8.265 -204.225 8.270 ;
        RECT -203.715 8.265 -202.365 8.270 ;
        RECT -195.655 9.170 -194.305 9.175 ;
        RECT -193.795 9.170 -192.445 9.175 ;
        RECT -195.655 8.270 -192.445 9.170 ;
        RECT -195.655 8.265 -194.305 8.270 ;
        RECT -193.795 8.265 -192.445 8.270 ;
        RECT -185.735 9.170 -184.385 9.175 ;
        RECT -183.875 9.170 -182.525 9.175 ;
        RECT -185.735 8.270 -182.525 9.170 ;
        RECT -185.735 8.265 -184.385 8.270 ;
        RECT -183.875 8.265 -182.525 8.270 ;
        RECT -175.815 9.170 -174.465 9.175 ;
        RECT -173.955 9.170 -172.605 9.175 ;
        RECT -175.815 8.270 -172.605 9.170 ;
        RECT -175.815 8.265 -174.465 8.270 ;
        RECT -173.955 8.265 -172.605 8.270 ;
        RECT -165.895 9.170 -164.545 9.175 ;
        RECT -164.035 9.170 -162.685 9.175 ;
        RECT -165.895 8.270 -162.685 9.170 ;
        RECT -165.895 8.265 -164.545 8.270 ;
        RECT -164.035 8.265 -162.685 8.270 ;
        RECT -155.975 9.170 -154.625 9.175 ;
        RECT -154.115 9.170 -152.765 9.175 ;
        RECT -155.975 8.270 -152.765 9.170 ;
        RECT -155.975 8.265 -154.625 8.270 ;
        RECT -154.115 8.265 -152.765 8.270 ;
        RECT -146.055 9.170 -144.705 9.175 ;
        RECT -144.195 9.170 -142.845 9.175 ;
        RECT -146.055 8.270 -142.845 9.170 ;
        RECT -146.055 8.265 -144.705 8.270 ;
        RECT -144.195 8.265 -142.845 8.270 ;
        RECT -136.135 9.170 -134.785 9.175 ;
        RECT -134.275 9.170 -132.925 9.175 ;
        RECT -136.135 8.270 -132.925 9.170 ;
        RECT -136.135 8.265 -134.785 8.270 ;
        RECT -134.275 8.265 -132.925 8.270 ;
        RECT -126.215 9.170 -124.865 9.175 ;
        RECT -124.355 9.170 -123.005 9.175 ;
        RECT -126.215 8.270 -123.005 9.170 ;
        RECT -126.215 8.265 -124.865 8.270 ;
        RECT -124.355 8.265 -123.005 8.270 ;
        RECT -116.295 9.170 -114.945 9.175 ;
        RECT -114.435 9.170 -113.085 9.175 ;
        RECT -116.295 8.270 -113.085 9.170 ;
        RECT -116.295 8.265 -114.945 8.270 ;
        RECT -114.435 8.265 -113.085 8.270 ;
        RECT -106.375 9.170 -105.025 9.175 ;
        RECT -104.515 9.170 -103.165 9.175 ;
        RECT -106.375 8.270 -103.165 9.170 ;
        RECT -106.375 8.265 -105.025 8.270 ;
        RECT -104.515 8.265 -103.165 8.270 ;
        RECT -96.455 9.170 -95.105 9.175 ;
        RECT -94.595 9.170 -93.245 9.175 ;
        RECT -96.455 8.270 -93.245 9.170 ;
        RECT -96.455 8.265 -95.105 8.270 ;
        RECT -94.595 8.265 -93.245 8.270 ;
        RECT -86.535 9.170 -85.185 9.175 ;
        RECT -84.675 9.170 -83.325 9.175 ;
        RECT -86.535 8.270 -83.325 9.170 ;
        RECT -86.535 8.265 -85.185 8.270 ;
        RECT -84.675 8.265 -83.325 8.270 ;
        RECT -76.615 9.170 -75.265 9.175 ;
        RECT -74.755 9.170 -73.405 9.175 ;
        RECT -76.615 8.270 -73.405 9.170 ;
        RECT -76.615 8.265 -75.265 8.270 ;
        RECT -74.755 8.265 -73.405 8.270 ;
        RECT -66.695 9.170 -65.345 9.175 ;
        RECT -64.835 9.170 -63.485 9.175 ;
        RECT -66.695 8.270 -63.485 9.170 ;
        RECT -66.695 8.265 -65.345 8.270 ;
        RECT -64.835 8.265 -63.485 8.270 ;
        RECT -56.775 9.170 -55.425 9.175 ;
        RECT -54.915 9.170 -53.565 9.175 ;
        RECT -56.775 8.270 -53.565 9.170 ;
        RECT -56.775 8.265 -55.425 8.270 ;
        RECT -54.915 8.265 -53.565 8.270 ;
        RECT -46.855 9.170 -45.505 9.175 ;
        RECT -44.995 9.170 -43.645 9.175 ;
        RECT -46.855 8.270 -43.645 9.170 ;
        RECT -46.855 8.265 -45.505 8.270 ;
        RECT -44.995 8.265 -43.645 8.270 ;
        RECT -36.935 9.170 -35.585 9.175 ;
        RECT -35.075 9.170 -33.725 9.175 ;
        RECT -36.935 8.270 -33.725 9.170 ;
        RECT -36.935 8.265 -35.585 8.270 ;
        RECT -35.075 8.265 -33.725 8.270 ;
        RECT -27.015 9.170 -25.665 9.175 ;
        RECT -25.155 9.170 -23.805 9.175 ;
        RECT -27.015 8.270 -23.805 9.170 ;
        RECT -27.015 8.265 -25.665 8.270 ;
        RECT -25.155 8.265 -23.805 8.270 ;
        RECT -17.095 9.170 -15.745 9.175 ;
        RECT -15.235 9.170 -13.885 9.175 ;
        RECT -17.095 8.270 -13.885 9.170 ;
        RECT -17.095 8.265 -15.745 8.270 ;
        RECT -15.235 8.265 -13.885 8.270 ;
        RECT -7.175 9.170 -5.825 9.175 ;
        RECT -5.315 9.170 -3.965 9.175 ;
        RECT -7.175 8.270 -3.965 9.170 ;
        RECT -7.175 8.265 -5.825 8.270 ;
        RECT -5.315 8.265 -3.965 8.270 ;
        RECT 2.745 9.170 4.095 9.175 ;
        RECT 4.605 9.170 5.955 9.175 ;
        RECT 2.745 8.270 5.955 9.170 ;
        RECT 2.745 8.265 4.095 8.270 ;
        RECT 4.605 8.265 5.955 8.270 ;
        RECT 12.665 9.170 14.015 9.175 ;
        RECT 14.525 9.170 15.875 9.175 ;
        RECT 12.665 8.270 15.875 9.170 ;
        RECT 12.665 8.265 14.015 8.270 ;
        RECT 14.525 8.265 15.875 8.270 ;
        RECT -289.895 7.570 -288.545 7.575 ;
        RECT -288.035 7.570 -286.685 7.575 ;
        RECT -289.895 6.670 -286.685 7.570 ;
        RECT -289.895 6.665 -288.545 6.670 ;
        RECT -288.035 6.665 -286.685 6.670 ;
        RECT -279.975 7.570 -278.625 7.575 ;
        RECT -278.115 7.570 -276.765 7.575 ;
        RECT -279.975 6.670 -276.765 7.570 ;
        RECT -279.975 6.665 -278.625 6.670 ;
        RECT -278.115 6.665 -276.765 6.670 ;
        RECT -270.055 7.570 -268.705 7.575 ;
        RECT -268.195 7.570 -266.845 7.575 ;
        RECT -270.055 6.670 -266.845 7.570 ;
        RECT -270.055 6.665 -268.705 6.670 ;
        RECT -268.195 6.665 -266.845 6.670 ;
        RECT -260.135 7.570 -258.785 7.575 ;
        RECT -258.275 7.570 -256.925 7.575 ;
        RECT -260.135 6.670 -256.925 7.570 ;
        RECT -260.135 6.665 -258.785 6.670 ;
        RECT -258.275 6.665 -256.925 6.670 ;
        RECT -250.215 7.570 -248.865 7.575 ;
        RECT -248.355 7.570 -247.005 7.575 ;
        RECT -250.215 6.670 -247.005 7.570 ;
        RECT -250.215 6.665 -248.865 6.670 ;
        RECT -248.355 6.665 -247.005 6.670 ;
        RECT -240.295 7.570 -238.945 7.575 ;
        RECT -238.435 7.570 -237.085 7.575 ;
        RECT -240.295 6.670 -237.085 7.570 ;
        RECT -240.295 6.665 -238.945 6.670 ;
        RECT -238.435 6.665 -237.085 6.670 ;
        RECT -230.375 7.570 -229.025 7.575 ;
        RECT -228.515 7.570 -227.165 7.575 ;
        RECT -230.375 6.670 -227.165 7.570 ;
        RECT -230.375 6.665 -229.025 6.670 ;
        RECT -228.515 6.665 -227.165 6.670 ;
        RECT -220.455 7.570 -219.105 7.575 ;
        RECT -218.595 7.570 -217.245 7.575 ;
        RECT -220.455 6.670 -217.245 7.570 ;
        RECT -220.455 6.665 -219.105 6.670 ;
        RECT -218.595 6.665 -217.245 6.670 ;
        RECT -210.535 7.570 -209.185 7.575 ;
        RECT -208.675 7.570 -207.325 7.575 ;
        RECT -210.535 6.670 -207.325 7.570 ;
        RECT -210.535 6.665 -209.185 6.670 ;
        RECT -208.675 6.665 -207.325 6.670 ;
        RECT -200.615 7.570 -199.265 7.575 ;
        RECT -198.755 7.570 -197.405 7.575 ;
        RECT -200.615 6.670 -197.405 7.570 ;
        RECT -200.615 6.665 -199.265 6.670 ;
        RECT -198.755 6.665 -197.405 6.670 ;
        RECT -190.695 7.570 -189.345 7.575 ;
        RECT -188.835 7.570 -187.485 7.575 ;
        RECT -190.695 6.670 -187.485 7.570 ;
        RECT -190.695 6.665 -189.345 6.670 ;
        RECT -188.835 6.665 -187.485 6.670 ;
        RECT -180.775 7.570 -179.425 7.575 ;
        RECT -178.915 7.570 -177.565 7.575 ;
        RECT -180.775 6.670 -177.565 7.570 ;
        RECT -180.775 6.665 -179.425 6.670 ;
        RECT -178.915 6.665 -177.565 6.670 ;
        RECT -170.855 7.570 -169.505 7.575 ;
        RECT -168.995 7.570 -167.645 7.575 ;
        RECT -170.855 6.670 -167.645 7.570 ;
        RECT -170.855 6.665 -169.505 6.670 ;
        RECT -168.995 6.665 -167.645 6.670 ;
        RECT -160.935 7.570 -159.585 7.575 ;
        RECT -159.075 7.570 -157.725 7.575 ;
        RECT -160.935 6.670 -157.725 7.570 ;
        RECT -160.935 6.665 -159.585 6.670 ;
        RECT -159.075 6.665 -157.725 6.670 ;
        RECT -151.015 7.570 -149.665 7.575 ;
        RECT -149.155 7.570 -147.805 7.575 ;
        RECT -151.015 6.670 -147.805 7.570 ;
        RECT -151.015 6.665 -149.665 6.670 ;
        RECT -149.155 6.665 -147.805 6.670 ;
        RECT -141.095 7.570 -139.745 7.575 ;
        RECT -139.235 7.570 -137.885 7.575 ;
        RECT -141.095 6.670 -137.885 7.570 ;
        RECT -141.095 6.665 -139.745 6.670 ;
        RECT -139.235 6.665 -137.885 6.670 ;
        RECT -131.175 7.570 -129.825 7.575 ;
        RECT -129.315 7.570 -127.965 7.575 ;
        RECT -131.175 6.670 -127.965 7.570 ;
        RECT -131.175 6.665 -129.825 6.670 ;
        RECT -129.315 6.665 -127.965 6.670 ;
        RECT -121.255 7.570 -119.905 7.575 ;
        RECT -119.395 7.570 -118.045 7.575 ;
        RECT -121.255 6.670 -118.045 7.570 ;
        RECT -121.255 6.665 -119.905 6.670 ;
        RECT -119.395 6.665 -118.045 6.670 ;
        RECT -111.335 7.570 -109.985 7.575 ;
        RECT -109.475 7.570 -108.125 7.575 ;
        RECT -111.335 6.670 -108.125 7.570 ;
        RECT -111.335 6.665 -109.985 6.670 ;
        RECT -109.475 6.665 -108.125 6.670 ;
        RECT -101.415 7.570 -100.065 7.575 ;
        RECT -99.555 7.570 -98.205 7.575 ;
        RECT -101.415 6.670 -98.205 7.570 ;
        RECT -101.415 6.665 -100.065 6.670 ;
        RECT -99.555 6.665 -98.205 6.670 ;
        RECT -91.495 7.570 -90.145 7.575 ;
        RECT -89.635 7.570 -88.285 7.575 ;
        RECT -91.495 6.670 -88.285 7.570 ;
        RECT -91.495 6.665 -90.145 6.670 ;
        RECT -89.635 6.665 -88.285 6.670 ;
        RECT -81.575 7.570 -80.225 7.575 ;
        RECT -79.715 7.570 -78.365 7.575 ;
        RECT -81.575 6.670 -78.365 7.570 ;
        RECT -81.575 6.665 -80.225 6.670 ;
        RECT -79.715 6.665 -78.365 6.670 ;
        RECT -71.655 7.570 -70.305 7.575 ;
        RECT -69.795 7.570 -68.445 7.575 ;
        RECT -71.655 6.670 -68.445 7.570 ;
        RECT -71.655 6.665 -70.305 6.670 ;
        RECT -69.795 6.665 -68.445 6.670 ;
        RECT -61.735 7.570 -60.385 7.575 ;
        RECT -59.875 7.570 -58.525 7.575 ;
        RECT -61.735 6.670 -58.525 7.570 ;
        RECT -61.735 6.665 -60.385 6.670 ;
        RECT -59.875 6.665 -58.525 6.670 ;
        RECT -51.815 7.570 -50.465 7.575 ;
        RECT -49.955 7.570 -48.605 7.575 ;
        RECT -51.815 6.670 -48.605 7.570 ;
        RECT -51.815 6.665 -50.465 6.670 ;
        RECT -49.955 6.665 -48.605 6.670 ;
        RECT -41.895 7.570 -40.545 7.575 ;
        RECT -40.035 7.570 -38.685 7.575 ;
        RECT -41.895 6.670 -38.685 7.570 ;
        RECT -41.895 6.665 -40.545 6.670 ;
        RECT -40.035 6.665 -38.685 6.670 ;
        RECT -31.975 7.570 -30.625 7.575 ;
        RECT -30.115 7.570 -28.765 7.575 ;
        RECT -31.975 6.670 -28.765 7.570 ;
        RECT -31.975 6.665 -30.625 6.670 ;
        RECT -30.115 6.665 -28.765 6.670 ;
        RECT -22.055 7.570 -20.705 7.575 ;
        RECT -20.195 7.570 -18.845 7.575 ;
        RECT -22.055 6.670 -18.845 7.570 ;
        RECT -22.055 6.665 -20.705 6.670 ;
        RECT -20.195 6.665 -18.845 6.670 ;
        RECT -12.135 7.570 -10.785 7.575 ;
        RECT -10.275 7.570 -8.925 7.575 ;
        RECT -12.135 6.670 -8.925 7.570 ;
        RECT -12.135 6.665 -10.785 6.670 ;
        RECT -10.275 6.665 -8.925 6.670 ;
        RECT -2.215 7.570 -0.865 7.575 ;
        RECT -0.355 7.570 0.995 7.575 ;
        RECT -2.215 6.670 0.995 7.570 ;
        RECT -2.215 6.665 -0.865 6.670 ;
        RECT -0.355 6.665 0.995 6.670 ;
        RECT 7.705 7.570 9.055 7.575 ;
        RECT 9.565 7.570 10.915 7.575 ;
        RECT 7.705 6.670 10.915 7.570 ;
        RECT 7.705 6.665 9.055 6.670 ;
        RECT 9.565 6.665 10.915 6.670 ;
        RECT 17.625 7.570 18.975 7.575 ;
        RECT 19.485 7.570 20.835 7.575 ;
        RECT 17.625 6.670 20.835 7.570 ;
        RECT 17.625 6.665 18.975 6.670 ;
        RECT 19.485 6.665 20.835 6.670 ;
        RECT -288.830 6.475 -288.660 6.665 ;
        RECT -287.920 6.475 -287.750 6.665 ;
        RECT -278.910 6.475 -278.740 6.665 ;
        RECT -278.000 6.475 -277.830 6.665 ;
        RECT -268.990 6.475 -268.820 6.665 ;
        RECT -268.080 6.475 -267.910 6.665 ;
        RECT -259.070 6.475 -258.900 6.665 ;
        RECT -258.160 6.475 -257.990 6.665 ;
        RECT -249.150 6.475 -248.980 6.665 ;
        RECT -248.240 6.475 -248.070 6.665 ;
        RECT -239.230 6.475 -239.060 6.665 ;
        RECT -238.320 6.475 -238.150 6.665 ;
        RECT -229.310 6.475 -229.140 6.665 ;
        RECT -228.400 6.475 -228.230 6.665 ;
        RECT -219.390 6.475 -219.220 6.665 ;
        RECT -218.480 6.475 -218.310 6.665 ;
        RECT -209.470 6.475 -209.300 6.665 ;
        RECT -208.560 6.475 -208.390 6.665 ;
        RECT -199.550 6.475 -199.380 6.665 ;
        RECT -198.640 6.475 -198.470 6.665 ;
        RECT -189.630 6.475 -189.460 6.665 ;
        RECT -188.720 6.475 -188.550 6.665 ;
        RECT -179.710 6.475 -179.540 6.665 ;
        RECT -178.800 6.475 -178.630 6.665 ;
        RECT -169.790 6.475 -169.620 6.665 ;
        RECT -168.880 6.475 -168.710 6.665 ;
        RECT -159.870 6.475 -159.700 6.665 ;
        RECT -158.960 6.475 -158.790 6.665 ;
        RECT -149.950 6.475 -149.780 6.665 ;
        RECT -149.040 6.475 -148.870 6.665 ;
        RECT -140.030 6.475 -139.860 6.665 ;
        RECT -139.120 6.475 -138.950 6.665 ;
        RECT -130.110 6.475 -129.940 6.665 ;
        RECT -129.200 6.475 -129.030 6.665 ;
        RECT -120.190 6.475 -120.020 6.665 ;
        RECT -119.280 6.475 -119.110 6.665 ;
        RECT -110.270 6.475 -110.100 6.665 ;
        RECT -109.360 6.475 -109.190 6.665 ;
        RECT -100.350 6.475 -100.180 6.665 ;
        RECT -99.440 6.475 -99.270 6.665 ;
        RECT -90.430 6.475 -90.260 6.665 ;
        RECT -89.520 6.475 -89.350 6.665 ;
        RECT -80.510 6.475 -80.340 6.665 ;
        RECT -79.600 6.475 -79.430 6.665 ;
        RECT -70.590 6.475 -70.420 6.665 ;
        RECT -69.680 6.475 -69.510 6.665 ;
        RECT -60.670 6.475 -60.500 6.665 ;
        RECT -59.760 6.475 -59.590 6.665 ;
        RECT -50.750 6.475 -50.580 6.665 ;
        RECT -49.840 6.475 -49.670 6.665 ;
        RECT -40.830 6.475 -40.660 6.665 ;
        RECT -39.920 6.475 -39.750 6.665 ;
        RECT -30.910 6.475 -30.740 6.665 ;
        RECT -30.000 6.475 -29.830 6.665 ;
        RECT -20.990 6.475 -20.820 6.665 ;
        RECT -20.080 6.475 -19.910 6.665 ;
        RECT -11.070 6.475 -10.900 6.665 ;
        RECT -10.160 6.475 -9.990 6.665 ;
        RECT -1.150 6.475 -0.980 6.665 ;
        RECT -0.240 6.475 -0.070 6.665 ;
        RECT 8.770 6.475 8.940 6.665 ;
        RECT 9.680 6.475 9.850 6.665 ;
        RECT 18.690 6.475 18.860 6.665 ;
        RECT 19.600 6.475 19.770 6.665 ;
        RECT -283.545 6.130 -283.115 6.145 ;
        RECT -273.625 6.130 -273.195 6.145 ;
        RECT -263.705 6.130 -263.275 6.145 ;
        RECT -253.785 6.130 -253.355 6.145 ;
        RECT -243.865 6.130 -243.435 6.145 ;
        RECT -233.945 6.130 -233.515 6.145 ;
        RECT -224.025 6.130 -223.595 6.145 ;
        RECT -214.105 6.130 -213.675 6.145 ;
        RECT -204.185 6.130 -203.755 6.145 ;
        RECT -194.265 6.130 -193.835 6.145 ;
        RECT -184.345 6.130 -183.915 6.145 ;
        RECT -174.425 6.130 -173.995 6.145 ;
        RECT -164.505 6.130 -164.075 6.145 ;
        RECT -154.585 6.130 -154.155 6.145 ;
        RECT -144.665 6.130 -144.235 6.145 ;
        RECT -134.745 6.130 -134.315 6.145 ;
        RECT -124.825 6.130 -124.395 6.145 ;
        RECT -114.905 6.130 -114.475 6.145 ;
        RECT -104.985 6.130 -104.555 6.145 ;
        RECT -95.065 6.130 -94.635 6.145 ;
        RECT -85.145 6.130 -84.715 6.145 ;
        RECT -75.225 6.130 -74.795 6.145 ;
        RECT -65.305 6.130 -64.875 6.145 ;
        RECT -55.385 6.130 -54.955 6.145 ;
        RECT -45.465 6.130 -45.035 6.145 ;
        RECT -35.545 6.130 -35.115 6.145 ;
        RECT -25.625 6.130 -25.195 6.145 ;
        RECT -15.705 6.130 -15.275 6.145 ;
        RECT -5.785 6.130 -5.355 6.145 ;
        RECT 4.135 6.130 4.565 6.145 ;
        RECT 14.055 6.130 14.485 6.145 ;
        RECT -285.380 6.125 -281.440 6.130 ;
        RECT -275.420 6.125 -271.400 6.130 ;
        RECT -265.540 6.125 -261.600 6.130 ;
        RECT -285.985 4.770 -280.675 6.125 ;
        RECT -285.985 4.755 -285.205 4.770 ;
        RECT -281.455 4.755 -280.675 4.770 ;
        RECT -276.065 4.755 -270.755 6.125 ;
        RECT -266.145 4.770 -260.835 6.125 ;
        RECT -266.145 4.755 -265.365 4.770 ;
        RECT -261.615 4.755 -260.835 4.770 ;
        RECT -256.225 6.120 -255.445 6.125 ;
        RECT -255.380 6.120 -251.930 6.130 ;
        RECT -245.700 6.125 -241.760 6.130 ;
        RECT -235.740 6.125 -231.720 6.130 ;
        RECT -225.860 6.125 -221.920 6.130 ;
        RECT -215.860 6.125 -211.790 6.130 ;
        RECT -206.020 6.125 -202.080 6.130 ;
        RECT -196.060 6.125 -192.040 6.130 ;
        RECT -186.180 6.125 -182.240 6.130 ;
        RECT -251.695 6.120 -250.915 6.125 ;
        RECT -256.225 4.755 -250.915 6.120 ;
        RECT -246.305 4.770 -240.995 6.125 ;
        RECT -246.305 4.755 -245.525 4.770 ;
        RECT -241.775 4.755 -240.995 4.770 ;
        RECT -236.385 4.755 -231.075 6.125 ;
        RECT -226.465 4.770 -221.155 6.125 ;
        RECT -226.465 4.755 -225.685 4.770 ;
        RECT -221.935 4.755 -221.155 4.770 ;
        RECT -216.545 4.760 -211.235 6.125 ;
        RECT -216.545 4.755 -215.765 4.760 ;
        RECT -212.015 4.755 -211.235 4.760 ;
        RECT -206.625 4.770 -201.315 6.125 ;
        RECT -206.625 4.755 -205.845 4.770 ;
        RECT -202.095 4.755 -201.315 4.770 ;
        RECT -196.705 4.755 -191.395 6.125 ;
        RECT -186.785 4.770 -181.475 6.125 ;
        RECT -186.785 4.755 -186.005 4.770 ;
        RECT -182.255 4.755 -181.475 4.770 ;
        RECT -176.865 6.120 -176.085 6.125 ;
        RECT -176.020 6.120 -172.570 6.130 ;
        RECT -166.340 6.125 -162.400 6.130 ;
        RECT -156.380 6.125 -152.360 6.130 ;
        RECT -146.500 6.125 -142.560 6.130 ;
        RECT -136.460 6.125 -132.520 6.130 ;
        RECT -126.660 6.125 -122.720 6.130 ;
        RECT -116.700 6.125 -112.680 6.130 ;
        RECT -106.820 6.125 -102.880 6.130 ;
        RECT -172.335 6.120 -171.555 6.125 ;
        RECT -176.865 4.755 -171.555 6.120 ;
        RECT -166.945 4.770 -161.635 6.125 ;
        RECT -166.945 4.755 -166.165 4.770 ;
        RECT -162.415 4.755 -161.635 4.770 ;
        RECT -157.025 4.755 -151.715 6.125 ;
        RECT -147.105 4.770 -141.795 6.125 ;
        RECT -147.105 4.755 -146.325 4.770 ;
        RECT -142.575 4.755 -141.795 4.770 ;
        RECT -137.185 4.770 -131.875 6.125 ;
        RECT -137.185 4.755 -136.405 4.770 ;
        RECT -132.655 4.755 -131.875 4.770 ;
        RECT -127.265 4.770 -121.955 6.125 ;
        RECT -127.265 4.755 -126.485 4.770 ;
        RECT -122.735 4.755 -121.955 4.770 ;
        RECT -117.345 4.755 -112.035 6.125 ;
        RECT -107.425 4.770 -102.115 6.125 ;
        RECT -107.425 4.755 -106.645 4.770 ;
        RECT -102.895 4.755 -102.115 4.770 ;
        RECT -97.505 6.120 -96.725 6.125 ;
        RECT -96.660 6.120 -93.210 6.130 ;
        RECT -86.980 6.125 -83.040 6.130 ;
        RECT -77.020 6.125 -73.000 6.130 ;
        RECT -67.140 6.125 -63.200 6.130 ;
        RECT -57.140 6.125 -53.070 6.130 ;
        RECT -47.300 6.125 -43.360 6.130 ;
        RECT -37.340 6.125 -33.320 6.130 ;
        RECT -27.460 6.125 -23.520 6.130 ;
        RECT -92.975 6.120 -92.195 6.125 ;
        RECT -97.505 4.755 -92.195 6.120 ;
        RECT -87.585 4.770 -82.275 6.125 ;
        RECT -87.585 4.755 -86.805 4.770 ;
        RECT -83.055 4.755 -82.275 4.770 ;
        RECT -77.665 4.755 -72.355 6.125 ;
        RECT -67.745 4.770 -62.435 6.125 ;
        RECT -67.745 4.755 -66.965 4.770 ;
        RECT -63.215 4.755 -62.435 4.770 ;
        RECT -57.825 4.760 -52.515 6.125 ;
        RECT -57.825 4.755 -57.045 4.760 ;
        RECT -53.295 4.755 -52.515 4.760 ;
        RECT -47.905 4.770 -42.595 6.125 ;
        RECT -47.905 4.755 -47.125 4.770 ;
        RECT -43.375 4.755 -42.595 4.770 ;
        RECT -37.985 4.755 -32.675 6.125 ;
        RECT -28.065 4.770 -22.755 6.125 ;
        RECT -28.065 4.755 -27.285 4.770 ;
        RECT -23.535 4.755 -22.755 4.770 ;
        RECT -18.145 6.120 -17.365 6.125 ;
        RECT -17.300 6.120 -13.850 6.130 ;
        RECT -7.620 6.125 -3.680 6.130 ;
        RECT 2.340 6.125 6.360 6.130 ;
        RECT 12.220 6.125 16.160 6.130 ;
        RECT -13.615 6.120 -12.835 6.125 ;
        RECT -18.145 4.755 -12.835 6.120 ;
        RECT -8.225 4.770 -2.915 6.125 ;
        RECT -8.225 4.755 -7.445 4.770 ;
        RECT -3.695 4.755 -2.915 4.770 ;
        RECT 1.695 4.755 7.005 6.125 ;
        RECT 11.615 4.770 16.925 6.125 ;
        RECT 11.615 4.755 12.395 4.770 ;
        RECT 16.145 4.755 16.925 4.770 ;
        RECT -275.420 4.750 -271.400 4.755 ;
        RECT -255.500 4.750 -251.660 4.755 ;
        RECT -235.740 4.750 -231.720 4.755 ;
        RECT -196.060 4.750 -192.040 4.755 ;
        RECT -176.140 4.750 -172.300 4.755 ;
        RECT -156.380 4.750 -152.360 4.755 ;
        RECT -116.700 4.750 -112.680 4.755 ;
        RECT -96.780 4.750 -92.940 4.755 ;
        RECT -77.020 4.750 -73.000 4.755 ;
        RECT -37.340 4.750 -33.320 4.755 ;
        RECT -17.420 4.750 -13.580 4.755 ;
        RECT 2.340 4.750 6.360 4.755 ;
        RECT -289.880 -77.865 -285.920 -77.860 ;
        RECT -279.960 -77.865 -276.000 -77.860 ;
        RECT -270.040 -77.865 -266.080 -77.860 ;
        RECT -260.120 -77.865 -256.160 -77.860 ;
        RECT -250.200 -77.865 -246.240 -77.860 ;
        RECT -240.280 -77.865 -236.320 -77.860 ;
        RECT -230.360 -77.865 -226.400 -77.860 ;
        RECT -220.440 -77.865 -216.480 -77.860 ;
        RECT -210.520 -77.865 -206.560 -77.860 ;
        RECT -200.600 -77.865 -196.640 -77.860 ;
        RECT -190.680 -77.865 -186.720 -77.860 ;
        RECT -180.760 -77.865 -176.800 -77.860 ;
        RECT -170.840 -77.865 -166.880 -77.860 ;
        RECT -160.920 -77.865 -156.960 -77.860 ;
        RECT -151.000 -77.865 -147.040 -77.860 ;
        RECT -141.080 -77.865 -137.120 -77.860 ;
        RECT -131.160 -77.865 -127.200 -77.860 ;
        RECT -121.240 -77.865 -117.280 -77.860 ;
        RECT -111.320 -77.865 -107.360 -77.860 ;
        RECT -101.400 -77.865 -97.440 -77.860 ;
        RECT -91.480 -77.865 -87.520 -77.860 ;
        RECT -81.560 -77.865 -77.600 -77.860 ;
        RECT -71.640 -77.865 -67.680 -77.860 ;
        RECT -61.720 -77.865 -57.760 -77.860 ;
        RECT -51.800 -77.865 -47.840 -77.860 ;
        RECT -41.880 -77.865 -37.920 -77.860 ;
        RECT -31.960 -77.865 -28.000 -77.860 ;
        RECT -22.040 -77.865 -18.080 -77.860 ;
        RECT -12.120 -77.865 -8.160 -77.860 ;
        RECT -2.200 -77.865 1.760 -77.860 ;
        RECT 7.720 -77.865 11.680 -77.860 ;
        RECT 17.640 -77.865 21.600 -77.860 ;
        RECT -290.585 -79.235 -285.275 -77.865 ;
        RECT -280.665 -79.235 -275.355 -77.865 ;
        RECT -270.745 -79.235 -265.435 -77.865 ;
        RECT -260.825 -79.235 -255.515 -77.865 ;
        RECT -250.905 -79.235 -245.595 -77.865 ;
        RECT -240.985 -79.235 -235.675 -77.865 ;
        RECT -231.065 -79.235 -225.755 -77.865 ;
        RECT -221.145 -79.235 -215.835 -77.865 ;
        RECT -211.225 -79.235 -205.915 -77.865 ;
        RECT -201.305 -79.235 -195.995 -77.865 ;
        RECT -191.385 -79.235 -186.075 -77.865 ;
        RECT -181.465 -79.235 -176.155 -77.865 ;
        RECT -171.545 -79.235 -166.235 -77.865 ;
        RECT -161.625 -79.235 -156.315 -77.865 ;
        RECT -151.705 -79.235 -146.395 -77.865 ;
        RECT -141.785 -79.235 -136.475 -77.865 ;
        RECT -131.865 -79.235 -126.555 -77.865 ;
        RECT -121.945 -79.235 -116.635 -77.865 ;
        RECT -112.025 -79.235 -106.715 -77.865 ;
        RECT -102.105 -79.235 -96.795 -77.865 ;
        RECT -92.185 -79.235 -86.875 -77.865 ;
        RECT -82.265 -79.235 -76.955 -77.865 ;
        RECT -72.345 -79.235 -67.035 -77.865 ;
        RECT -62.425 -79.235 -57.115 -77.865 ;
        RECT -52.505 -79.235 -47.195 -77.865 ;
        RECT -42.585 -79.235 -37.275 -77.865 ;
        RECT -32.665 -79.235 -27.355 -77.865 ;
        RECT -22.745 -79.235 -17.435 -77.865 ;
        RECT -12.825 -79.235 -7.515 -77.865 ;
        RECT -2.905 -79.235 2.405 -77.865 ;
        RECT 7.015 -79.235 12.325 -77.865 ;
        RECT 16.935 -79.235 22.245 -77.865 ;
        RECT -289.880 -79.240 -285.920 -79.235 ;
        RECT -279.960 -79.240 -276.000 -79.235 ;
        RECT -270.040 -79.240 -266.080 -79.235 ;
        RECT -260.120 -79.240 -256.160 -79.235 ;
        RECT -250.200 -79.240 -246.240 -79.235 ;
        RECT -240.280 -79.240 -236.320 -79.235 ;
        RECT -230.360 -79.240 -226.400 -79.235 ;
        RECT -220.440 -79.240 -216.480 -79.235 ;
        RECT -210.520 -79.240 -206.560 -79.235 ;
        RECT -200.600 -79.240 -196.640 -79.235 ;
        RECT -190.680 -79.240 -186.720 -79.235 ;
        RECT -180.760 -79.240 -176.800 -79.235 ;
        RECT -170.840 -79.240 -166.880 -79.235 ;
        RECT -160.920 -79.240 -156.960 -79.235 ;
        RECT -151.000 -79.240 -147.040 -79.235 ;
        RECT -141.080 -79.240 -137.120 -79.235 ;
        RECT -131.160 -79.240 -127.200 -79.235 ;
        RECT -121.240 -79.240 -117.280 -79.235 ;
        RECT -111.320 -79.240 -107.360 -79.235 ;
        RECT -101.400 -79.240 -97.440 -79.235 ;
        RECT -91.480 -79.240 -87.520 -79.235 ;
        RECT -81.560 -79.240 -77.600 -79.235 ;
        RECT -71.640 -79.240 -67.680 -79.235 ;
        RECT -61.720 -79.240 -57.760 -79.235 ;
        RECT -51.800 -79.240 -47.840 -79.235 ;
        RECT -41.880 -79.240 -37.920 -79.235 ;
        RECT -31.960 -79.240 -28.000 -79.235 ;
        RECT -22.040 -79.240 -18.080 -79.235 ;
        RECT -12.120 -79.240 -8.160 -79.235 ;
        RECT -2.200 -79.240 1.760 -79.235 ;
        RECT 7.720 -79.240 11.680 -79.235 ;
        RECT 17.640 -79.240 21.600 -79.235 ;
        RECT -283.510 -79.775 -283.340 -79.585 ;
        RECT -282.600 -79.775 -282.430 -79.585 ;
        RECT -273.590 -79.775 -273.420 -79.585 ;
        RECT -272.680 -79.775 -272.510 -79.585 ;
        RECT -263.670 -79.775 -263.500 -79.585 ;
        RECT -262.760 -79.775 -262.590 -79.585 ;
        RECT -253.750 -79.775 -253.580 -79.585 ;
        RECT -252.840 -79.775 -252.670 -79.585 ;
        RECT -243.830 -79.775 -243.660 -79.585 ;
        RECT -242.920 -79.775 -242.750 -79.585 ;
        RECT -233.910 -79.775 -233.740 -79.585 ;
        RECT -233.000 -79.775 -232.830 -79.585 ;
        RECT -223.990 -79.775 -223.820 -79.585 ;
        RECT -223.080 -79.775 -222.910 -79.585 ;
        RECT -214.070 -79.775 -213.900 -79.585 ;
        RECT -213.160 -79.775 -212.990 -79.585 ;
        RECT -204.150 -79.775 -203.980 -79.585 ;
        RECT -203.240 -79.775 -203.070 -79.585 ;
        RECT -194.230 -79.775 -194.060 -79.585 ;
        RECT -193.320 -79.775 -193.150 -79.585 ;
        RECT -184.310 -79.775 -184.140 -79.585 ;
        RECT -183.400 -79.775 -183.230 -79.585 ;
        RECT -174.390 -79.775 -174.220 -79.585 ;
        RECT -173.480 -79.775 -173.310 -79.585 ;
        RECT -164.470 -79.775 -164.300 -79.585 ;
        RECT -163.560 -79.775 -163.390 -79.585 ;
        RECT -154.550 -79.775 -154.380 -79.585 ;
        RECT -153.640 -79.775 -153.470 -79.585 ;
        RECT -144.630 -79.775 -144.460 -79.585 ;
        RECT -143.720 -79.775 -143.550 -79.585 ;
        RECT -134.710 -79.775 -134.540 -79.585 ;
        RECT -133.800 -79.775 -133.630 -79.585 ;
        RECT -124.790 -79.775 -124.620 -79.585 ;
        RECT -123.880 -79.775 -123.710 -79.585 ;
        RECT -114.870 -79.775 -114.700 -79.585 ;
        RECT -113.960 -79.775 -113.790 -79.585 ;
        RECT -104.950 -79.775 -104.780 -79.585 ;
        RECT -104.040 -79.775 -103.870 -79.585 ;
        RECT -95.030 -79.775 -94.860 -79.585 ;
        RECT -94.120 -79.775 -93.950 -79.585 ;
        RECT -85.110 -79.775 -84.940 -79.585 ;
        RECT -84.200 -79.775 -84.030 -79.585 ;
        RECT -75.190 -79.775 -75.020 -79.585 ;
        RECT -74.280 -79.775 -74.110 -79.585 ;
        RECT -65.270 -79.775 -65.100 -79.585 ;
        RECT -64.360 -79.775 -64.190 -79.585 ;
        RECT -55.350 -79.775 -55.180 -79.585 ;
        RECT -54.440 -79.775 -54.270 -79.585 ;
        RECT -45.430 -79.775 -45.260 -79.585 ;
        RECT -44.520 -79.775 -44.350 -79.585 ;
        RECT -35.510 -79.775 -35.340 -79.585 ;
        RECT -34.600 -79.775 -34.430 -79.585 ;
        RECT -25.590 -79.775 -25.420 -79.585 ;
        RECT -24.680 -79.775 -24.510 -79.585 ;
        RECT -15.670 -79.775 -15.500 -79.585 ;
        RECT -14.760 -79.775 -14.590 -79.585 ;
        RECT -5.750 -79.775 -5.580 -79.585 ;
        RECT -4.840 -79.775 -4.670 -79.585 ;
        RECT 4.170 -79.775 4.340 -79.585 ;
        RECT 5.080 -79.775 5.250 -79.585 ;
        RECT 14.090 -79.775 14.260 -79.585 ;
        RECT 15.000 -79.775 15.170 -79.585 ;
        RECT -284.575 -79.780 -283.225 -79.775 ;
        RECT -282.715 -79.780 -281.365 -79.775 ;
        RECT -284.575 -80.680 -281.365 -79.780 ;
        RECT -284.575 -80.685 -283.225 -80.680 ;
        RECT -282.715 -80.685 -281.365 -80.680 ;
        RECT -274.655 -79.780 -273.305 -79.775 ;
        RECT -272.795 -79.780 -271.445 -79.775 ;
        RECT -274.655 -80.680 -271.445 -79.780 ;
        RECT -274.655 -80.685 -273.305 -80.680 ;
        RECT -272.795 -80.685 -271.445 -80.680 ;
        RECT -264.735 -79.780 -263.385 -79.775 ;
        RECT -262.875 -79.780 -261.525 -79.775 ;
        RECT -264.735 -80.680 -261.525 -79.780 ;
        RECT -264.735 -80.685 -263.385 -80.680 ;
        RECT -262.875 -80.685 -261.525 -80.680 ;
        RECT -254.815 -79.780 -253.465 -79.775 ;
        RECT -252.955 -79.780 -251.605 -79.775 ;
        RECT -254.815 -80.680 -251.605 -79.780 ;
        RECT -254.815 -80.685 -253.465 -80.680 ;
        RECT -252.955 -80.685 -251.605 -80.680 ;
        RECT -244.895 -79.780 -243.545 -79.775 ;
        RECT -243.035 -79.780 -241.685 -79.775 ;
        RECT -244.895 -80.680 -241.685 -79.780 ;
        RECT -244.895 -80.685 -243.545 -80.680 ;
        RECT -243.035 -80.685 -241.685 -80.680 ;
        RECT -234.975 -79.780 -233.625 -79.775 ;
        RECT -233.115 -79.780 -231.765 -79.775 ;
        RECT -234.975 -80.680 -231.765 -79.780 ;
        RECT -234.975 -80.685 -233.625 -80.680 ;
        RECT -233.115 -80.685 -231.765 -80.680 ;
        RECT -225.055 -79.780 -223.705 -79.775 ;
        RECT -223.195 -79.780 -221.845 -79.775 ;
        RECT -225.055 -80.680 -221.845 -79.780 ;
        RECT -225.055 -80.685 -223.705 -80.680 ;
        RECT -223.195 -80.685 -221.845 -80.680 ;
        RECT -215.135 -79.780 -213.785 -79.775 ;
        RECT -213.275 -79.780 -211.925 -79.775 ;
        RECT -215.135 -80.680 -211.925 -79.780 ;
        RECT -215.135 -80.685 -213.785 -80.680 ;
        RECT -213.275 -80.685 -211.925 -80.680 ;
        RECT -205.215 -79.780 -203.865 -79.775 ;
        RECT -203.355 -79.780 -202.005 -79.775 ;
        RECT -205.215 -80.680 -202.005 -79.780 ;
        RECT -205.215 -80.685 -203.865 -80.680 ;
        RECT -203.355 -80.685 -202.005 -80.680 ;
        RECT -195.295 -79.780 -193.945 -79.775 ;
        RECT -193.435 -79.780 -192.085 -79.775 ;
        RECT -195.295 -80.680 -192.085 -79.780 ;
        RECT -195.295 -80.685 -193.945 -80.680 ;
        RECT -193.435 -80.685 -192.085 -80.680 ;
        RECT -185.375 -79.780 -184.025 -79.775 ;
        RECT -183.515 -79.780 -182.165 -79.775 ;
        RECT -185.375 -80.680 -182.165 -79.780 ;
        RECT -185.375 -80.685 -184.025 -80.680 ;
        RECT -183.515 -80.685 -182.165 -80.680 ;
        RECT -175.455 -79.780 -174.105 -79.775 ;
        RECT -173.595 -79.780 -172.245 -79.775 ;
        RECT -175.455 -80.680 -172.245 -79.780 ;
        RECT -175.455 -80.685 -174.105 -80.680 ;
        RECT -173.595 -80.685 -172.245 -80.680 ;
        RECT -165.535 -79.780 -164.185 -79.775 ;
        RECT -163.675 -79.780 -162.325 -79.775 ;
        RECT -165.535 -80.680 -162.325 -79.780 ;
        RECT -165.535 -80.685 -164.185 -80.680 ;
        RECT -163.675 -80.685 -162.325 -80.680 ;
        RECT -155.615 -79.780 -154.265 -79.775 ;
        RECT -153.755 -79.780 -152.405 -79.775 ;
        RECT -155.615 -80.680 -152.405 -79.780 ;
        RECT -155.615 -80.685 -154.265 -80.680 ;
        RECT -153.755 -80.685 -152.405 -80.680 ;
        RECT -145.695 -79.780 -144.345 -79.775 ;
        RECT -143.835 -79.780 -142.485 -79.775 ;
        RECT -145.695 -80.680 -142.485 -79.780 ;
        RECT -145.695 -80.685 -144.345 -80.680 ;
        RECT -143.835 -80.685 -142.485 -80.680 ;
        RECT -135.775 -79.780 -134.425 -79.775 ;
        RECT -133.915 -79.780 -132.565 -79.775 ;
        RECT -135.775 -80.680 -132.565 -79.780 ;
        RECT -135.775 -80.685 -134.425 -80.680 ;
        RECT -133.915 -80.685 -132.565 -80.680 ;
        RECT -125.855 -79.780 -124.505 -79.775 ;
        RECT -123.995 -79.780 -122.645 -79.775 ;
        RECT -125.855 -80.680 -122.645 -79.780 ;
        RECT -125.855 -80.685 -124.505 -80.680 ;
        RECT -123.995 -80.685 -122.645 -80.680 ;
        RECT -115.935 -79.780 -114.585 -79.775 ;
        RECT -114.075 -79.780 -112.725 -79.775 ;
        RECT -115.935 -80.680 -112.725 -79.780 ;
        RECT -115.935 -80.685 -114.585 -80.680 ;
        RECT -114.075 -80.685 -112.725 -80.680 ;
        RECT -106.015 -79.780 -104.665 -79.775 ;
        RECT -104.155 -79.780 -102.805 -79.775 ;
        RECT -106.015 -80.680 -102.805 -79.780 ;
        RECT -106.015 -80.685 -104.665 -80.680 ;
        RECT -104.155 -80.685 -102.805 -80.680 ;
        RECT -96.095 -79.780 -94.745 -79.775 ;
        RECT -94.235 -79.780 -92.885 -79.775 ;
        RECT -96.095 -80.680 -92.885 -79.780 ;
        RECT -96.095 -80.685 -94.745 -80.680 ;
        RECT -94.235 -80.685 -92.885 -80.680 ;
        RECT -86.175 -79.780 -84.825 -79.775 ;
        RECT -84.315 -79.780 -82.965 -79.775 ;
        RECT -86.175 -80.680 -82.965 -79.780 ;
        RECT -86.175 -80.685 -84.825 -80.680 ;
        RECT -84.315 -80.685 -82.965 -80.680 ;
        RECT -76.255 -79.780 -74.905 -79.775 ;
        RECT -74.395 -79.780 -73.045 -79.775 ;
        RECT -76.255 -80.680 -73.045 -79.780 ;
        RECT -76.255 -80.685 -74.905 -80.680 ;
        RECT -74.395 -80.685 -73.045 -80.680 ;
        RECT -66.335 -79.780 -64.985 -79.775 ;
        RECT -64.475 -79.780 -63.125 -79.775 ;
        RECT -66.335 -80.680 -63.125 -79.780 ;
        RECT -66.335 -80.685 -64.985 -80.680 ;
        RECT -64.475 -80.685 -63.125 -80.680 ;
        RECT -56.415 -79.780 -55.065 -79.775 ;
        RECT -54.555 -79.780 -53.205 -79.775 ;
        RECT -56.415 -80.680 -53.205 -79.780 ;
        RECT -56.415 -80.685 -55.065 -80.680 ;
        RECT -54.555 -80.685 -53.205 -80.680 ;
        RECT -46.495 -79.780 -45.145 -79.775 ;
        RECT -44.635 -79.780 -43.285 -79.775 ;
        RECT -46.495 -80.680 -43.285 -79.780 ;
        RECT -46.495 -80.685 -45.145 -80.680 ;
        RECT -44.635 -80.685 -43.285 -80.680 ;
        RECT -36.575 -79.780 -35.225 -79.775 ;
        RECT -34.715 -79.780 -33.365 -79.775 ;
        RECT -36.575 -80.680 -33.365 -79.780 ;
        RECT -36.575 -80.685 -35.225 -80.680 ;
        RECT -34.715 -80.685 -33.365 -80.680 ;
        RECT -26.655 -79.780 -25.305 -79.775 ;
        RECT -24.795 -79.780 -23.445 -79.775 ;
        RECT -26.655 -80.680 -23.445 -79.780 ;
        RECT -26.655 -80.685 -25.305 -80.680 ;
        RECT -24.795 -80.685 -23.445 -80.680 ;
        RECT -16.735 -79.780 -15.385 -79.775 ;
        RECT -14.875 -79.780 -13.525 -79.775 ;
        RECT -16.735 -80.680 -13.525 -79.780 ;
        RECT -16.735 -80.685 -15.385 -80.680 ;
        RECT -14.875 -80.685 -13.525 -80.680 ;
        RECT -6.815 -79.780 -5.465 -79.775 ;
        RECT -4.955 -79.780 -3.605 -79.775 ;
        RECT -6.815 -80.680 -3.605 -79.780 ;
        RECT -6.815 -80.685 -5.465 -80.680 ;
        RECT -4.955 -80.685 -3.605 -80.680 ;
        RECT 3.105 -79.780 4.455 -79.775 ;
        RECT 4.965 -79.780 6.315 -79.775 ;
        RECT 3.105 -80.680 6.315 -79.780 ;
        RECT 3.105 -80.685 4.455 -80.680 ;
        RECT 4.965 -80.685 6.315 -80.680 ;
        RECT 13.025 -79.780 14.375 -79.775 ;
        RECT 14.885 -79.780 16.235 -79.775 ;
        RECT 13.025 -80.680 16.235 -79.780 ;
        RECT 13.025 -80.685 14.375 -80.680 ;
        RECT 14.885 -80.685 16.235 -80.680 ;
        RECT -289.535 -81.380 -288.185 -81.375 ;
        RECT -287.675 -81.380 -286.325 -81.375 ;
        RECT -289.535 -82.280 -286.325 -81.380 ;
        RECT -289.535 -82.285 -288.185 -82.280 ;
        RECT -287.675 -82.285 -286.325 -82.280 ;
        RECT -279.615 -81.380 -278.265 -81.375 ;
        RECT -277.755 -81.380 -276.405 -81.375 ;
        RECT -279.615 -82.280 -276.405 -81.380 ;
        RECT -279.615 -82.285 -278.265 -82.280 ;
        RECT -277.755 -82.285 -276.405 -82.280 ;
        RECT -269.695 -81.380 -268.345 -81.375 ;
        RECT -267.835 -81.380 -266.485 -81.375 ;
        RECT -269.695 -82.280 -266.485 -81.380 ;
        RECT -269.695 -82.285 -268.345 -82.280 ;
        RECT -267.835 -82.285 -266.485 -82.280 ;
        RECT -259.775 -81.380 -258.425 -81.375 ;
        RECT -257.915 -81.380 -256.565 -81.375 ;
        RECT -259.775 -82.280 -256.565 -81.380 ;
        RECT -259.775 -82.285 -258.425 -82.280 ;
        RECT -257.915 -82.285 -256.565 -82.280 ;
        RECT -249.855 -81.380 -248.505 -81.375 ;
        RECT -247.995 -81.380 -246.645 -81.375 ;
        RECT -249.855 -82.280 -246.645 -81.380 ;
        RECT -249.855 -82.285 -248.505 -82.280 ;
        RECT -247.995 -82.285 -246.645 -82.280 ;
        RECT -239.935 -81.380 -238.585 -81.375 ;
        RECT -238.075 -81.380 -236.725 -81.375 ;
        RECT -239.935 -82.280 -236.725 -81.380 ;
        RECT -239.935 -82.285 -238.585 -82.280 ;
        RECT -238.075 -82.285 -236.725 -82.280 ;
        RECT -230.015 -81.380 -228.665 -81.375 ;
        RECT -228.155 -81.380 -226.805 -81.375 ;
        RECT -230.015 -82.280 -226.805 -81.380 ;
        RECT -230.015 -82.285 -228.665 -82.280 ;
        RECT -228.155 -82.285 -226.805 -82.280 ;
        RECT -220.095 -81.380 -218.745 -81.375 ;
        RECT -218.235 -81.380 -216.885 -81.375 ;
        RECT -220.095 -82.280 -216.885 -81.380 ;
        RECT -220.095 -82.285 -218.745 -82.280 ;
        RECT -218.235 -82.285 -216.885 -82.280 ;
        RECT -210.175 -81.380 -208.825 -81.375 ;
        RECT -208.315 -81.380 -206.965 -81.375 ;
        RECT -210.175 -82.280 -206.965 -81.380 ;
        RECT -210.175 -82.285 -208.825 -82.280 ;
        RECT -208.315 -82.285 -206.965 -82.280 ;
        RECT -200.255 -81.380 -198.905 -81.375 ;
        RECT -198.395 -81.380 -197.045 -81.375 ;
        RECT -200.255 -82.280 -197.045 -81.380 ;
        RECT -200.255 -82.285 -198.905 -82.280 ;
        RECT -198.395 -82.285 -197.045 -82.280 ;
        RECT -190.335 -81.380 -188.985 -81.375 ;
        RECT -188.475 -81.380 -187.125 -81.375 ;
        RECT -190.335 -82.280 -187.125 -81.380 ;
        RECT -190.335 -82.285 -188.985 -82.280 ;
        RECT -188.475 -82.285 -187.125 -82.280 ;
        RECT -180.415 -81.380 -179.065 -81.375 ;
        RECT -178.555 -81.380 -177.205 -81.375 ;
        RECT -180.415 -82.280 -177.205 -81.380 ;
        RECT -180.415 -82.285 -179.065 -82.280 ;
        RECT -178.555 -82.285 -177.205 -82.280 ;
        RECT -170.495 -81.380 -169.145 -81.375 ;
        RECT -168.635 -81.380 -167.285 -81.375 ;
        RECT -170.495 -82.280 -167.285 -81.380 ;
        RECT -170.495 -82.285 -169.145 -82.280 ;
        RECT -168.635 -82.285 -167.285 -82.280 ;
        RECT -160.575 -81.380 -159.225 -81.375 ;
        RECT -158.715 -81.380 -157.365 -81.375 ;
        RECT -160.575 -82.280 -157.365 -81.380 ;
        RECT -160.575 -82.285 -159.225 -82.280 ;
        RECT -158.715 -82.285 -157.365 -82.280 ;
        RECT -150.655 -81.380 -149.305 -81.375 ;
        RECT -148.795 -81.380 -147.445 -81.375 ;
        RECT -150.655 -82.280 -147.445 -81.380 ;
        RECT -150.655 -82.285 -149.305 -82.280 ;
        RECT -148.795 -82.285 -147.445 -82.280 ;
        RECT -140.735 -81.380 -139.385 -81.375 ;
        RECT -138.875 -81.380 -137.525 -81.375 ;
        RECT -140.735 -82.280 -137.525 -81.380 ;
        RECT -140.735 -82.285 -139.385 -82.280 ;
        RECT -138.875 -82.285 -137.525 -82.280 ;
        RECT -130.815 -81.380 -129.465 -81.375 ;
        RECT -128.955 -81.380 -127.605 -81.375 ;
        RECT -130.815 -82.280 -127.605 -81.380 ;
        RECT -130.815 -82.285 -129.465 -82.280 ;
        RECT -128.955 -82.285 -127.605 -82.280 ;
        RECT -120.895 -81.380 -119.545 -81.375 ;
        RECT -119.035 -81.380 -117.685 -81.375 ;
        RECT -120.895 -82.280 -117.685 -81.380 ;
        RECT -120.895 -82.285 -119.545 -82.280 ;
        RECT -119.035 -82.285 -117.685 -82.280 ;
        RECT -110.975 -81.380 -109.625 -81.375 ;
        RECT -109.115 -81.380 -107.765 -81.375 ;
        RECT -110.975 -82.280 -107.765 -81.380 ;
        RECT -110.975 -82.285 -109.625 -82.280 ;
        RECT -109.115 -82.285 -107.765 -82.280 ;
        RECT -101.055 -81.380 -99.705 -81.375 ;
        RECT -99.195 -81.380 -97.845 -81.375 ;
        RECT -101.055 -82.280 -97.845 -81.380 ;
        RECT -101.055 -82.285 -99.705 -82.280 ;
        RECT -99.195 -82.285 -97.845 -82.280 ;
        RECT -91.135 -81.380 -89.785 -81.375 ;
        RECT -89.275 -81.380 -87.925 -81.375 ;
        RECT -91.135 -82.280 -87.925 -81.380 ;
        RECT -91.135 -82.285 -89.785 -82.280 ;
        RECT -89.275 -82.285 -87.925 -82.280 ;
        RECT -81.215 -81.380 -79.865 -81.375 ;
        RECT -79.355 -81.380 -78.005 -81.375 ;
        RECT -81.215 -82.280 -78.005 -81.380 ;
        RECT -81.215 -82.285 -79.865 -82.280 ;
        RECT -79.355 -82.285 -78.005 -82.280 ;
        RECT -71.295 -81.380 -69.945 -81.375 ;
        RECT -69.435 -81.380 -68.085 -81.375 ;
        RECT -71.295 -82.280 -68.085 -81.380 ;
        RECT -71.295 -82.285 -69.945 -82.280 ;
        RECT -69.435 -82.285 -68.085 -82.280 ;
        RECT -61.375 -81.380 -60.025 -81.375 ;
        RECT -59.515 -81.380 -58.165 -81.375 ;
        RECT -61.375 -82.280 -58.165 -81.380 ;
        RECT -61.375 -82.285 -60.025 -82.280 ;
        RECT -59.515 -82.285 -58.165 -82.280 ;
        RECT -51.455 -81.380 -50.105 -81.375 ;
        RECT -49.595 -81.380 -48.245 -81.375 ;
        RECT -51.455 -82.280 -48.245 -81.380 ;
        RECT -51.455 -82.285 -50.105 -82.280 ;
        RECT -49.595 -82.285 -48.245 -82.280 ;
        RECT -41.535 -81.380 -40.185 -81.375 ;
        RECT -39.675 -81.380 -38.325 -81.375 ;
        RECT -41.535 -82.280 -38.325 -81.380 ;
        RECT -41.535 -82.285 -40.185 -82.280 ;
        RECT -39.675 -82.285 -38.325 -82.280 ;
        RECT -31.615 -81.380 -30.265 -81.375 ;
        RECT -29.755 -81.380 -28.405 -81.375 ;
        RECT -31.615 -82.280 -28.405 -81.380 ;
        RECT -31.615 -82.285 -30.265 -82.280 ;
        RECT -29.755 -82.285 -28.405 -82.280 ;
        RECT -21.695 -81.380 -20.345 -81.375 ;
        RECT -19.835 -81.380 -18.485 -81.375 ;
        RECT -21.695 -82.280 -18.485 -81.380 ;
        RECT -21.695 -82.285 -20.345 -82.280 ;
        RECT -19.835 -82.285 -18.485 -82.280 ;
        RECT -11.775 -81.380 -10.425 -81.375 ;
        RECT -9.915 -81.380 -8.565 -81.375 ;
        RECT -11.775 -82.280 -8.565 -81.380 ;
        RECT -11.775 -82.285 -10.425 -82.280 ;
        RECT -9.915 -82.285 -8.565 -82.280 ;
        RECT -1.855 -81.380 -0.505 -81.375 ;
        RECT 0.005 -81.380 1.355 -81.375 ;
        RECT -1.855 -82.280 1.355 -81.380 ;
        RECT -1.855 -82.285 -0.505 -82.280 ;
        RECT 0.005 -82.285 1.355 -82.280 ;
        RECT 8.065 -81.380 9.415 -81.375 ;
        RECT 9.925 -81.380 11.275 -81.375 ;
        RECT 8.065 -82.280 11.275 -81.380 ;
        RECT 8.065 -82.285 9.415 -82.280 ;
        RECT 9.925 -82.285 11.275 -82.280 ;
        RECT 17.985 -81.380 19.335 -81.375 ;
        RECT 19.845 -81.380 21.195 -81.375 ;
        RECT 17.985 -82.280 21.195 -81.380 ;
        RECT 17.985 -82.285 19.335 -82.280 ;
        RECT 19.845 -82.285 21.195 -82.280 ;
        RECT -288.470 -82.475 -288.300 -82.285 ;
        RECT -287.560 -82.475 -287.390 -82.285 ;
        RECT -278.550 -82.475 -278.380 -82.285 ;
        RECT -277.640 -82.475 -277.470 -82.285 ;
        RECT -268.630 -82.475 -268.460 -82.285 ;
        RECT -267.720 -82.475 -267.550 -82.285 ;
        RECT -258.710 -82.475 -258.540 -82.285 ;
        RECT -257.800 -82.475 -257.630 -82.285 ;
        RECT -248.790 -82.475 -248.620 -82.285 ;
        RECT -247.880 -82.475 -247.710 -82.285 ;
        RECT -238.870 -82.475 -238.700 -82.285 ;
        RECT -237.960 -82.475 -237.790 -82.285 ;
        RECT -228.950 -82.475 -228.780 -82.285 ;
        RECT -228.040 -82.475 -227.870 -82.285 ;
        RECT -219.030 -82.475 -218.860 -82.285 ;
        RECT -218.120 -82.475 -217.950 -82.285 ;
        RECT -209.110 -82.475 -208.940 -82.285 ;
        RECT -208.200 -82.475 -208.030 -82.285 ;
        RECT -199.190 -82.475 -199.020 -82.285 ;
        RECT -198.280 -82.475 -198.110 -82.285 ;
        RECT -189.270 -82.475 -189.100 -82.285 ;
        RECT -188.360 -82.475 -188.190 -82.285 ;
        RECT -179.350 -82.475 -179.180 -82.285 ;
        RECT -178.440 -82.475 -178.270 -82.285 ;
        RECT -169.430 -82.475 -169.260 -82.285 ;
        RECT -168.520 -82.475 -168.350 -82.285 ;
        RECT -159.510 -82.475 -159.340 -82.285 ;
        RECT -158.600 -82.475 -158.430 -82.285 ;
        RECT -149.590 -82.475 -149.420 -82.285 ;
        RECT -148.680 -82.475 -148.510 -82.285 ;
        RECT -139.670 -82.475 -139.500 -82.285 ;
        RECT -138.760 -82.475 -138.590 -82.285 ;
        RECT -129.750 -82.475 -129.580 -82.285 ;
        RECT -128.840 -82.475 -128.670 -82.285 ;
        RECT -119.830 -82.475 -119.660 -82.285 ;
        RECT -118.920 -82.475 -118.750 -82.285 ;
        RECT -109.910 -82.475 -109.740 -82.285 ;
        RECT -109.000 -82.475 -108.830 -82.285 ;
        RECT -99.990 -82.475 -99.820 -82.285 ;
        RECT -99.080 -82.475 -98.910 -82.285 ;
        RECT -90.070 -82.475 -89.900 -82.285 ;
        RECT -89.160 -82.475 -88.990 -82.285 ;
        RECT -80.150 -82.475 -79.980 -82.285 ;
        RECT -79.240 -82.475 -79.070 -82.285 ;
        RECT -70.230 -82.475 -70.060 -82.285 ;
        RECT -69.320 -82.475 -69.150 -82.285 ;
        RECT -60.310 -82.475 -60.140 -82.285 ;
        RECT -59.400 -82.475 -59.230 -82.285 ;
        RECT -50.390 -82.475 -50.220 -82.285 ;
        RECT -49.480 -82.475 -49.310 -82.285 ;
        RECT -40.470 -82.475 -40.300 -82.285 ;
        RECT -39.560 -82.475 -39.390 -82.285 ;
        RECT -30.550 -82.475 -30.380 -82.285 ;
        RECT -29.640 -82.475 -29.470 -82.285 ;
        RECT -20.630 -82.475 -20.460 -82.285 ;
        RECT -19.720 -82.475 -19.550 -82.285 ;
        RECT -10.710 -82.475 -10.540 -82.285 ;
        RECT -9.800 -82.475 -9.630 -82.285 ;
        RECT -0.790 -82.475 -0.620 -82.285 ;
        RECT 0.120 -82.475 0.290 -82.285 ;
        RECT 9.130 -82.475 9.300 -82.285 ;
        RECT 10.040 -82.475 10.210 -82.285 ;
        RECT 19.050 -82.475 19.220 -82.285 ;
        RECT 19.960 -82.475 20.130 -82.285 ;
        RECT -283.185 -82.820 -282.755 -82.805 ;
        RECT -273.265 -82.820 -272.835 -82.805 ;
        RECT -263.345 -82.820 -262.915 -82.805 ;
        RECT -253.425 -82.820 -252.995 -82.805 ;
        RECT -243.505 -82.820 -243.075 -82.805 ;
        RECT -233.585 -82.820 -233.155 -82.805 ;
        RECT -223.665 -82.820 -223.235 -82.805 ;
        RECT -213.745 -82.820 -213.315 -82.805 ;
        RECT -203.825 -82.820 -203.395 -82.805 ;
        RECT -193.905 -82.820 -193.475 -82.805 ;
        RECT -183.985 -82.820 -183.555 -82.805 ;
        RECT -174.065 -82.820 -173.635 -82.805 ;
        RECT -164.145 -82.820 -163.715 -82.805 ;
        RECT -154.225 -82.820 -153.795 -82.805 ;
        RECT -144.305 -82.820 -143.875 -82.805 ;
        RECT -134.385 -82.820 -133.955 -82.805 ;
        RECT -124.465 -82.820 -124.035 -82.805 ;
        RECT -114.545 -82.820 -114.115 -82.805 ;
        RECT -104.625 -82.820 -104.195 -82.805 ;
        RECT -94.705 -82.820 -94.275 -82.805 ;
        RECT -84.785 -82.820 -84.355 -82.805 ;
        RECT -74.865 -82.820 -74.435 -82.805 ;
        RECT -64.945 -82.820 -64.515 -82.805 ;
        RECT -55.025 -82.820 -54.595 -82.805 ;
        RECT -45.105 -82.820 -44.675 -82.805 ;
        RECT -35.185 -82.820 -34.755 -82.805 ;
        RECT -25.265 -82.820 -24.835 -82.805 ;
        RECT -15.345 -82.820 -14.915 -82.805 ;
        RECT -5.425 -82.820 -4.995 -82.805 ;
        RECT 4.495 -82.820 4.925 -82.805 ;
        RECT 14.415 -82.820 14.845 -82.805 ;
        RECT -285.020 -82.825 -281.080 -82.820 ;
        RECT -275.060 -82.825 -271.040 -82.820 ;
        RECT -265.180 -82.825 -261.240 -82.820 ;
        RECT -285.625 -84.180 -280.315 -82.825 ;
        RECT -285.625 -84.195 -284.845 -84.180 ;
        RECT -281.095 -84.195 -280.315 -84.180 ;
        RECT -275.705 -84.195 -270.395 -82.825 ;
        RECT -265.785 -84.180 -260.475 -82.825 ;
        RECT -265.785 -84.195 -265.005 -84.180 ;
        RECT -261.255 -84.195 -260.475 -84.180 ;
        RECT -255.865 -82.830 -255.085 -82.825 ;
        RECT -255.020 -82.830 -251.570 -82.820 ;
        RECT -245.340 -82.825 -241.400 -82.820 ;
        RECT -235.380 -82.825 -231.360 -82.820 ;
        RECT -225.500 -82.825 -221.560 -82.820 ;
        RECT -215.500 -82.825 -211.430 -82.820 ;
        RECT -205.660 -82.825 -201.720 -82.820 ;
        RECT -195.700 -82.825 -191.680 -82.820 ;
        RECT -185.820 -82.825 -181.880 -82.820 ;
        RECT -251.335 -82.830 -250.555 -82.825 ;
        RECT -255.865 -84.195 -250.555 -82.830 ;
        RECT -245.945 -84.180 -240.635 -82.825 ;
        RECT -245.945 -84.195 -245.165 -84.180 ;
        RECT -241.415 -84.195 -240.635 -84.180 ;
        RECT -236.025 -84.195 -230.715 -82.825 ;
        RECT -226.105 -84.180 -220.795 -82.825 ;
        RECT -226.105 -84.195 -225.325 -84.180 ;
        RECT -221.575 -84.195 -220.795 -84.180 ;
        RECT -216.185 -84.190 -210.875 -82.825 ;
        RECT -216.185 -84.195 -215.405 -84.190 ;
        RECT -211.655 -84.195 -210.875 -84.190 ;
        RECT -206.265 -84.180 -200.955 -82.825 ;
        RECT -206.265 -84.195 -205.485 -84.180 ;
        RECT -201.735 -84.195 -200.955 -84.180 ;
        RECT -196.345 -84.195 -191.035 -82.825 ;
        RECT -186.425 -84.180 -181.115 -82.825 ;
        RECT -186.425 -84.195 -185.645 -84.180 ;
        RECT -181.895 -84.195 -181.115 -84.180 ;
        RECT -176.505 -82.830 -175.725 -82.825 ;
        RECT -175.660 -82.830 -172.210 -82.820 ;
        RECT -165.980 -82.825 -162.040 -82.820 ;
        RECT -156.020 -82.825 -152.000 -82.820 ;
        RECT -146.140 -82.825 -142.200 -82.820 ;
        RECT -136.100 -82.825 -132.160 -82.820 ;
        RECT -126.300 -82.825 -122.360 -82.820 ;
        RECT -116.340 -82.825 -112.320 -82.820 ;
        RECT -106.460 -82.825 -102.520 -82.820 ;
        RECT -171.975 -82.830 -171.195 -82.825 ;
        RECT -176.505 -84.195 -171.195 -82.830 ;
        RECT -166.585 -84.180 -161.275 -82.825 ;
        RECT -166.585 -84.195 -165.805 -84.180 ;
        RECT -162.055 -84.195 -161.275 -84.180 ;
        RECT -156.665 -84.195 -151.355 -82.825 ;
        RECT -146.745 -84.180 -141.435 -82.825 ;
        RECT -146.745 -84.195 -145.965 -84.180 ;
        RECT -142.215 -84.195 -141.435 -84.180 ;
        RECT -136.825 -84.180 -131.515 -82.825 ;
        RECT -136.825 -84.195 -136.045 -84.180 ;
        RECT -132.295 -84.195 -131.515 -84.180 ;
        RECT -126.905 -84.180 -121.595 -82.825 ;
        RECT -126.905 -84.195 -126.125 -84.180 ;
        RECT -122.375 -84.195 -121.595 -84.180 ;
        RECT -116.985 -84.195 -111.675 -82.825 ;
        RECT -107.065 -84.180 -101.755 -82.825 ;
        RECT -107.065 -84.195 -106.285 -84.180 ;
        RECT -102.535 -84.195 -101.755 -84.180 ;
        RECT -97.145 -82.830 -96.365 -82.825 ;
        RECT -96.300 -82.830 -92.850 -82.820 ;
        RECT -86.620 -82.825 -82.680 -82.820 ;
        RECT -76.660 -82.825 -72.640 -82.820 ;
        RECT -66.780 -82.825 -62.840 -82.820 ;
        RECT -56.780 -82.825 -52.710 -82.820 ;
        RECT -46.940 -82.825 -43.000 -82.820 ;
        RECT -36.980 -82.825 -32.960 -82.820 ;
        RECT -27.100 -82.825 -23.160 -82.820 ;
        RECT -92.615 -82.830 -91.835 -82.825 ;
        RECT -97.145 -84.195 -91.835 -82.830 ;
        RECT -87.225 -84.180 -81.915 -82.825 ;
        RECT -87.225 -84.195 -86.445 -84.180 ;
        RECT -82.695 -84.195 -81.915 -84.180 ;
        RECT -77.305 -84.195 -71.995 -82.825 ;
        RECT -67.385 -84.180 -62.075 -82.825 ;
        RECT -67.385 -84.195 -66.605 -84.180 ;
        RECT -62.855 -84.195 -62.075 -84.180 ;
        RECT -57.465 -84.190 -52.155 -82.825 ;
        RECT -57.465 -84.195 -56.685 -84.190 ;
        RECT -52.935 -84.195 -52.155 -84.190 ;
        RECT -47.545 -84.180 -42.235 -82.825 ;
        RECT -47.545 -84.195 -46.765 -84.180 ;
        RECT -43.015 -84.195 -42.235 -84.180 ;
        RECT -37.625 -84.195 -32.315 -82.825 ;
        RECT -27.705 -84.180 -22.395 -82.825 ;
        RECT -27.705 -84.195 -26.925 -84.180 ;
        RECT -23.175 -84.195 -22.395 -84.180 ;
        RECT -17.785 -82.830 -17.005 -82.825 ;
        RECT -16.940 -82.830 -13.490 -82.820 ;
        RECT -7.260 -82.825 -3.320 -82.820 ;
        RECT 2.700 -82.825 6.720 -82.820 ;
        RECT 12.580 -82.825 16.520 -82.820 ;
        RECT -13.255 -82.830 -12.475 -82.825 ;
        RECT -17.785 -84.195 -12.475 -82.830 ;
        RECT -7.865 -84.180 -2.555 -82.825 ;
        RECT -7.865 -84.195 -7.085 -84.180 ;
        RECT -3.335 -84.195 -2.555 -84.180 ;
        RECT 2.055 -84.195 7.365 -82.825 ;
        RECT 11.975 -84.180 17.285 -82.825 ;
        RECT 11.975 -84.195 12.755 -84.180 ;
        RECT 16.505 -84.195 17.285 -84.180 ;
        RECT -275.060 -84.200 -271.040 -84.195 ;
        RECT -255.140 -84.200 -251.300 -84.195 ;
        RECT -235.380 -84.200 -231.360 -84.195 ;
        RECT -195.700 -84.200 -191.680 -84.195 ;
        RECT -175.780 -84.200 -171.940 -84.195 ;
        RECT -156.020 -84.200 -152.000 -84.195 ;
        RECT -116.340 -84.200 -112.320 -84.195 ;
        RECT -96.420 -84.200 -92.580 -84.195 ;
        RECT -76.660 -84.200 -72.640 -84.195 ;
        RECT -36.980 -84.200 -32.960 -84.195 ;
        RECT -17.060 -84.200 -13.220 -84.195 ;
        RECT 2.700 -84.200 6.720 -84.195 ;
        RECT -291.640 -172.445 -287.680 -172.440 ;
        RECT -281.720 -172.445 -277.760 -172.440 ;
        RECT -271.800 -172.445 -267.840 -172.440 ;
        RECT -261.880 -172.445 -257.920 -172.440 ;
        RECT -251.960 -172.445 -248.000 -172.440 ;
        RECT -242.040 -172.445 -238.080 -172.440 ;
        RECT -232.120 -172.445 -228.160 -172.440 ;
        RECT -222.200 -172.445 -218.240 -172.440 ;
        RECT -212.280 -172.445 -208.320 -172.440 ;
        RECT -202.360 -172.445 -198.400 -172.440 ;
        RECT -192.440 -172.445 -188.480 -172.440 ;
        RECT -182.520 -172.445 -178.560 -172.440 ;
        RECT -172.600 -172.445 -168.640 -172.440 ;
        RECT -162.680 -172.445 -158.720 -172.440 ;
        RECT -152.760 -172.445 -148.800 -172.440 ;
        RECT -142.840 -172.445 -138.880 -172.440 ;
        RECT -132.920 -172.445 -128.960 -172.440 ;
        RECT -123.000 -172.445 -119.040 -172.440 ;
        RECT -113.080 -172.445 -109.120 -172.440 ;
        RECT -103.160 -172.445 -99.200 -172.440 ;
        RECT -93.240 -172.445 -89.280 -172.440 ;
        RECT -83.320 -172.445 -79.360 -172.440 ;
        RECT -73.400 -172.445 -69.440 -172.440 ;
        RECT -63.480 -172.445 -59.520 -172.440 ;
        RECT -53.560 -172.445 -49.600 -172.440 ;
        RECT -43.640 -172.445 -39.680 -172.440 ;
        RECT -33.720 -172.445 -29.760 -172.440 ;
        RECT -23.800 -172.445 -19.840 -172.440 ;
        RECT -13.880 -172.445 -9.920 -172.440 ;
        RECT -3.960 -172.445 0.000 -172.440 ;
        RECT 5.960 -172.445 9.920 -172.440 ;
        RECT 15.880 -172.445 19.840 -172.440 ;
        RECT -292.345 -173.815 -287.035 -172.445 ;
        RECT -282.425 -173.815 -277.115 -172.445 ;
        RECT -272.505 -173.815 -267.195 -172.445 ;
        RECT -262.585 -173.815 -257.275 -172.445 ;
        RECT -252.665 -173.815 -247.355 -172.445 ;
        RECT -242.745 -173.815 -237.435 -172.445 ;
        RECT -232.825 -173.815 -227.515 -172.445 ;
        RECT -222.905 -173.815 -217.595 -172.445 ;
        RECT -212.985 -173.815 -207.675 -172.445 ;
        RECT -203.065 -173.815 -197.755 -172.445 ;
        RECT -193.145 -173.815 -187.835 -172.445 ;
        RECT -183.225 -173.815 -177.915 -172.445 ;
        RECT -173.305 -173.815 -167.995 -172.445 ;
        RECT -163.385 -173.815 -158.075 -172.445 ;
        RECT -153.465 -173.815 -148.155 -172.445 ;
        RECT -143.545 -173.815 -138.235 -172.445 ;
        RECT -133.625 -173.815 -128.315 -172.445 ;
        RECT -123.705 -173.815 -118.395 -172.445 ;
        RECT -113.785 -173.815 -108.475 -172.445 ;
        RECT -103.865 -173.815 -98.555 -172.445 ;
        RECT -93.945 -173.815 -88.635 -172.445 ;
        RECT -84.025 -173.815 -78.715 -172.445 ;
        RECT -74.105 -173.815 -68.795 -172.445 ;
        RECT -64.185 -173.815 -58.875 -172.445 ;
        RECT -54.265 -173.815 -48.955 -172.445 ;
        RECT -44.345 -173.815 -39.035 -172.445 ;
        RECT -34.425 -173.815 -29.115 -172.445 ;
        RECT -24.505 -173.815 -19.195 -172.445 ;
        RECT -14.585 -173.815 -9.275 -172.445 ;
        RECT -4.665 -173.815 0.645 -172.445 ;
        RECT 5.255 -173.815 10.565 -172.445 ;
        RECT 15.175 -173.815 20.485 -172.445 ;
        RECT -291.640 -173.820 -287.680 -173.815 ;
        RECT -281.720 -173.820 -277.760 -173.815 ;
        RECT -271.800 -173.820 -267.840 -173.815 ;
        RECT -261.880 -173.820 -257.920 -173.815 ;
        RECT -251.960 -173.820 -248.000 -173.815 ;
        RECT -242.040 -173.820 -238.080 -173.815 ;
        RECT -232.120 -173.820 -228.160 -173.815 ;
        RECT -222.200 -173.820 -218.240 -173.815 ;
        RECT -212.280 -173.820 -208.320 -173.815 ;
        RECT -202.360 -173.820 -198.400 -173.815 ;
        RECT -192.440 -173.820 -188.480 -173.815 ;
        RECT -182.520 -173.820 -178.560 -173.815 ;
        RECT -172.600 -173.820 -168.640 -173.815 ;
        RECT -162.680 -173.820 -158.720 -173.815 ;
        RECT -152.760 -173.820 -148.800 -173.815 ;
        RECT -142.840 -173.820 -138.880 -173.815 ;
        RECT -132.920 -173.820 -128.960 -173.815 ;
        RECT -123.000 -173.820 -119.040 -173.815 ;
        RECT -113.080 -173.820 -109.120 -173.815 ;
        RECT -103.160 -173.820 -99.200 -173.815 ;
        RECT -93.240 -173.820 -89.280 -173.815 ;
        RECT -83.320 -173.820 -79.360 -173.815 ;
        RECT -73.400 -173.820 -69.440 -173.815 ;
        RECT -63.480 -173.820 -59.520 -173.815 ;
        RECT -53.560 -173.820 -49.600 -173.815 ;
        RECT -43.640 -173.820 -39.680 -173.815 ;
        RECT -33.720 -173.820 -29.760 -173.815 ;
        RECT -23.800 -173.820 -19.840 -173.815 ;
        RECT -13.880 -173.820 -9.920 -173.815 ;
        RECT -3.960 -173.820 0.000 -173.815 ;
        RECT 5.960 -173.820 9.920 -173.815 ;
        RECT 15.880 -173.820 19.840 -173.815 ;
        RECT -285.270 -174.355 -285.100 -174.165 ;
        RECT -284.360 -174.355 -284.190 -174.165 ;
        RECT -275.350 -174.355 -275.180 -174.165 ;
        RECT -274.440 -174.355 -274.270 -174.165 ;
        RECT -265.430 -174.355 -265.260 -174.165 ;
        RECT -264.520 -174.355 -264.350 -174.165 ;
        RECT -255.510 -174.355 -255.340 -174.165 ;
        RECT -254.600 -174.355 -254.430 -174.165 ;
        RECT -245.590 -174.355 -245.420 -174.165 ;
        RECT -244.680 -174.355 -244.510 -174.165 ;
        RECT -235.670 -174.355 -235.500 -174.165 ;
        RECT -234.760 -174.355 -234.590 -174.165 ;
        RECT -225.750 -174.355 -225.580 -174.165 ;
        RECT -224.840 -174.355 -224.670 -174.165 ;
        RECT -215.830 -174.355 -215.660 -174.165 ;
        RECT -214.920 -174.355 -214.750 -174.165 ;
        RECT -205.910 -174.355 -205.740 -174.165 ;
        RECT -205.000 -174.355 -204.830 -174.165 ;
        RECT -195.990 -174.355 -195.820 -174.165 ;
        RECT -195.080 -174.355 -194.910 -174.165 ;
        RECT -186.070 -174.355 -185.900 -174.165 ;
        RECT -185.160 -174.355 -184.990 -174.165 ;
        RECT -176.150 -174.355 -175.980 -174.165 ;
        RECT -175.240 -174.355 -175.070 -174.165 ;
        RECT -166.230 -174.355 -166.060 -174.165 ;
        RECT -165.320 -174.355 -165.150 -174.165 ;
        RECT -156.310 -174.355 -156.140 -174.165 ;
        RECT -155.400 -174.355 -155.230 -174.165 ;
        RECT -146.390 -174.355 -146.220 -174.165 ;
        RECT -145.480 -174.355 -145.310 -174.165 ;
        RECT -136.470 -174.355 -136.300 -174.165 ;
        RECT -135.560 -174.355 -135.390 -174.165 ;
        RECT -126.550 -174.355 -126.380 -174.165 ;
        RECT -125.640 -174.355 -125.470 -174.165 ;
        RECT -116.630 -174.355 -116.460 -174.165 ;
        RECT -115.720 -174.355 -115.550 -174.165 ;
        RECT -106.710 -174.355 -106.540 -174.165 ;
        RECT -105.800 -174.355 -105.630 -174.165 ;
        RECT -96.790 -174.355 -96.620 -174.165 ;
        RECT -95.880 -174.355 -95.710 -174.165 ;
        RECT -86.870 -174.355 -86.700 -174.165 ;
        RECT -85.960 -174.355 -85.790 -174.165 ;
        RECT -76.950 -174.355 -76.780 -174.165 ;
        RECT -76.040 -174.355 -75.870 -174.165 ;
        RECT -67.030 -174.355 -66.860 -174.165 ;
        RECT -66.120 -174.355 -65.950 -174.165 ;
        RECT -57.110 -174.355 -56.940 -174.165 ;
        RECT -56.200 -174.355 -56.030 -174.165 ;
        RECT -47.190 -174.355 -47.020 -174.165 ;
        RECT -46.280 -174.355 -46.110 -174.165 ;
        RECT -37.270 -174.355 -37.100 -174.165 ;
        RECT -36.360 -174.355 -36.190 -174.165 ;
        RECT -27.350 -174.355 -27.180 -174.165 ;
        RECT -26.440 -174.355 -26.270 -174.165 ;
        RECT -17.430 -174.355 -17.260 -174.165 ;
        RECT -16.520 -174.355 -16.350 -174.165 ;
        RECT -7.510 -174.355 -7.340 -174.165 ;
        RECT -6.600 -174.355 -6.430 -174.165 ;
        RECT 2.410 -174.355 2.580 -174.165 ;
        RECT 3.320 -174.355 3.490 -174.165 ;
        RECT 12.330 -174.355 12.500 -174.165 ;
        RECT 13.240 -174.355 13.410 -174.165 ;
        RECT -286.335 -174.360 -284.985 -174.355 ;
        RECT -284.475 -174.360 -283.125 -174.355 ;
        RECT -286.335 -175.260 -283.125 -174.360 ;
        RECT -286.335 -175.265 -284.985 -175.260 ;
        RECT -284.475 -175.265 -283.125 -175.260 ;
        RECT -276.415 -174.360 -275.065 -174.355 ;
        RECT -274.555 -174.360 -273.205 -174.355 ;
        RECT -276.415 -175.260 -273.205 -174.360 ;
        RECT -276.415 -175.265 -275.065 -175.260 ;
        RECT -274.555 -175.265 -273.205 -175.260 ;
        RECT -266.495 -174.360 -265.145 -174.355 ;
        RECT -264.635 -174.360 -263.285 -174.355 ;
        RECT -266.495 -175.260 -263.285 -174.360 ;
        RECT -266.495 -175.265 -265.145 -175.260 ;
        RECT -264.635 -175.265 -263.285 -175.260 ;
        RECT -256.575 -174.360 -255.225 -174.355 ;
        RECT -254.715 -174.360 -253.365 -174.355 ;
        RECT -256.575 -175.260 -253.365 -174.360 ;
        RECT -256.575 -175.265 -255.225 -175.260 ;
        RECT -254.715 -175.265 -253.365 -175.260 ;
        RECT -246.655 -174.360 -245.305 -174.355 ;
        RECT -244.795 -174.360 -243.445 -174.355 ;
        RECT -246.655 -175.260 -243.445 -174.360 ;
        RECT -246.655 -175.265 -245.305 -175.260 ;
        RECT -244.795 -175.265 -243.445 -175.260 ;
        RECT -236.735 -174.360 -235.385 -174.355 ;
        RECT -234.875 -174.360 -233.525 -174.355 ;
        RECT -236.735 -175.260 -233.525 -174.360 ;
        RECT -236.735 -175.265 -235.385 -175.260 ;
        RECT -234.875 -175.265 -233.525 -175.260 ;
        RECT -226.815 -174.360 -225.465 -174.355 ;
        RECT -224.955 -174.360 -223.605 -174.355 ;
        RECT -226.815 -175.260 -223.605 -174.360 ;
        RECT -226.815 -175.265 -225.465 -175.260 ;
        RECT -224.955 -175.265 -223.605 -175.260 ;
        RECT -216.895 -174.360 -215.545 -174.355 ;
        RECT -215.035 -174.360 -213.685 -174.355 ;
        RECT -216.895 -175.260 -213.685 -174.360 ;
        RECT -216.895 -175.265 -215.545 -175.260 ;
        RECT -215.035 -175.265 -213.685 -175.260 ;
        RECT -206.975 -174.360 -205.625 -174.355 ;
        RECT -205.115 -174.360 -203.765 -174.355 ;
        RECT -206.975 -175.260 -203.765 -174.360 ;
        RECT -206.975 -175.265 -205.625 -175.260 ;
        RECT -205.115 -175.265 -203.765 -175.260 ;
        RECT -197.055 -174.360 -195.705 -174.355 ;
        RECT -195.195 -174.360 -193.845 -174.355 ;
        RECT -197.055 -175.260 -193.845 -174.360 ;
        RECT -197.055 -175.265 -195.705 -175.260 ;
        RECT -195.195 -175.265 -193.845 -175.260 ;
        RECT -187.135 -174.360 -185.785 -174.355 ;
        RECT -185.275 -174.360 -183.925 -174.355 ;
        RECT -187.135 -175.260 -183.925 -174.360 ;
        RECT -187.135 -175.265 -185.785 -175.260 ;
        RECT -185.275 -175.265 -183.925 -175.260 ;
        RECT -177.215 -174.360 -175.865 -174.355 ;
        RECT -175.355 -174.360 -174.005 -174.355 ;
        RECT -177.215 -175.260 -174.005 -174.360 ;
        RECT -177.215 -175.265 -175.865 -175.260 ;
        RECT -175.355 -175.265 -174.005 -175.260 ;
        RECT -167.295 -174.360 -165.945 -174.355 ;
        RECT -165.435 -174.360 -164.085 -174.355 ;
        RECT -167.295 -175.260 -164.085 -174.360 ;
        RECT -167.295 -175.265 -165.945 -175.260 ;
        RECT -165.435 -175.265 -164.085 -175.260 ;
        RECT -157.375 -174.360 -156.025 -174.355 ;
        RECT -155.515 -174.360 -154.165 -174.355 ;
        RECT -157.375 -175.260 -154.165 -174.360 ;
        RECT -157.375 -175.265 -156.025 -175.260 ;
        RECT -155.515 -175.265 -154.165 -175.260 ;
        RECT -147.455 -174.360 -146.105 -174.355 ;
        RECT -145.595 -174.360 -144.245 -174.355 ;
        RECT -147.455 -175.260 -144.245 -174.360 ;
        RECT -147.455 -175.265 -146.105 -175.260 ;
        RECT -145.595 -175.265 -144.245 -175.260 ;
        RECT -137.535 -174.360 -136.185 -174.355 ;
        RECT -135.675 -174.360 -134.325 -174.355 ;
        RECT -137.535 -175.260 -134.325 -174.360 ;
        RECT -137.535 -175.265 -136.185 -175.260 ;
        RECT -135.675 -175.265 -134.325 -175.260 ;
        RECT -127.615 -174.360 -126.265 -174.355 ;
        RECT -125.755 -174.360 -124.405 -174.355 ;
        RECT -127.615 -175.260 -124.405 -174.360 ;
        RECT -127.615 -175.265 -126.265 -175.260 ;
        RECT -125.755 -175.265 -124.405 -175.260 ;
        RECT -117.695 -174.360 -116.345 -174.355 ;
        RECT -115.835 -174.360 -114.485 -174.355 ;
        RECT -117.695 -175.260 -114.485 -174.360 ;
        RECT -117.695 -175.265 -116.345 -175.260 ;
        RECT -115.835 -175.265 -114.485 -175.260 ;
        RECT -107.775 -174.360 -106.425 -174.355 ;
        RECT -105.915 -174.360 -104.565 -174.355 ;
        RECT -107.775 -175.260 -104.565 -174.360 ;
        RECT -107.775 -175.265 -106.425 -175.260 ;
        RECT -105.915 -175.265 -104.565 -175.260 ;
        RECT -97.855 -174.360 -96.505 -174.355 ;
        RECT -95.995 -174.360 -94.645 -174.355 ;
        RECT -97.855 -175.260 -94.645 -174.360 ;
        RECT -97.855 -175.265 -96.505 -175.260 ;
        RECT -95.995 -175.265 -94.645 -175.260 ;
        RECT -87.935 -174.360 -86.585 -174.355 ;
        RECT -86.075 -174.360 -84.725 -174.355 ;
        RECT -87.935 -175.260 -84.725 -174.360 ;
        RECT -87.935 -175.265 -86.585 -175.260 ;
        RECT -86.075 -175.265 -84.725 -175.260 ;
        RECT -78.015 -174.360 -76.665 -174.355 ;
        RECT -76.155 -174.360 -74.805 -174.355 ;
        RECT -78.015 -175.260 -74.805 -174.360 ;
        RECT -78.015 -175.265 -76.665 -175.260 ;
        RECT -76.155 -175.265 -74.805 -175.260 ;
        RECT -68.095 -174.360 -66.745 -174.355 ;
        RECT -66.235 -174.360 -64.885 -174.355 ;
        RECT -68.095 -175.260 -64.885 -174.360 ;
        RECT -68.095 -175.265 -66.745 -175.260 ;
        RECT -66.235 -175.265 -64.885 -175.260 ;
        RECT -58.175 -174.360 -56.825 -174.355 ;
        RECT -56.315 -174.360 -54.965 -174.355 ;
        RECT -58.175 -175.260 -54.965 -174.360 ;
        RECT -58.175 -175.265 -56.825 -175.260 ;
        RECT -56.315 -175.265 -54.965 -175.260 ;
        RECT -48.255 -174.360 -46.905 -174.355 ;
        RECT -46.395 -174.360 -45.045 -174.355 ;
        RECT -48.255 -175.260 -45.045 -174.360 ;
        RECT -48.255 -175.265 -46.905 -175.260 ;
        RECT -46.395 -175.265 -45.045 -175.260 ;
        RECT -38.335 -174.360 -36.985 -174.355 ;
        RECT -36.475 -174.360 -35.125 -174.355 ;
        RECT -38.335 -175.260 -35.125 -174.360 ;
        RECT -38.335 -175.265 -36.985 -175.260 ;
        RECT -36.475 -175.265 -35.125 -175.260 ;
        RECT -28.415 -174.360 -27.065 -174.355 ;
        RECT -26.555 -174.360 -25.205 -174.355 ;
        RECT -28.415 -175.260 -25.205 -174.360 ;
        RECT -28.415 -175.265 -27.065 -175.260 ;
        RECT -26.555 -175.265 -25.205 -175.260 ;
        RECT -18.495 -174.360 -17.145 -174.355 ;
        RECT -16.635 -174.360 -15.285 -174.355 ;
        RECT -18.495 -175.260 -15.285 -174.360 ;
        RECT -18.495 -175.265 -17.145 -175.260 ;
        RECT -16.635 -175.265 -15.285 -175.260 ;
        RECT -8.575 -174.360 -7.225 -174.355 ;
        RECT -6.715 -174.360 -5.365 -174.355 ;
        RECT -8.575 -175.260 -5.365 -174.360 ;
        RECT -8.575 -175.265 -7.225 -175.260 ;
        RECT -6.715 -175.265 -5.365 -175.260 ;
        RECT 1.345 -174.360 2.695 -174.355 ;
        RECT 3.205 -174.360 4.555 -174.355 ;
        RECT 1.345 -175.260 4.555 -174.360 ;
        RECT 1.345 -175.265 2.695 -175.260 ;
        RECT 3.205 -175.265 4.555 -175.260 ;
        RECT 11.265 -174.360 12.615 -174.355 ;
        RECT 13.125 -174.360 14.475 -174.355 ;
        RECT 11.265 -175.260 14.475 -174.360 ;
        RECT 11.265 -175.265 12.615 -175.260 ;
        RECT 13.125 -175.265 14.475 -175.260 ;
        RECT -291.295 -175.960 -289.945 -175.955 ;
        RECT -289.435 -175.960 -288.085 -175.955 ;
        RECT -291.295 -176.860 -288.085 -175.960 ;
        RECT -291.295 -176.865 -289.945 -176.860 ;
        RECT -289.435 -176.865 -288.085 -176.860 ;
        RECT -281.375 -175.960 -280.025 -175.955 ;
        RECT -279.515 -175.960 -278.165 -175.955 ;
        RECT -281.375 -176.860 -278.165 -175.960 ;
        RECT -281.375 -176.865 -280.025 -176.860 ;
        RECT -279.515 -176.865 -278.165 -176.860 ;
        RECT -271.455 -175.960 -270.105 -175.955 ;
        RECT -269.595 -175.960 -268.245 -175.955 ;
        RECT -271.455 -176.860 -268.245 -175.960 ;
        RECT -271.455 -176.865 -270.105 -176.860 ;
        RECT -269.595 -176.865 -268.245 -176.860 ;
        RECT -261.535 -175.960 -260.185 -175.955 ;
        RECT -259.675 -175.960 -258.325 -175.955 ;
        RECT -261.535 -176.860 -258.325 -175.960 ;
        RECT -261.535 -176.865 -260.185 -176.860 ;
        RECT -259.675 -176.865 -258.325 -176.860 ;
        RECT -251.615 -175.960 -250.265 -175.955 ;
        RECT -249.755 -175.960 -248.405 -175.955 ;
        RECT -251.615 -176.860 -248.405 -175.960 ;
        RECT -251.615 -176.865 -250.265 -176.860 ;
        RECT -249.755 -176.865 -248.405 -176.860 ;
        RECT -241.695 -175.960 -240.345 -175.955 ;
        RECT -239.835 -175.960 -238.485 -175.955 ;
        RECT -241.695 -176.860 -238.485 -175.960 ;
        RECT -241.695 -176.865 -240.345 -176.860 ;
        RECT -239.835 -176.865 -238.485 -176.860 ;
        RECT -231.775 -175.960 -230.425 -175.955 ;
        RECT -229.915 -175.960 -228.565 -175.955 ;
        RECT -231.775 -176.860 -228.565 -175.960 ;
        RECT -231.775 -176.865 -230.425 -176.860 ;
        RECT -229.915 -176.865 -228.565 -176.860 ;
        RECT -221.855 -175.960 -220.505 -175.955 ;
        RECT -219.995 -175.960 -218.645 -175.955 ;
        RECT -221.855 -176.860 -218.645 -175.960 ;
        RECT -221.855 -176.865 -220.505 -176.860 ;
        RECT -219.995 -176.865 -218.645 -176.860 ;
        RECT -211.935 -175.960 -210.585 -175.955 ;
        RECT -210.075 -175.960 -208.725 -175.955 ;
        RECT -211.935 -176.860 -208.725 -175.960 ;
        RECT -211.935 -176.865 -210.585 -176.860 ;
        RECT -210.075 -176.865 -208.725 -176.860 ;
        RECT -202.015 -175.960 -200.665 -175.955 ;
        RECT -200.155 -175.960 -198.805 -175.955 ;
        RECT -202.015 -176.860 -198.805 -175.960 ;
        RECT -202.015 -176.865 -200.665 -176.860 ;
        RECT -200.155 -176.865 -198.805 -176.860 ;
        RECT -192.095 -175.960 -190.745 -175.955 ;
        RECT -190.235 -175.960 -188.885 -175.955 ;
        RECT -192.095 -176.860 -188.885 -175.960 ;
        RECT -192.095 -176.865 -190.745 -176.860 ;
        RECT -190.235 -176.865 -188.885 -176.860 ;
        RECT -182.175 -175.960 -180.825 -175.955 ;
        RECT -180.315 -175.960 -178.965 -175.955 ;
        RECT -182.175 -176.860 -178.965 -175.960 ;
        RECT -182.175 -176.865 -180.825 -176.860 ;
        RECT -180.315 -176.865 -178.965 -176.860 ;
        RECT -172.255 -175.960 -170.905 -175.955 ;
        RECT -170.395 -175.960 -169.045 -175.955 ;
        RECT -172.255 -176.860 -169.045 -175.960 ;
        RECT -172.255 -176.865 -170.905 -176.860 ;
        RECT -170.395 -176.865 -169.045 -176.860 ;
        RECT -162.335 -175.960 -160.985 -175.955 ;
        RECT -160.475 -175.960 -159.125 -175.955 ;
        RECT -162.335 -176.860 -159.125 -175.960 ;
        RECT -162.335 -176.865 -160.985 -176.860 ;
        RECT -160.475 -176.865 -159.125 -176.860 ;
        RECT -152.415 -175.960 -151.065 -175.955 ;
        RECT -150.555 -175.960 -149.205 -175.955 ;
        RECT -152.415 -176.860 -149.205 -175.960 ;
        RECT -152.415 -176.865 -151.065 -176.860 ;
        RECT -150.555 -176.865 -149.205 -176.860 ;
        RECT -142.495 -175.960 -141.145 -175.955 ;
        RECT -140.635 -175.960 -139.285 -175.955 ;
        RECT -142.495 -176.860 -139.285 -175.960 ;
        RECT -142.495 -176.865 -141.145 -176.860 ;
        RECT -140.635 -176.865 -139.285 -176.860 ;
        RECT -132.575 -175.960 -131.225 -175.955 ;
        RECT -130.715 -175.960 -129.365 -175.955 ;
        RECT -132.575 -176.860 -129.365 -175.960 ;
        RECT -132.575 -176.865 -131.225 -176.860 ;
        RECT -130.715 -176.865 -129.365 -176.860 ;
        RECT -122.655 -175.960 -121.305 -175.955 ;
        RECT -120.795 -175.960 -119.445 -175.955 ;
        RECT -122.655 -176.860 -119.445 -175.960 ;
        RECT -122.655 -176.865 -121.305 -176.860 ;
        RECT -120.795 -176.865 -119.445 -176.860 ;
        RECT -112.735 -175.960 -111.385 -175.955 ;
        RECT -110.875 -175.960 -109.525 -175.955 ;
        RECT -112.735 -176.860 -109.525 -175.960 ;
        RECT -112.735 -176.865 -111.385 -176.860 ;
        RECT -110.875 -176.865 -109.525 -176.860 ;
        RECT -102.815 -175.960 -101.465 -175.955 ;
        RECT -100.955 -175.960 -99.605 -175.955 ;
        RECT -102.815 -176.860 -99.605 -175.960 ;
        RECT -102.815 -176.865 -101.465 -176.860 ;
        RECT -100.955 -176.865 -99.605 -176.860 ;
        RECT -92.895 -175.960 -91.545 -175.955 ;
        RECT -91.035 -175.960 -89.685 -175.955 ;
        RECT -92.895 -176.860 -89.685 -175.960 ;
        RECT -92.895 -176.865 -91.545 -176.860 ;
        RECT -91.035 -176.865 -89.685 -176.860 ;
        RECT -82.975 -175.960 -81.625 -175.955 ;
        RECT -81.115 -175.960 -79.765 -175.955 ;
        RECT -82.975 -176.860 -79.765 -175.960 ;
        RECT -82.975 -176.865 -81.625 -176.860 ;
        RECT -81.115 -176.865 -79.765 -176.860 ;
        RECT -73.055 -175.960 -71.705 -175.955 ;
        RECT -71.195 -175.960 -69.845 -175.955 ;
        RECT -73.055 -176.860 -69.845 -175.960 ;
        RECT -73.055 -176.865 -71.705 -176.860 ;
        RECT -71.195 -176.865 -69.845 -176.860 ;
        RECT -63.135 -175.960 -61.785 -175.955 ;
        RECT -61.275 -175.960 -59.925 -175.955 ;
        RECT -63.135 -176.860 -59.925 -175.960 ;
        RECT -63.135 -176.865 -61.785 -176.860 ;
        RECT -61.275 -176.865 -59.925 -176.860 ;
        RECT -53.215 -175.960 -51.865 -175.955 ;
        RECT -51.355 -175.960 -50.005 -175.955 ;
        RECT -53.215 -176.860 -50.005 -175.960 ;
        RECT -53.215 -176.865 -51.865 -176.860 ;
        RECT -51.355 -176.865 -50.005 -176.860 ;
        RECT -43.295 -175.960 -41.945 -175.955 ;
        RECT -41.435 -175.960 -40.085 -175.955 ;
        RECT -43.295 -176.860 -40.085 -175.960 ;
        RECT -43.295 -176.865 -41.945 -176.860 ;
        RECT -41.435 -176.865 -40.085 -176.860 ;
        RECT -33.375 -175.960 -32.025 -175.955 ;
        RECT -31.515 -175.960 -30.165 -175.955 ;
        RECT -33.375 -176.860 -30.165 -175.960 ;
        RECT -33.375 -176.865 -32.025 -176.860 ;
        RECT -31.515 -176.865 -30.165 -176.860 ;
        RECT -23.455 -175.960 -22.105 -175.955 ;
        RECT -21.595 -175.960 -20.245 -175.955 ;
        RECT -23.455 -176.860 -20.245 -175.960 ;
        RECT -23.455 -176.865 -22.105 -176.860 ;
        RECT -21.595 -176.865 -20.245 -176.860 ;
        RECT -13.535 -175.960 -12.185 -175.955 ;
        RECT -11.675 -175.960 -10.325 -175.955 ;
        RECT -13.535 -176.860 -10.325 -175.960 ;
        RECT -13.535 -176.865 -12.185 -176.860 ;
        RECT -11.675 -176.865 -10.325 -176.860 ;
        RECT -3.615 -175.960 -2.265 -175.955 ;
        RECT -1.755 -175.960 -0.405 -175.955 ;
        RECT -3.615 -176.860 -0.405 -175.960 ;
        RECT -3.615 -176.865 -2.265 -176.860 ;
        RECT -1.755 -176.865 -0.405 -176.860 ;
        RECT 6.305 -175.960 7.655 -175.955 ;
        RECT 8.165 -175.960 9.515 -175.955 ;
        RECT 6.305 -176.860 9.515 -175.960 ;
        RECT 6.305 -176.865 7.655 -176.860 ;
        RECT 8.165 -176.865 9.515 -176.860 ;
        RECT 16.225 -175.960 17.575 -175.955 ;
        RECT 18.085 -175.960 19.435 -175.955 ;
        RECT 16.225 -176.860 19.435 -175.960 ;
        RECT 16.225 -176.865 17.575 -176.860 ;
        RECT 18.085 -176.865 19.435 -176.860 ;
        RECT -290.230 -177.055 -290.060 -176.865 ;
        RECT -289.320 -177.055 -289.150 -176.865 ;
        RECT -280.310 -177.055 -280.140 -176.865 ;
        RECT -279.400 -177.055 -279.230 -176.865 ;
        RECT -270.390 -177.055 -270.220 -176.865 ;
        RECT -269.480 -177.055 -269.310 -176.865 ;
        RECT -260.470 -177.055 -260.300 -176.865 ;
        RECT -259.560 -177.055 -259.390 -176.865 ;
        RECT -250.550 -177.055 -250.380 -176.865 ;
        RECT -249.640 -177.055 -249.470 -176.865 ;
        RECT -240.630 -177.055 -240.460 -176.865 ;
        RECT -239.720 -177.055 -239.550 -176.865 ;
        RECT -230.710 -177.055 -230.540 -176.865 ;
        RECT -229.800 -177.055 -229.630 -176.865 ;
        RECT -220.790 -177.055 -220.620 -176.865 ;
        RECT -219.880 -177.055 -219.710 -176.865 ;
        RECT -210.870 -177.055 -210.700 -176.865 ;
        RECT -209.960 -177.055 -209.790 -176.865 ;
        RECT -200.950 -177.055 -200.780 -176.865 ;
        RECT -200.040 -177.055 -199.870 -176.865 ;
        RECT -191.030 -177.055 -190.860 -176.865 ;
        RECT -190.120 -177.055 -189.950 -176.865 ;
        RECT -181.110 -177.055 -180.940 -176.865 ;
        RECT -180.200 -177.055 -180.030 -176.865 ;
        RECT -171.190 -177.055 -171.020 -176.865 ;
        RECT -170.280 -177.055 -170.110 -176.865 ;
        RECT -161.270 -177.055 -161.100 -176.865 ;
        RECT -160.360 -177.055 -160.190 -176.865 ;
        RECT -151.350 -177.055 -151.180 -176.865 ;
        RECT -150.440 -177.055 -150.270 -176.865 ;
        RECT -141.430 -177.055 -141.260 -176.865 ;
        RECT -140.520 -177.055 -140.350 -176.865 ;
        RECT -131.510 -177.055 -131.340 -176.865 ;
        RECT -130.600 -177.055 -130.430 -176.865 ;
        RECT -121.590 -177.055 -121.420 -176.865 ;
        RECT -120.680 -177.055 -120.510 -176.865 ;
        RECT -111.670 -177.055 -111.500 -176.865 ;
        RECT -110.760 -177.055 -110.590 -176.865 ;
        RECT -101.750 -177.055 -101.580 -176.865 ;
        RECT -100.840 -177.055 -100.670 -176.865 ;
        RECT -91.830 -177.055 -91.660 -176.865 ;
        RECT -90.920 -177.055 -90.750 -176.865 ;
        RECT -81.910 -177.055 -81.740 -176.865 ;
        RECT -81.000 -177.055 -80.830 -176.865 ;
        RECT -71.990 -177.055 -71.820 -176.865 ;
        RECT -71.080 -177.055 -70.910 -176.865 ;
        RECT -62.070 -177.055 -61.900 -176.865 ;
        RECT -61.160 -177.055 -60.990 -176.865 ;
        RECT -52.150 -177.055 -51.980 -176.865 ;
        RECT -51.240 -177.055 -51.070 -176.865 ;
        RECT -42.230 -177.055 -42.060 -176.865 ;
        RECT -41.320 -177.055 -41.150 -176.865 ;
        RECT -32.310 -177.055 -32.140 -176.865 ;
        RECT -31.400 -177.055 -31.230 -176.865 ;
        RECT -22.390 -177.055 -22.220 -176.865 ;
        RECT -21.480 -177.055 -21.310 -176.865 ;
        RECT -12.470 -177.055 -12.300 -176.865 ;
        RECT -11.560 -177.055 -11.390 -176.865 ;
        RECT -2.550 -177.055 -2.380 -176.865 ;
        RECT -1.640 -177.055 -1.470 -176.865 ;
        RECT 7.370 -177.055 7.540 -176.865 ;
        RECT 8.280 -177.055 8.450 -176.865 ;
        RECT 17.290 -177.055 17.460 -176.865 ;
        RECT 18.200 -177.055 18.370 -176.865 ;
        RECT -284.945 -177.400 -284.515 -177.385 ;
        RECT -275.025 -177.400 -274.595 -177.385 ;
        RECT -265.105 -177.400 -264.675 -177.385 ;
        RECT -255.185 -177.400 -254.755 -177.385 ;
        RECT -245.265 -177.400 -244.835 -177.385 ;
        RECT -235.345 -177.400 -234.915 -177.385 ;
        RECT -225.425 -177.400 -224.995 -177.385 ;
        RECT -215.505 -177.400 -215.075 -177.385 ;
        RECT -205.585 -177.400 -205.155 -177.385 ;
        RECT -195.665 -177.400 -195.235 -177.385 ;
        RECT -185.745 -177.400 -185.315 -177.385 ;
        RECT -175.825 -177.400 -175.395 -177.385 ;
        RECT -165.905 -177.400 -165.475 -177.385 ;
        RECT -155.985 -177.400 -155.555 -177.385 ;
        RECT -146.065 -177.400 -145.635 -177.385 ;
        RECT -136.145 -177.400 -135.715 -177.385 ;
        RECT -126.225 -177.400 -125.795 -177.385 ;
        RECT -116.305 -177.400 -115.875 -177.385 ;
        RECT -106.385 -177.400 -105.955 -177.385 ;
        RECT -96.465 -177.400 -96.035 -177.385 ;
        RECT -86.545 -177.400 -86.115 -177.385 ;
        RECT -76.625 -177.400 -76.195 -177.385 ;
        RECT -66.705 -177.400 -66.275 -177.385 ;
        RECT -56.785 -177.400 -56.355 -177.385 ;
        RECT -46.865 -177.400 -46.435 -177.385 ;
        RECT -36.945 -177.400 -36.515 -177.385 ;
        RECT -27.025 -177.400 -26.595 -177.385 ;
        RECT -17.105 -177.400 -16.675 -177.385 ;
        RECT -7.185 -177.400 -6.755 -177.385 ;
        RECT 2.735 -177.400 3.165 -177.385 ;
        RECT 12.655 -177.400 13.085 -177.385 ;
        RECT -286.780 -177.405 -282.840 -177.400 ;
        RECT -276.820 -177.405 -272.800 -177.400 ;
        RECT -266.940 -177.405 -263.000 -177.400 ;
        RECT -287.385 -178.760 -282.075 -177.405 ;
        RECT -287.385 -178.775 -286.605 -178.760 ;
        RECT -282.855 -178.775 -282.075 -178.760 ;
        RECT -277.465 -178.775 -272.155 -177.405 ;
        RECT -267.545 -178.760 -262.235 -177.405 ;
        RECT -267.545 -178.775 -266.765 -178.760 ;
        RECT -263.015 -178.775 -262.235 -178.760 ;
        RECT -257.625 -177.410 -256.845 -177.405 ;
        RECT -256.780 -177.410 -253.330 -177.400 ;
        RECT -247.100 -177.405 -243.160 -177.400 ;
        RECT -237.140 -177.405 -233.120 -177.400 ;
        RECT -227.260 -177.405 -223.320 -177.400 ;
        RECT -217.260 -177.405 -213.190 -177.400 ;
        RECT -207.420 -177.405 -203.480 -177.400 ;
        RECT -197.460 -177.405 -193.440 -177.400 ;
        RECT -187.580 -177.405 -183.640 -177.400 ;
        RECT -253.095 -177.410 -252.315 -177.405 ;
        RECT -257.625 -178.775 -252.315 -177.410 ;
        RECT -247.705 -178.760 -242.395 -177.405 ;
        RECT -247.705 -178.775 -246.925 -178.760 ;
        RECT -243.175 -178.775 -242.395 -178.760 ;
        RECT -237.785 -178.775 -232.475 -177.405 ;
        RECT -227.865 -178.760 -222.555 -177.405 ;
        RECT -227.865 -178.775 -227.085 -178.760 ;
        RECT -223.335 -178.775 -222.555 -178.760 ;
        RECT -217.945 -178.770 -212.635 -177.405 ;
        RECT -217.945 -178.775 -217.165 -178.770 ;
        RECT -213.415 -178.775 -212.635 -178.770 ;
        RECT -208.025 -178.760 -202.715 -177.405 ;
        RECT -208.025 -178.775 -207.245 -178.760 ;
        RECT -203.495 -178.775 -202.715 -178.760 ;
        RECT -198.105 -178.775 -192.795 -177.405 ;
        RECT -188.185 -178.760 -182.875 -177.405 ;
        RECT -188.185 -178.775 -187.405 -178.760 ;
        RECT -183.655 -178.775 -182.875 -178.760 ;
        RECT -178.265 -177.410 -177.485 -177.405 ;
        RECT -177.420 -177.410 -173.970 -177.400 ;
        RECT -167.740 -177.405 -163.800 -177.400 ;
        RECT -157.780 -177.405 -153.760 -177.400 ;
        RECT -147.900 -177.405 -143.960 -177.400 ;
        RECT -137.860 -177.405 -133.920 -177.400 ;
        RECT -128.060 -177.405 -124.120 -177.400 ;
        RECT -118.100 -177.405 -114.080 -177.400 ;
        RECT -108.220 -177.405 -104.280 -177.400 ;
        RECT -173.735 -177.410 -172.955 -177.405 ;
        RECT -178.265 -178.775 -172.955 -177.410 ;
        RECT -168.345 -178.760 -163.035 -177.405 ;
        RECT -168.345 -178.775 -167.565 -178.760 ;
        RECT -163.815 -178.775 -163.035 -178.760 ;
        RECT -158.425 -178.775 -153.115 -177.405 ;
        RECT -148.505 -178.760 -143.195 -177.405 ;
        RECT -148.505 -178.775 -147.725 -178.760 ;
        RECT -143.975 -178.775 -143.195 -178.760 ;
        RECT -138.585 -178.760 -133.275 -177.405 ;
        RECT -138.585 -178.775 -137.805 -178.760 ;
        RECT -134.055 -178.775 -133.275 -178.760 ;
        RECT -128.665 -178.760 -123.355 -177.405 ;
        RECT -128.665 -178.775 -127.885 -178.760 ;
        RECT -124.135 -178.775 -123.355 -178.760 ;
        RECT -118.745 -178.775 -113.435 -177.405 ;
        RECT -108.825 -178.760 -103.515 -177.405 ;
        RECT -108.825 -178.775 -108.045 -178.760 ;
        RECT -104.295 -178.775 -103.515 -178.760 ;
        RECT -98.905 -177.410 -98.125 -177.405 ;
        RECT -98.060 -177.410 -94.610 -177.400 ;
        RECT -88.380 -177.405 -84.440 -177.400 ;
        RECT -78.420 -177.405 -74.400 -177.400 ;
        RECT -68.540 -177.405 -64.600 -177.400 ;
        RECT -58.540 -177.405 -54.470 -177.400 ;
        RECT -48.700 -177.405 -44.760 -177.400 ;
        RECT -38.740 -177.405 -34.720 -177.400 ;
        RECT -28.860 -177.405 -24.920 -177.400 ;
        RECT -94.375 -177.410 -93.595 -177.405 ;
        RECT -98.905 -178.775 -93.595 -177.410 ;
        RECT -88.985 -178.760 -83.675 -177.405 ;
        RECT -88.985 -178.775 -88.205 -178.760 ;
        RECT -84.455 -178.775 -83.675 -178.760 ;
        RECT -79.065 -178.775 -73.755 -177.405 ;
        RECT -69.145 -178.760 -63.835 -177.405 ;
        RECT -69.145 -178.775 -68.365 -178.760 ;
        RECT -64.615 -178.775 -63.835 -178.760 ;
        RECT -59.225 -178.770 -53.915 -177.405 ;
        RECT -59.225 -178.775 -58.445 -178.770 ;
        RECT -54.695 -178.775 -53.915 -178.770 ;
        RECT -49.305 -178.760 -43.995 -177.405 ;
        RECT -49.305 -178.775 -48.525 -178.760 ;
        RECT -44.775 -178.775 -43.995 -178.760 ;
        RECT -39.385 -178.775 -34.075 -177.405 ;
        RECT -29.465 -178.760 -24.155 -177.405 ;
        RECT -29.465 -178.775 -28.685 -178.760 ;
        RECT -24.935 -178.775 -24.155 -178.760 ;
        RECT -19.545 -177.410 -18.765 -177.405 ;
        RECT -18.700 -177.410 -15.250 -177.400 ;
        RECT -9.020 -177.405 -5.080 -177.400 ;
        RECT 0.940 -177.405 4.960 -177.400 ;
        RECT 10.820 -177.405 14.760 -177.400 ;
        RECT -15.015 -177.410 -14.235 -177.405 ;
        RECT -19.545 -178.775 -14.235 -177.410 ;
        RECT -9.625 -178.760 -4.315 -177.405 ;
        RECT -9.625 -178.775 -8.845 -178.760 ;
        RECT -5.095 -178.775 -4.315 -178.760 ;
        RECT 0.295 -178.775 5.605 -177.405 ;
        RECT 10.215 -178.760 15.525 -177.405 ;
        RECT 10.215 -178.775 10.995 -178.760 ;
        RECT 14.745 -178.775 15.525 -178.760 ;
        RECT -276.820 -178.780 -272.800 -178.775 ;
        RECT -256.900 -178.780 -253.060 -178.775 ;
        RECT -237.140 -178.780 -233.120 -178.775 ;
        RECT -197.460 -178.780 -193.440 -178.775 ;
        RECT -177.540 -178.780 -173.700 -178.775 ;
        RECT -157.780 -178.780 -153.760 -178.775 ;
        RECT -118.100 -178.780 -114.080 -178.775 ;
        RECT -98.180 -178.780 -94.340 -178.775 ;
        RECT -78.420 -178.780 -74.400 -178.775 ;
        RECT -38.740 -178.780 -34.720 -178.775 ;
        RECT -18.820 -178.780 -14.980 -178.775 ;
        RECT 0.940 -178.780 4.960 -178.775 ;
      LAYER li1 ;
        RECT -288.125 94.615 -287.955 95.140 ;
        RECT -286.500 94.725 -286.040 94.895 ;
        RECT -288.505 94.285 -287.955 94.615 ;
        RECT -288.125 93.760 -287.955 94.285 ;
        RECT -286.415 94.000 -286.125 94.725 ;
        RECT -284.585 94.615 -284.415 95.140 ;
        RECT -278.205 94.615 -278.035 95.140 ;
        RECT -276.580 94.725 -276.120 94.895 ;
        RECT -284.585 94.285 -284.035 94.615 ;
        RECT -278.585 94.285 -278.035 94.615 ;
        RECT -284.585 93.760 -284.415 94.285 ;
        RECT -278.205 93.760 -278.035 94.285 ;
        RECT -276.495 94.000 -276.205 94.725 ;
        RECT -274.665 94.615 -274.495 95.140 ;
        RECT -268.285 94.615 -268.115 95.140 ;
        RECT -266.660 94.725 -266.200 94.895 ;
        RECT -274.665 94.285 -274.115 94.615 ;
        RECT -268.665 94.285 -268.115 94.615 ;
        RECT -274.665 93.760 -274.495 94.285 ;
        RECT -268.285 93.760 -268.115 94.285 ;
        RECT -266.575 94.000 -266.285 94.725 ;
        RECT -264.745 94.615 -264.575 95.140 ;
        RECT -258.365 94.615 -258.195 95.140 ;
        RECT -256.740 94.725 -256.280 94.895 ;
        RECT -264.745 94.285 -264.195 94.615 ;
        RECT -258.745 94.285 -258.195 94.615 ;
        RECT -264.745 93.760 -264.575 94.285 ;
        RECT -258.365 93.760 -258.195 94.285 ;
        RECT -256.655 94.000 -256.365 94.725 ;
        RECT -254.825 94.615 -254.655 95.140 ;
        RECT -248.445 94.615 -248.275 95.140 ;
        RECT -246.820 94.725 -246.360 94.895 ;
        RECT -254.825 94.285 -254.275 94.615 ;
        RECT -248.825 94.285 -248.275 94.615 ;
        RECT -254.825 93.760 -254.655 94.285 ;
        RECT -248.445 93.760 -248.275 94.285 ;
        RECT -246.735 94.000 -246.445 94.725 ;
        RECT -244.905 94.615 -244.735 95.140 ;
        RECT -238.525 94.615 -238.355 95.140 ;
        RECT -236.900 94.725 -236.440 94.895 ;
        RECT -244.905 94.285 -244.355 94.615 ;
        RECT -238.905 94.285 -238.355 94.615 ;
        RECT -244.905 93.760 -244.735 94.285 ;
        RECT -238.525 93.760 -238.355 94.285 ;
        RECT -236.815 94.000 -236.525 94.725 ;
        RECT -234.985 94.615 -234.815 95.140 ;
        RECT -228.605 94.615 -228.435 95.140 ;
        RECT -226.980 94.725 -226.520 94.895 ;
        RECT -234.985 94.285 -234.435 94.615 ;
        RECT -228.985 94.285 -228.435 94.615 ;
        RECT -234.985 93.760 -234.815 94.285 ;
        RECT -228.605 93.760 -228.435 94.285 ;
        RECT -226.895 94.000 -226.605 94.725 ;
        RECT -225.065 94.615 -224.895 95.140 ;
        RECT -218.685 94.615 -218.515 95.140 ;
        RECT -217.060 94.725 -216.600 94.895 ;
        RECT -225.065 94.285 -224.515 94.615 ;
        RECT -219.065 94.285 -218.515 94.615 ;
        RECT -225.065 93.760 -224.895 94.285 ;
        RECT -218.685 93.760 -218.515 94.285 ;
        RECT -216.975 94.000 -216.685 94.725 ;
        RECT -215.145 94.615 -214.975 95.140 ;
        RECT -208.765 94.615 -208.595 95.140 ;
        RECT -207.140 94.725 -206.680 94.895 ;
        RECT -215.145 94.285 -214.595 94.615 ;
        RECT -209.145 94.285 -208.595 94.615 ;
        RECT -215.145 93.760 -214.975 94.285 ;
        RECT -208.765 93.760 -208.595 94.285 ;
        RECT -207.055 94.000 -206.765 94.725 ;
        RECT -205.225 94.615 -205.055 95.140 ;
        RECT -198.845 94.615 -198.675 95.140 ;
        RECT -197.220 94.725 -196.760 94.895 ;
        RECT -205.225 94.285 -204.675 94.615 ;
        RECT -199.225 94.285 -198.675 94.615 ;
        RECT -205.225 93.760 -205.055 94.285 ;
        RECT -198.845 93.760 -198.675 94.285 ;
        RECT -197.135 94.000 -196.845 94.725 ;
        RECT -195.305 94.615 -195.135 95.140 ;
        RECT -188.925 94.615 -188.755 95.140 ;
        RECT -187.300 94.725 -186.840 94.895 ;
        RECT -195.305 94.285 -194.755 94.615 ;
        RECT -189.305 94.285 -188.755 94.615 ;
        RECT -195.305 93.760 -195.135 94.285 ;
        RECT -188.925 93.760 -188.755 94.285 ;
        RECT -187.215 94.000 -186.925 94.725 ;
        RECT -185.385 94.615 -185.215 95.140 ;
        RECT -179.005 94.615 -178.835 95.140 ;
        RECT -177.380 94.725 -176.920 94.895 ;
        RECT -185.385 94.285 -184.835 94.615 ;
        RECT -179.385 94.285 -178.835 94.615 ;
        RECT -185.385 93.760 -185.215 94.285 ;
        RECT -179.005 93.760 -178.835 94.285 ;
        RECT -177.295 94.000 -177.005 94.725 ;
        RECT -175.465 94.615 -175.295 95.140 ;
        RECT -169.085 94.615 -168.915 95.140 ;
        RECT -167.460 94.725 -167.000 94.895 ;
        RECT -175.465 94.285 -174.915 94.615 ;
        RECT -169.465 94.285 -168.915 94.615 ;
        RECT -175.465 93.760 -175.295 94.285 ;
        RECT -169.085 93.760 -168.915 94.285 ;
        RECT -167.375 94.000 -167.085 94.725 ;
        RECT -165.545 94.615 -165.375 95.140 ;
        RECT -159.165 94.615 -158.995 95.140 ;
        RECT -157.540 94.725 -157.080 94.895 ;
        RECT -165.545 94.285 -164.995 94.615 ;
        RECT -159.545 94.285 -158.995 94.615 ;
        RECT -165.545 93.760 -165.375 94.285 ;
        RECT -159.165 93.760 -158.995 94.285 ;
        RECT -157.455 94.000 -157.165 94.725 ;
        RECT -155.625 94.615 -155.455 95.140 ;
        RECT -149.245 94.615 -149.075 95.140 ;
        RECT -147.620 94.725 -147.160 94.895 ;
        RECT -155.625 94.285 -155.075 94.615 ;
        RECT -149.625 94.285 -149.075 94.615 ;
        RECT -155.625 93.760 -155.455 94.285 ;
        RECT -149.245 93.760 -149.075 94.285 ;
        RECT -147.535 94.000 -147.245 94.725 ;
        RECT -145.705 94.615 -145.535 95.140 ;
        RECT -139.325 94.615 -139.155 95.140 ;
        RECT -137.700 94.725 -137.240 94.895 ;
        RECT -145.705 94.285 -145.155 94.615 ;
        RECT -139.705 94.285 -139.155 94.615 ;
        RECT -145.705 93.760 -145.535 94.285 ;
        RECT -139.325 93.760 -139.155 94.285 ;
        RECT -137.615 94.000 -137.325 94.725 ;
        RECT -135.785 94.615 -135.615 95.140 ;
        RECT -129.405 94.615 -129.235 95.140 ;
        RECT -127.780 94.725 -127.320 94.895 ;
        RECT -135.785 94.285 -135.235 94.615 ;
        RECT -129.785 94.285 -129.235 94.615 ;
        RECT -135.785 93.760 -135.615 94.285 ;
        RECT -129.405 93.760 -129.235 94.285 ;
        RECT -127.695 94.000 -127.405 94.725 ;
        RECT -125.865 94.615 -125.695 95.140 ;
        RECT -119.485 94.615 -119.315 95.140 ;
        RECT -117.860 94.725 -117.400 94.895 ;
        RECT -125.865 94.285 -125.315 94.615 ;
        RECT -119.865 94.285 -119.315 94.615 ;
        RECT -125.865 93.760 -125.695 94.285 ;
        RECT -119.485 93.760 -119.315 94.285 ;
        RECT -117.775 94.000 -117.485 94.725 ;
        RECT -115.945 94.615 -115.775 95.140 ;
        RECT -109.565 94.615 -109.395 95.140 ;
        RECT -107.940 94.725 -107.480 94.895 ;
        RECT -115.945 94.285 -115.395 94.615 ;
        RECT -109.945 94.285 -109.395 94.615 ;
        RECT -115.945 93.760 -115.775 94.285 ;
        RECT -109.565 93.760 -109.395 94.285 ;
        RECT -107.855 94.000 -107.565 94.725 ;
        RECT -106.025 94.615 -105.855 95.140 ;
        RECT -99.645 94.615 -99.475 95.140 ;
        RECT -98.020 94.725 -97.560 94.895 ;
        RECT -106.025 94.285 -105.475 94.615 ;
        RECT -100.025 94.285 -99.475 94.615 ;
        RECT -106.025 93.760 -105.855 94.285 ;
        RECT -99.645 93.760 -99.475 94.285 ;
        RECT -97.935 94.000 -97.645 94.725 ;
        RECT -96.105 94.615 -95.935 95.140 ;
        RECT -89.725 94.615 -89.555 95.140 ;
        RECT -88.100 94.725 -87.640 94.895 ;
        RECT -96.105 94.285 -95.555 94.615 ;
        RECT -90.105 94.285 -89.555 94.615 ;
        RECT -96.105 93.760 -95.935 94.285 ;
        RECT -89.725 93.760 -89.555 94.285 ;
        RECT -88.015 94.000 -87.725 94.725 ;
        RECT -86.185 94.615 -86.015 95.140 ;
        RECT -79.805 94.615 -79.635 95.140 ;
        RECT -78.180 94.725 -77.720 94.895 ;
        RECT -86.185 94.285 -85.635 94.615 ;
        RECT -80.185 94.285 -79.635 94.615 ;
        RECT -86.185 93.760 -86.015 94.285 ;
        RECT -79.805 93.760 -79.635 94.285 ;
        RECT -78.095 94.000 -77.805 94.725 ;
        RECT -76.265 94.615 -76.095 95.140 ;
        RECT -69.885 94.615 -69.715 95.140 ;
        RECT -68.260 94.725 -67.800 94.895 ;
        RECT -76.265 94.285 -75.715 94.615 ;
        RECT -70.265 94.285 -69.715 94.615 ;
        RECT -76.265 93.760 -76.095 94.285 ;
        RECT -69.885 93.760 -69.715 94.285 ;
        RECT -68.175 94.000 -67.885 94.725 ;
        RECT -66.345 94.615 -66.175 95.140 ;
        RECT -59.965 94.615 -59.795 95.140 ;
        RECT -58.340 94.725 -57.880 94.895 ;
        RECT -66.345 94.285 -65.795 94.615 ;
        RECT -60.345 94.285 -59.795 94.615 ;
        RECT -66.345 93.760 -66.175 94.285 ;
        RECT -59.965 93.760 -59.795 94.285 ;
        RECT -58.255 94.000 -57.965 94.725 ;
        RECT -56.425 94.615 -56.255 95.140 ;
        RECT -50.045 94.615 -49.875 95.140 ;
        RECT -48.420 94.725 -47.960 94.895 ;
        RECT -56.425 94.285 -55.875 94.615 ;
        RECT -50.425 94.285 -49.875 94.615 ;
        RECT -56.425 93.760 -56.255 94.285 ;
        RECT -50.045 93.760 -49.875 94.285 ;
        RECT -48.335 94.000 -48.045 94.725 ;
        RECT -46.505 94.615 -46.335 95.140 ;
        RECT -40.125 94.615 -39.955 95.140 ;
        RECT -38.500 94.725 -38.040 94.895 ;
        RECT -46.505 94.285 -45.955 94.615 ;
        RECT -40.505 94.285 -39.955 94.615 ;
        RECT -46.505 93.760 -46.335 94.285 ;
        RECT -40.125 93.760 -39.955 94.285 ;
        RECT -38.415 94.000 -38.125 94.725 ;
        RECT -36.585 94.615 -36.415 95.140 ;
        RECT -30.205 94.615 -30.035 95.140 ;
        RECT -28.580 94.725 -28.120 94.895 ;
        RECT -36.585 94.285 -36.035 94.615 ;
        RECT -30.585 94.285 -30.035 94.615 ;
        RECT -36.585 93.760 -36.415 94.285 ;
        RECT -30.205 93.760 -30.035 94.285 ;
        RECT -28.495 94.000 -28.205 94.725 ;
        RECT -26.665 94.615 -26.495 95.140 ;
        RECT -20.285 94.615 -20.115 95.140 ;
        RECT -18.660 94.725 -18.200 94.895 ;
        RECT -26.665 94.285 -26.115 94.615 ;
        RECT -20.665 94.285 -20.115 94.615 ;
        RECT -26.665 93.760 -26.495 94.285 ;
        RECT -20.285 93.760 -20.115 94.285 ;
        RECT -18.575 94.000 -18.285 94.725 ;
        RECT -16.745 94.615 -16.575 95.140 ;
        RECT -10.365 94.615 -10.195 95.140 ;
        RECT -8.740 94.725 -8.280 94.895 ;
        RECT -16.745 94.285 -16.195 94.615 ;
        RECT -10.745 94.285 -10.195 94.615 ;
        RECT -16.745 93.760 -16.575 94.285 ;
        RECT -10.365 93.760 -10.195 94.285 ;
        RECT -8.655 94.000 -8.365 94.725 ;
        RECT -6.825 94.615 -6.655 95.140 ;
        RECT -0.445 94.615 -0.275 95.140 ;
        RECT 1.180 94.725 1.640 94.895 ;
        RECT -6.825 94.285 -6.275 94.615 ;
        RECT -0.825 94.285 -0.275 94.615 ;
        RECT -6.825 93.760 -6.655 94.285 ;
        RECT -0.445 93.760 -0.275 94.285 ;
        RECT 1.265 94.000 1.555 94.725 ;
        RECT 3.095 94.615 3.265 95.140 ;
        RECT 9.475 94.615 9.645 95.140 ;
        RECT 11.100 94.725 11.560 94.895 ;
        RECT 3.095 94.285 3.645 94.615 ;
        RECT 9.095 94.285 9.645 94.615 ;
        RECT 3.095 93.760 3.265 94.285 ;
        RECT 9.475 93.760 9.645 94.285 ;
        RECT 11.185 94.000 11.475 94.725 ;
        RECT 13.015 94.615 13.185 95.140 ;
        RECT 19.395 94.615 19.565 95.140 ;
        RECT 21.020 94.725 21.480 94.895 ;
        RECT 13.015 94.285 13.565 94.615 ;
        RECT 19.015 94.285 19.565 94.615 ;
        RECT 13.015 93.760 13.185 94.285 ;
        RECT 19.395 93.760 19.565 94.285 ;
        RECT 21.105 94.000 21.395 94.725 ;
        RECT 22.935 94.615 23.105 95.140 ;
        RECT 22.935 94.285 23.485 94.615 ;
        RECT 22.935 93.760 23.105 94.285 ;
        RECT -282.920 93.245 -279.700 93.415 ;
        RECT -273.000 93.245 -269.780 93.415 ;
        RECT -263.080 93.245 -259.860 93.415 ;
        RECT -253.160 93.245 -249.940 93.415 ;
        RECT -243.240 93.245 -240.020 93.415 ;
        RECT -233.320 93.245 -230.100 93.415 ;
        RECT -223.400 93.245 -220.180 93.415 ;
        RECT -213.480 93.245 -210.260 93.415 ;
        RECT -203.560 93.245 -200.340 93.415 ;
        RECT -193.640 93.245 -190.420 93.415 ;
        RECT -183.720 93.245 -180.500 93.415 ;
        RECT -173.800 93.245 -170.580 93.415 ;
        RECT -163.880 93.245 -160.660 93.415 ;
        RECT -153.960 93.245 -150.740 93.415 ;
        RECT -144.040 93.245 -140.820 93.415 ;
        RECT -134.120 93.245 -130.900 93.415 ;
        RECT -124.200 93.245 -120.980 93.415 ;
        RECT -114.280 93.245 -111.060 93.415 ;
        RECT -104.360 93.245 -101.140 93.415 ;
        RECT -94.440 93.245 -91.220 93.415 ;
        RECT -84.520 93.245 -81.300 93.415 ;
        RECT -74.600 93.245 -71.380 93.415 ;
        RECT -64.680 93.245 -61.460 93.415 ;
        RECT -54.760 93.245 -51.540 93.415 ;
        RECT -44.840 93.245 -41.620 93.415 ;
        RECT -34.920 93.245 -31.700 93.415 ;
        RECT -25.000 93.245 -21.780 93.415 ;
        RECT -15.080 93.245 -11.860 93.415 ;
        RECT -5.160 93.245 -1.940 93.415 ;
        RECT 4.760 93.245 7.980 93.415 ;
        RECT 14.680 93.245 17.900 93.415 ;
        RECT -281.935 92.445 -281.625 93.245 ;
        RECT -281.455 92.520 -281.165 93.245 ;
        RECT -280.995 92.445 -280.685 93.245 ;
        RECT -272.015 92.445 -271.705 93.245 ;
        RECT -271.535 92.520 -271.245 93.245 ;
        RECT -271.075 92.445 -270.765 93.245 ;
        RECT -262.095 92.445 -261.785 93.245 ;
        RECT -261.615 92.520 -261.325 93.245 ;
        RECT -261.155 92.445 -260.845 93.245 ;
        RECT -252.175 92.445 -251.865 93.245 ;
        RECT -251.695 92.520 -251.405 93.245 ;
        RECT -251.235 92.445 -250.925 93.245 ;
        RECT -242.255 92.445 -241.945 93.245 ;
        RECT -241.775 92.520 -241.485 93.245 ;
        RECT -241.315 92.445 -241.005 93.245 ;
        RECT -232.335 92.445 -232.025 93.245 ;
        RECT -231.855 92.520 -231.565 93.245 ;
        RECT -231.395 92.445 -231.085 93.245 ;
        RECT -222.415 92.445 -222.105 93.245 ;
        RECT -221.935 92.520 -221.645 93.245 ;
        RECT -221.475 92.445 -221.165 93.245 ;
        RECT -212.495 92.445 -212.185 93.245 ;
        RECT -212.015 92.520 -211.725 93.245 ;
        RECT -211.555 92.445 -211.245 93.245 ;
        RECT -202.575 92.445 -202.265 93.245 ;
        RECT -202.095 92.520 -201.805 93.245 ;
        RECT -201.635 92.445 -201.325 93.245 ;
        RECT -192.655 92.445 -192.345 93.245 ;
        RECT -192.175 92.520 -191.885 93.245 ;
        RECT -191.715 92.445 -191.405 93.245 ;
        RECT -182.735 92.445 -182.425 93.245 ;
        RECT -182.255 92.520 -181.965 93.245 ;
        RECT -181.795 92.445 -181.485 93.245 ;
        RECT -172.815 92.445 -172.505 93.245 ;
        RECT -172.335 92.520 -172.045 93.245 ;
        RECT -171.875 92.445 -171.565 93.245 ;
        RECT -162.895 92.445 -162.585 93.245 ;
        RECT -162.415 92.520 -162.125 93.245 ;
        RECT -161.955 92.445 -161.645 93.245 ;
        RECT -152.975 92.445 -152.665 93.245 ;
        RECT -152.495 92.520 -152.205 93.245 ;
        RECT -152.035 92.445 -151.725 93.245 ;
        RECT -143.055 92.445 -142.745 93.245 ;
        RECT -142.575 92.520 -142.285 93.245 ;
        RECT -142.115 92.445 -141.805 93.245 ;
        RECT -133.135 92.445 -132.825 93.245 ;
        RECT -132.655 92.520 -132.365 93.245 ;
        RECT -132.195 92.445 -131.885 93.245 ;
        RECT -123.215 92.445 -122.905 93.245 ;
        RECT -122.735 92.520 -122.445 93.245 ;
        RECT -122.275 92.445 -121.965 93.245 ;
        RECT -113.295 92.445 -112.985 93.245 ;
        RECT -112.815 92.520 -112.525 93.245 ;
        RECT -112.355 92.445 -112.045 93.245 ;
        RECT -103.375 92.445 -103.065 93.245 ;
        RECT -102.895 92.520 -102.605 93.245 ;
        RECT -102.435 92.445 -102.125 93.245 ;
        RECT -93.455 92.445 -93.145 93.245 ;
        RECT -92.975 92.520 -92.685 93.245 ;
        RECT -92.515 92.445 -92.205 93.245 ;
        RECT -83.535 92.445 -83.225 93.245 ;
        RECT -83.055 92.520 -82.765 93.245 ;
        RECT -82.595 92.445 -82.285 93.245 ;
        RECT -73.615 92.445 -73.305 93.245 ;
        RECT -73.135 92.520 -72.845 93.245 ;
        RECT -72.675 92.445 -72.365 93.245 ;
        RECT -63.695 92.445 -63.385 93.245 ;
        RECT -63.215 92.520 -62.925 93.245 ;
        RECT -62.755 92.445 -62.445 93.245 ;
        RECT -53.775 92.445 -53.465 93.245 ;
        RECT -53.295 92.520 -53.005 93.245 ;
        RECT -52.835 92.445 -52.525 93.245 ;
        RECT -43.855 92.445 -43.545 93.245 ;
        RECT -43.375 92.520 -43.085 93.245 ;
        RECT -42.915 92.445 -42.605 93.245 ;
        RECT -33.935 92.445 -33.625 93.245 ;
        RECT -33.455 92.520 -33.165 93.245 ;
        RECT -32.995 92.445 -32.685 93.245 ;
        RECT -24.015 92.445 -23.705 93.245 ;
        RECT -23.535 92.520 -23.245 93.245 ;
        RECT -23.075 92.445 -22.765 93.245 ;
        RECT -14.095 92.445 -13.785 93.245 ;
        RECT -13.615 92.520 -13.325 93.245 ;
        RECT -13.155 92.445 -12.845 93.245 ;
        RECT -4.175 92.445 -3.865 93.245 ;
        RECT -3.695 92.520 -3.405 93.245 ;
        RECT -3.235 92.445 -2.925 93.245 ;
        RECT 5.745 92.445 6.055 93.245 ;
        RECT 6.225 92.520 6.515 93.245 ;
        RECT 6.685 92.445 6.995 93.245 ;
        RECT 15.665 92.445 15.975 93.245 ;
        RECT 16.145 92.520 16.435 93.245 ;
        RECT 16.605 92.445 16.915 93.245 ;
        RECT -286.895 90.695 -286.585 91.495 ;
        RECT -286.415 90.695 -286.125 91.420 ;
        RECT -285.955 90.695 -285.645 91.495 ;
        RECT -276.975 90.695 -276.665 91.495 ;
        RECT -276.495 90.695 -276.205 91.420 ;
        RECT -276.035 90.695 -275.725 91.495 ;
        RECT -267.055 90.695 -266.745 91.495 ;
        RECT -266.575 90.695 -266.285 91.420 ;
        RECT -266.115 90.695 -265.805 91.495 ;
        RECT -257.135 90.695 -256.825 91.495 ;
        RECT -256.655 90.695 -256.365 91.420 ;
        RECT -256.195 90.695 -255.885 91.495 ;
        RECT -247.215 90.695 -246.905 91.495 ;
        RECT -246.735 90.695 -246.445 91.420 ;
        RECT -246.275 90.695 -245.965 91.495 ;
        RECT -237.295 90.695 -236.985 91.495 ;
        RECT -236.815 90.695 -236.525 91.420 ;
        RECT -236.355 90.695 -236.045 91.495 ;
        RECT -227.375 90.695 -227.065 91.495 ;
        RECT -226.895 90.695 -226.605 91.420 ;
        RECT -226.435 90.695 -226.125 91.495 ;
        RECT -217.455 90.695 -217.145 91.495 ;
        RECT -216.975 90.695 -216.685 91.420 ;
        RECT -216.515 90.695 -216.205 91.495 ;
        RECT -207.535 90.695 -207.225 91.495 ;
        RECT -207.055 90.695 -206.765 91.420 ;
        RECT -206.595 90.695 -206.285 91.495 ;
        RECT -197.615 90.695 -197.305 91.495 ;
        RECT -197.135 90.695 -196.845 91.420 ;
        RECT -196.675 90.695 -196.365 91.495 ;
        RECT -187.695 90.695 -187.385 91.495 ;
        RECT -187.215 90.695 -186.925 91.420 ;
        RECT -186.755 90.695 -186.445 91.495 ;
        RECT -177.775 90.695 -177.465 91.495 ;
        RECT -177.295 90.695 -177.005 91.420 ;
        RECT -176.835 90.695 -176.525 91.495 ;
        RECT -167.855 90.695 -167.545 91.495 ;
        RECT -167.375 90.695 -167.085 91.420 ;
        RECT -166.915 90.695 -166.605 91.495 ;
        RECT -157.935 90.695 -157.625 91.495 ;
        RECT -157.455 90.695 -157.165 91.420 ;
        RECT -156.995 90.695 -156.685 91.495 ;
        RECT -148.015 90.695 -147.705 91.495 ;
        RECT -147.535 90.695 -147.245 91.420 ;
        RECT -147.075 90.695 -146.765 91.495 ;
        RECT -138.095 90.695 -137.785 91.495 ;
        RECT -137.615 90.695 -137.325 91.420 ;
        RECT -137.155 90.695 -136.845 91.495 ;
        RECT -128.175 90.695 -127.865 91.495 ;
        RECT -127.695 90.695 -127.405 91.420 ;
        RECT -127.235 90.695 -126.925 91.495 ;
        RECT -118.255 90.695 -117.945 91.495 ;
        RECT -117.775 90.695 -117.485 91.420 ;
        RECT -117.315 90.695 -117.005 91.495 ;
        RECT -108.335 90.695 -108.025 91.495 ;
        RECT -107.855 90.695 -107.565 91.420 ;
        RECT -107.395 90.695 -107.085 91.495 ;
        RECT -98.415 90.695 -98.105 91.495 ;
        RECT -97.935 90.695 -97.645 91.420 ;
        RECT -97.475 90.695 -97.165 91.495 ;
        RECT -88.495 90.695 -88.185 91.495 ;
        RECT -88.015 90.695 -87.725 91.420 ;
        RECT -87.555 90.695 -87.245 91.495 ;
        RECT -78.575 90.695 -78.265 91.495 ;
        RECT -78.095 90.695 -77.805 91.420 ;
        RECT -77.635 90.695 -77.325 91.495 ;
        RECT -68.655 90.695 -68.345 91.495 ;
        RECT -68.175 90.695 -67.885 91.420 ;
        RECT -67.715 90.695 -67.405 91.495 ;
        RECT -58.735 90.695 -58.425 91.495 ;
        RECT -58.255 90.695 -57.965 91.420 ;
        RECT -57.795 90.695 -57.485 91.495 ;
        RECT -48.815 90.695 -48.505 91.495 ;
        RECT -48.335 90.695 -48.045 91.420 ;
        RECT -47.875 90.695 -47.565 91.495 ;
        RECT -38.895 90.695 -38.585 91.495 ;
        RECT -38.415 90.695 -38.125 91.420 ;
        RECT -37.955 90.695 -37.645 91.495 ;
        RECT -28.975 90.695 -28.665 91.495 ;
        RECT -28.495 90.695 -28.205 91.420 ;
        RECT -28.035 90.695 -27.725 91.495 ;
        RECT -19.055 90.695 -18.745 91.495 ;
        RECT -18.575 90.695 -18.285 91.420 ;
        RECT -18.115 90.695 -17.805 91.495 ;
        RECT -9.135 90.695 -8.825 91.495 ;
        RECT -8.655 90.695 -8.365 91.420 ;
        RECT -8.195 90.695 -7.885 91.495 ;
        RECT 0.785 90.695 1.095 91.495 ;
        RECT 1.265 90.695 1.555 91.420 ;
        RECT 1.725 90.695 2.035 91.495 ;
        RECT 10.705 90.695 11.015 91.495 ;
        RECT 11.185 90.695 11.475 91.420 ;
        RECT 11.645 90.695 11.955 91.495 ;
        RECT 20.625 90.695 20.935 91.495 ;
        RECT 21.105 90.695 21.395 91.420 ;
        RECT 21.565 90.695 21.875 91.495 ;
        RECT -287.880 90.525 -284.660 90.695 ;
        RECT -277.960 90.525 -274.740 90.695 ;
        RECT -268.040 90.525 -264.820 90.695 ;
        RECT -258.120 90.525 -254.900 90.695 ;
        RECT -248.200 90.525 -244.980 90.695 ;
        RECT -238.280 90.525 -235.060 90.695 ;
        RECT -228.360 90.525 -225.140 90.695 ;
        RECT -218.440 90.525 -215.220 90.695 ;
        RECT -208.520 90.525 -205.300 90.695 ;
        RECT -198.600 90.525 -195.380 90.695 ;
        RECT -188.680 90.525 -185.460 90.695 ;
        RECT -178.760 90.525 -175.540 90.695 ;
        RECT -168.840 90.525 -165.620 90.695 ;
        RECT -158.920 90.525 -155.700 90.695 ;
        RECT -149.000 90.525 -145.780 90.695 ;
        RECT -139.080 90.525 -135.860 90.695 ;
        RECT -129.160 90.525 -125.940 90.695 ;
        RECT -119.240 90.525 -116.020 90.695 ;
        RECT -109.320 90.525 -106.100 90.695 ;
        RECT -99.400 90.525 -96.180 90.695 ;
        RECT -89.480 90.525 -86.260 90.695 ;
        RECT -79.560 90.525 -76.340 90.695 ;
        RECT -69.640 90.525 -66.420 90.695 ;
        RECT -59.720 90.525 -56.500 90.695 ;
        RECT -49.800 90.525 -46.580 90.695 ;
        RECT -39.880 90.525 -36.660 90.695 ;
        RECT -29.960 90.525 -26.740 90.695 ;
        RECT -20.040 90.525 -16.820 90.695 ;
        RECT -10.120 90.525 -6.900 90.695 ;
        RECT -0.200 90.525 3.020 90.695 ;
        RECT 9.720 90.525 12.940 90.695 ;
        RECT 19.640 90.525 22.860 90.695 ;
        RECT -283.165 89.655 -282.995 90.180 ;
        RECT -283.545 89.325 -282.995 89.655 ;
        RECT -283.165 88.800 -282.995 89.325 ;
        RECT -281.455 89.305 -281.165 90.030 ;
        RECT -279.625 89.655 -279.455 90.180 ;
        RECT -273.245 89.655 -273.075 90.180 ;
        RECT -279.625 89.325 -279.075 89.655 ;
        RECT -273.625 89.325 -273.075 89.655 ;
        RECT -281.540 89.135 -281.080 89.305 ;
        RECT -279.625 88.800 -279.455 89.325 ;
        RECT -273.245 88.800 -273.075 89.325 ;
        RECT -271.535 89.305 -271.245 90.030 ;
        RECT -269.705 89.655 -269.535 90.180 ;
        RECT -263.325 89.655 -263.155 90.180 ;
        RECT -269.705 89.325 -269.155 89.655 ;
        RECT -263.705 89.325 -263.155 89.655 ;
        RECT -271.620 89.135 -271.160 89.305 ;
        RECT -269.705 88.800 -269.535 89.325 ;
        RECT -263.325 88.800 -263.155 89.325 ;
        RECT -261.615 89.305 -261.325 90.030 ;
        RECT -259.785 89.655 -259.615 90.180 ;
        RECT -253.405 89.655 -253.235 90.180 ;
        RECT -259.785 89.325 -259.235 89.655 ;
        RECT -253.785 89.325 -253.235 89.655 ;
        RECT -261.700 89.135 -261.240 89.305 ;
        RECT -259.785 88.800 -259.615 89.325 ;
        RECT -253.405 88.800 -253.235 89.325 ;
        RECT -251.695 89.305 -251.405 90.030 ;
        RECT -249.865 89.655 -249.695 90.180 ;
        RECT -243.485 89.655 -243.315 90.180 ;
        RECT -249.865 89.325 -249.315 89.655 ;
        RECT -243.865 89.325 -243.315 89.655 ;
        RECT -251.780 89.135 -251.320 89.305 ;
        RECT -249.865 88.800 -249.695 89.325 ;
        RECT -243.485 88.800 -243.315 89.325 ;
        RECT -241.775 89.305 -241.485 90.030 ;
        RECT -239.945 89.655 -239.775 90.180 ;
        RECT -233.565 89.655 -233.395 90.180 ;
        RECT -239.945 89.325 -239.395 89.655 ;
        RECT -233.945 89.325 -233.395 89.655 ;
        RECT -241.860 89.135 -241.400 89.305 ;
        RECT -239.945 88.800 -239.775 89.325 ;
        RECT -233.565 88.800 -233.395 89.325 ;
        RECT -231.855 89.305 -231.565 90.030 ;
        RECT -230.025 89.655 -229.855 90.180 ;
        RECT -223.645 89.655 -223.475 90.180 ;
        RECT -230.025 89.325 -229.475 89.655 ;
        RECT -224.025 89.325 -223.475 89.655 ;
        RECT -231.940 89.135 -231.480 89.305 ;
        RECT -230.025 88.800 -229.855 89.325 ;
        RECT -223.645 88.800 -223.475 89.325 ;
        RECT -221.935 89.305 -221.645 90.030 ;
        RECT -220.105 89.655 -219.935 90.180 ;
        RECT -213.725 89.655 -213.555 90.180 ;
        RECT -220.105 89.325 -219.555 89.655 ;
        RECT -214.105 89.325 -213.555 89.655 ;
        RECT -222.020 89.135 -221.560 89.305 ;
        RECT -220.105 88.800 -219.935 89.325 ;
        RECT -213.725 88.800 -213.555 89.325 ;
        RECT -212.015 89.305 -211.725 90.030 ;
        RECT -210.185 89.655 -210.015 90.180 ;
        RECT -203.805 89.655 -203.635 90.180 ;
        RECT -210.185 89.325 -209.635 89.655 ;
        RECT -204.185 89.325 -203.635 89.655 ;
        RECT -212.100 89.135 -211.640 89.305 ;
        RECT -210.185 88.800 -210.015 89.325 ;
        RECT -203.805 88.800 -203.635 89.325 ;
        RECT -202.095 89.305 -201.805 90.030 ;
        RECT -200.265 89.655 -200.095 90.180 ;
        RECT -193.885 89.655 -193.715 90.180 ;
        RECT -200.265 89.325 -199.715 89.655 ;
        RECT -194.265 89.325 -193.715 89.655 ;
        RECT -202.180 89.135 -201.720 89.305 ;
        RECT -200.265 88.800 -200.095 89.325 ;
        RECT -193.885 88.800 -193.715 89.325 ;
        RECT -192.175 89.305 -191.885 90.030 ;
        RECT -190.345 89.655 -190.175 90.180 ;
        RECT -183.965 89.655 -183.795 90.180 ;
        RECT -190.345 89.325 -189.795 89.655 ;
        RECT -184.345 89.325 -183.795 89.655 ;
        RECT -192.260 89.135 -191.800 89.305 ;
        RECT -190.345 88.800 -190.175 89.325 ;
        RECT -183.965 88.800 -183.795 89.325 ;
        RECT -182.255 89.305 -181.965 90.030 ;
        RECT -180.425 89.655 -180.255 90.180 ;
        RECT -174.045 89.655 -173.875 90.180 ;
        RECT -180.425 89.325 -179.875 89.655 ;
        RECT -174.425 89.325 -173.875 89.655 ;
        RECT -182.340 89.135 -181.880 89.305 ;
        RECT -180.425 88.800 -180.255 89.325 ;
        RECT -174.045 88.800 -173.875 89.325 ;
        RECT -172.335 89.305 -172.045 90.030 ;
        RECT -170.505 89.655 -170.335 90.180 ;
        RECT -164.125 89.655 -163.955 90.180 ;
        RECT -170.505 89.325 -169.955 89.655 ;
        RECT -164.505 89.325 -163.955 89.655 ;
        RECT -172.420 89.135 -171.960 89.305 ;
        RECT -170.505 88.800 -170.335 89.325 ;
        RECT -164.125 88.800 -163.955 89.325 ;
        RECT -162.415 89.305 -162.125 90.030 ;
        RECT -160.585 89.655 -160.415 90.180 ;
        RECT -154.205 89.655 -154.035 90.180 ;
        RECT -160.585 89.325 -160.035 89.655 ;
        RECT -154.585 89.325 -154.035 89.655 ;
        RECT -162.500 89.135 -162.040 89.305 ;
        RECT -160.585 88.800 -160.415 89.325 ;
        RECT -154.205 88.800 -154.035 89.325 ;
        RECT -152.495 89.305 -152.205 90.030 ;
        RECT -150.665 89.655 -150.495 90.180 ;
        RECT -144.285 89.655 -144.115 90.180 ;
        RECT -150.665 89.325 -150.115 89.655 ;
        RECT -144.665 89.325 -144.115 89.655 ;
        RECT -152.580 89.135 -152.120 89.305 ;
        RECT -150.665 88.800 -150.495 89.325 ;
        RECT -144.285 88.800 -144.115 89.325 ;
        RECT -142.575 89.305 -142.285 90.030 ;
        RECT -140.745 89.655 -140.575 90.180 ;
        RECT -134.365 89.655 -134.195 90.180 ;
        RECT -140.745 89.325 -140.195 89.655 ;
        RECT -134.745 89.325 -134.195 89.655 ;
        RECT -142.660 89.135 -142.200 89.305 ;
        RECT -140.745 88.800 -140.575 89.325 ;
        RECT -134.365 88.800 -134.195 89.325 ;
        RECT -132.655 89.305 -132.365 90.030 ;
        RECT -130.825 89.655 -130.655 90.180 ;
        RECT -124.445 89.655 -124.275 90.180 ;
        RECT -130.825 89.325 -130.275 89.655 ;
        RECT -124.825 89.325 -124.275 89.655 ;
        RECT -132.740 89.135 -132.280 89.305 ;
        RECT -130.825 88.800 -130.655 89.325 ;
        RECT -124.445 88.800 -124.275 89.325 ;
        RECT -122.735 89.305 -122.445 90.030 ;
        RECT -120.905 89.655 -120.735 90.180 ;
        RECT -114.525 89.655 -114.355 90.180 ;
        RECT -120.905 89.325 -120.355 89.655 ;
        RECT -114.905 89.325 -114.355 89.655 ;
        RECT -122.820 89.135 -122.360 89.305 ;
        RECT -120.905 88.800 -120.735 89.325 ;
        RECT -114.525 88.800 -114.355 89.325 ;
        RECT -112.815 89.305 -112.525 90.030 ;
        RECT -110.985 89.655 -110.815 90.180 ;
        RECT -104.605 89.655 -104.435 90.180 ;
        RECT -110.985 89.325 -110.435 89.655 ;
        RECT -104.985 89.325 -104.435 89.655 ;
        RECT -112.900 89.135 -112.440 89.305 ;
        RECT -110.985 88.800 -110.815 89.325 ;
        RECT -104.605 88.800 -104.435 89.325 ;
        RECT -102.895 89.305 -102.605 90.030 ;
        RECT -101.065 89.655 -100.895 90.180 ;
        RECT -94.685 89.655 -94.515 90.180 ;
        RECT -101.065 89.325 -100.515 89.655 ;
        RECT -95.065 89.325 -94.515 89.655 ;
        RECT -102.980 89.135 -102.520 89.305 ;
        RECT -101.065 88.800 -100.895 89.325 ;
        RECT -94.685 88.800 -94.515 89.325 ;
        RECT -92.975 89.305 -92.685 90.030 ;
        RECT -91.145 89.655 -90.975 90.180 ;
        RECT -84.765 89.655 -84.595 90.180 ;
        RECT -91.145 89.325 -90.595 89.655 ;
        RECT -85.145 89.325 -84.595 89.655 ;
        RECT -93.060 89.135 -92.600 89.305 ;
        RECT -91.145 88.800 -90.975 89.325 ;
        RECT -84.765 88.800 -84.595 89.325 ;
        RECT -83.055 89.305 -82.765 90.030 ;
        RECT -81.225 89.655 -81.055 90.180 ;
        RECT -74.845 89.655 -74.675 90.180 ;
        RECT -81.225 89.325 -80.675 89.655 ;
        RECT -75.225 89.325 -74.675 89.655 ;
        RECT -83.140 89.135 -82.680 89.305 ;
        RECT -81.225 88.800 -81.055 89.325 ;
        RECT -74.845 88.800 -74.675 89.325 ;
        RECT -73.135 89.305 -72.845 90.030 ;
        RECT -71.305 89.655 -71.135 90.180 ;
        RECT -64.925 89.655 -64.755 90.180 ;
        RECT -71.305 89.325 -70.755 89.655 ;
        RECT -65.305 89.325 -64.755 89.655 ;
        RECT -73.220 89.135 -72.760 89.305 ;
        RECT -71.305 88.800 -71.135 89.325 ;
        RECT -64.925 88.800 -64.755 89.325 ;
        RECT -63.215 89.305 -62.925 90.030 ;
        RECT -61.385 89.655 -61.215 90.180 ;
        RECT -55.005 89.655 -54.835 90.180 ;
        RECT -61.385 89.325 -60.835 89.655 ;
        RECT -55.385 89.325 -54.835 89.655 ;
        RECT -63.300 89.135 -62.840 89.305 ;
        RECT -61.385 88.800 -61.215 89.325 ;
        RECT -55.005 88.800 -54.835 89.325 ;
        RECT -53.295 89.305 -53.005 90.030 ;
        RECT -51.465 89.655 -51.295 90.180 ;
        RECT -45.085 89.655 -44.915 90.180 ;
        RECT -51.465 89.325 -50.915 89.655 ;
        RECT -45.465 89.325 -44.915 89.655 ;
        RECT -53.380 89.135 -52.920 89.305 ;
        RECT -51.465 88.800 -51.295 89.325 ;
        RECT -45.085 88.800 -44.915 89.325 ;
        RECT -43.375 89.305 -43.085 90.030 ;
        RECT -41.545 89.655 -41.375 90.180 ;
        RECT -35.165 89.655 -34.995 90.180 ;
        RECT -41.545 89.325 -40.995 89.655 ;
        RECT -35.545 89.325 -34.995 89.655 ;
        RECT -43.460 89.135 -43.000 89.305 ;
        RECT -41.545 88.800 -41.375 89.325 ;
        RECT -35.165 88.800 -34.995 89.325 ;
        RECT -33.455 89.305 -33.165 90.030 ;
        RECT -31.625 89.655 -31.455 90.180 ;
        RECT -25.245 89.655 -25.075 90.180 ;
        RECT -31.625 89.325 -31.075 89.655 ;
        RECT -25.625 89.325 -25.075 89.655 ;
        RECT -33.540 89.135 -33.080 89.305 ;
        RECT -31.625 88.800 -31.455 89.325 ;
        RECT -25.245 88.800 -25.075 89.325 ;
        RECT -23.535 89.305 -23.245 90.030 ;
        RECT -21.705 89.655 -21.535 90.180 ;
        RECT -15.325 89.655 -15.155 90.180 ;
        RECT -21.705 89.325 -21.155 89.655 ;
        RECT -15.705 89.325 -15.155 89.655 ;
        RECT -23.620 89.135 -23.160 89.305 ;
        RECT -21.705 88.800 -21.535 89.325 ;
        RECT -15.325 88.800 -15.155 89.325 ;
        RECT -13.615 89.305 -13.325 90.030 ;
        RECT -11.785 89.655 -11.615 90.180 ;
        RECT -5.405 89.655 -5.235 90.180 ;
        RECT -11.785 89.325 -11.235 89.655 ;
        RECT -5.785 89.325 -5.235 89.655 ;
        RECT -13.700 89.135 -13.240 89.305 ;
        RECT -11.785 88.800 -11.615 89.325 ;
        RECT -5.405 88.800 -5.235 89.325 ;
        RECT -3.695 89.305 -3.405 90.030 ;
        RECT -1.865 89.655 -1.695 90.180 ;
        RECT 4.515 89.655 4.685 90.180 ;
        RECT -1.865 89.325 -1.315 89.655 ;
        RECT 4.135 89.325 4.685 89.655 ;
        RECT -3.780 89.135 -3.320 89.305 ;
        RECT -1.865 88.800 -1.695 89.325 ;
        RECT 4.515 88.800 4.685 89.325 ;
        RECT 6.225 89.305 6.515 90.030 ;
        RECT 8.055 89.655 8.225 90.180 ;
        RECT 14.435 89.655 14.605 90.180 ;
        RECT 8.055 89.325 8.605 89.655 ;
        RECT 14.055 89.325 14.605 89.655 ;
        RECT 6.140 89.135 6.600 89.305 ;
        RECT 8.055 88.800 8.225 89.325 ;
        RECT 14.435 88.800 14.605 89.325 ;
        RECT 16.145 89.305 16.435 90.030 ;
        RECT 17.975 89.655 18.145 90.180 ;
        RECT 17.975 89.325 18.525 89.655 ;
        RECT 16.060 89.135 16.520 89.305 ;
        RECT 17.975 88.800 18.145 89.325 ;
        RECT -290.145 10.565 -289.975 11.090 ;
        RECT -288.520 10.675 -288.060 10.845 ;
        RECT -290.525 10.235 -289.975 10.565 ;
        RECT -290.145 9.710 -289.975 10.235 ;
        RECT -288.435 9.950 -288.145 10.675 ;
        RECT -286.605 10.565 -286.435 11.090 ;
        RECT -280.225 10.565 -280.055 11.090 ;
        RECT -278.600 10.675 -278.140 10.845 ;
        RECT -286.605 10.235 -286.055 10.565 ;
        RECT -280.605 10.235 -280.055 10.565 ;
        RECT -286.605 9.710 -286.435 10.235 ;
        RECT -280.225 9.710 -280.055 10.235 ;
        RECT -278.515 9.950 -278.225 10.675 ;
        RECT -276.685 10.565 -276.515 11.090 ;
        RECT -270.305 10.565 -270.135 11.090 ;
        RECT -268.680 10.675 -268.220 10.845 ;
        RECT -276.685 10.235 -276.135 10.565 ;
        RECT -270.685 10.235 -270.135 10.565 ;
        RECT -276.685 9.710 -276.515 10.235 ;
        RECT -270.305 9.710 -270.135 10.235 ;
        RECT -268.595 9.950 -268.305 10.675 ;
        RECT -266.765 10.565 -266.595 11.090 ;
        RECT -260.385 10.565 -260.215 11.090 ;
        RECT -258.760 10.675 -258.300 10.845 ;
        RECT -266.765 10.235 -266.215 10.565 ;
        RECT -260.765 10.235 -260.215 10.565 ;
        RECT -266.765 9.710 -266.595 10.235 ;
        RECT -260.385 9.710 -260.215 10.235 ;
        RECT -258.675 9.950 -258.385 10.675 ;
        RECT -256.845 10.565 -256.675 11.090 ;
        RECT -250.465 10.565 -250.295 11.090 ;
        RECT -248.840 10.675 -248.380 10.845 ;
        RECT -256.845 10.235 -256.295 10.565 ;
        RECT -250.845 10.235 -250.295 10.565 ;
        RECT -256.845 9.710 -256.675 10.235 ;
        RECT -250.465 9.710 -250.295 10.235 ;
        RECT -248.755 9.950 -248.465 10.675 ;
        RECT -246.925 10.565 -246.755 11.090 ;
        RECT -240.545 10.565 -240.375 11.090 ;
        RECT -238.920 10.675 -238.460 10.845 ;
        RECT -246.925 10.235 -246.375 10.565 ;
        RECT -240.925 10.235 -240.375 10.565 ;
        RECT -246.925 9.710 -246.755 10.235 ;
        RECT -240.545 9.710 -240.375 10.235 ;
        RECT -238.835 9.950 -238.545 10.675 ;
        RECT -237.005 10.565 -236.835 11.090 ;
        RECT -230.625 10.565 -230.455 11.090 ;
        RECT -229.000 10.675 -228.540 10.845 ;
        RECT -237.005 10.235 -236.455 10.565 ;
        RECT -231.005 10.235 -230.455 10.565 ;
        RECT -237.005 9.710 -236.835 10.235 ;
        RECT -230.625 9.710 -230.455 10.235 ;
        RECT -228.915 9.950 -228.625 10.675 ;
        RECT -227.085 10.565 -226.915 11.090 ;
        RECT -220.705 10.565 -220.535 11.090 ;
        RECT -219.080 10.675 -218.620 10.845 ;
        RECT -227.085 10.235 -226.535 10.565 ;
        RECT -221.085 10.235 -220.535 10.565 ;
        RECT -227.085 9.710 -226.915 10.235 ;
        RECT -220.705 9.710 -220.535 10.235 ;
        RECT -218.995 9.950 -218.705 10.675 ;
        RECT -217.165 10.565 -216.995 11.090 ;
        RECT -210.785 10.565 -210.615 11.090 ;
        RECT -209.160 10.675 -208.700 10.845 ;
        RECT -217.165 10.235 -216.615 10.565 ;
        RECT -211.165 10.235 -210.615 10.565 ;
        RECT -217.165 9.710 -216.995 10.235 ;
        RECT -210.785 9.710 -210.615 10.235 ;
        RECT -209.075 9.950 -208.785 10.675 ;
        RECT -207.245 10.565 -207.075 11.090 ;
        RECT -200.865 10.565 -200.695 11.090 ;
        RECT -199.240 10.675 -198.780 10.845 ;
        RECT -207.245 10.235 -206.695 10.565 ;
        RECT -201.245 10.235 -200.695 10.565 ;
        RECT -207.245 9.710 -207.075 10.235 ;
        RECT -200.865 9.710 -200.695 10.235 ;
        RECT -199.155 9.950 -198.865 10.675 ;
        RECT -197.325 10.565 -197.155 11.090 ;
        RECT -190.945 10.565 -190.775 11.090 ;
        RECT -189.320 10.675 -188.860 10.845 ;
        RECT -197.325 10.235 -196.775 10.565 ;
        RECT -191.325 10.235 -190.775 10.565 ;
        RECT -197.325 9.710 -197.155 10.235 ;
        RECT -190.945 9.710 -190.775 10.235 ;
        RECT -189.235 9.950 -188.945 10.675 ;
        RECT -187.405 10.565 -187.235 11.090 ;
        RECT -181.025 10.565 -180.855 11.090 ;
        RECT -179.400 10.675 -178.940 10.845 ;
        RECT -187.405 10.235 -186.855 10.565 ;
        RECT -181.405 10.235 -180.855 10.565 ;
        RECT -187.405 9.710 -187.235 10.235 ;
        RECT -181.025 9.710 -180.855 10.235 ;
        RECT -179.315 9.950 -179.025 10.675 ;
        RECT -177.485 10.565 -177.315 11.090 ;
        RECT -171.105 10.565 -170.935 11.090 ;
        RECT -169.480 10.675 -169.020 10.845 ;
        RECT -177.485 10.235 -176.935 10.565 ;
        RECT -171.485 10.235 -170.935 10.565 ;
        RECT -177.485 9.710 -177.315 10.235 ;
        RECT -171.105 9.710 -170.935 10.235 ;
        RECT -169.395 9.950 -169.105 10.675 ;
        RECT -167.565 10.565 -167.395 11.090 ;
        RECT -161.185 10.565 -161.015 11.090 ;
        RECT -159.560 10.675 -159.100 10.845 ;
        RECT -167.565 10.235 -167.015 10.565 ;
        RECT -161.565 10.235 -161.015 10.565 ;
        RECT -167.565 9.710 -167.395 10.235 ;
        RECT -161.185 9.710 -161.015 10.235 ;
        RECT -159.475 9.950 -159.185 10.675 ;
        RECT -157.645 10.565 -157.475 11.090 ;
        RECT -151.265 10.565 -151.095 11.090 ;
        RECT -149.640 10.675 -149.180 10.845 ;
        RECT -157.645 10.235 -157.095 10.565 ;
        RECT -151.645 10.235 -151.095 10.565 ;
        RECT -157.645 9.710 -157.475 10.235 ;
        RECT -151.265 9.710 -151.095 10.235 ;
        RECT -149.555 9.950 -149.265 10.675 ;
        RECT -147.725 10.565 -147.555 11.090 ;
        RECT -141.345 10.565 -141.175 11.090 ;
        RECT -139.720 10.675 -139.260 10.845 ;
        RECT -147.725 10.235 -147.175 10.565 ;
        RECT -141.725 10.235 -141.175 10.565 ;
        RECT -147.725 9.710 -147.555 10.235 ;
        RECT -141.345 9.710 -141.175 10.235 ;
        RECT -139.635 9.950 -139.345 10.675 ;
        RECT -137.805 10.565 -137.635 11.090 ;
        RECT -131.425 10.565 -131.255 11.090 ;
        RECT -129.800 10.675 -129.340 10.845 ;
        RECT -137.805 10.235 -137.255 10.565 ;
        RECT -131.805 10.235 -131.255 10.565 ;
        RECT -137.805 9.710 -137.635 10.235 ;
        RECT -131.425 9.710 -131.255 10.235 ;
        RECT -129.715 9.950 -129.425 10.675 ;
        RECT -127.885 10.565 -127.715 11.090 ;
        RECT -121.505 10.565 -121.335 11.090 ;
        RECT -119.880 10.675 -119.420 10.845 ;
        RECT -127.885 10.235 -127.335 10.565 ;
        RECT -121.885 10.235 -121.335 10.565 ;
        RECT -127.885 9.710 -127.715 10.235 ;
        RECT -121.505 9.710 -121.335 10.235 ;
        RECT -119.795 9.950 -119.505 10.675 ;
        RECT -117.965 10.565 -117.795 11.090 ;
        RECT -111.585 10.565 -111.415 11.090 ;
        RECT -109.960 10.675 -109.500 10.845 ;
        RECT -117.965 10.235 -117.415 10.565 ;
        RECT -111.965 10.235 -111.415 10.565 ;
        RECT -117.965 9.710 -117.795 10.235 ;
        RECT -111.585 9.710 -111.415 10.235 ;
        RECT -109.875 9.950 -109.585 10.675 ;
        RECT -108.045 10.565 -107.875 11.090 ;
        RECT -101.665 10.565 -101.495 11.090 ;
        RECT -100.040 10.675 -99.580 10.845 ;
        RECT -108.045 10.235 -107.495 10.565 ;
        RECT -102.045 10.235 -101.495 10.565 ;
        RECT -108.045 9.710 -107.875 10.235 ;
        RECT -101.665 9.710 -101.495 10.235 ;
        RECT -99.955 9.950 -99.665 10.675 ;
        RECT -98.125 10.565 -97.955 11.090 ;
        RECT -91.745 10.565 -91.575 11.090 ;
        RECT -90.120 10.675 -89.660 10.845 ;
        RECT -98.125 10.235 -97.575 10.565 ;
        RECT -92.125 10.235 -91.575 10.565 ;
        RECT -98.125 9.710 -97.955 10.235 ;
        RECT -91.745 9.710 -91.575 10.235 ;
        RECT -90.035 9.950 -89.745 10.675 ;
        RECT -88.205 10.565 -88.035 11.090 ;
        RECT -81.825 10.565 -81.655 11.090 ;
        RECT -80.200 10.675 -79.740 10.845 ;
        RECT -88.205 10.235 -87.655 10.565 ;
        RECT -82.205 10.235 -81.655 10.565 ;
        RECT -88.205 9.710 -88.035 10.235 ;
        RECT -81.825 9.710 -81.655 10.235 ;
        RECT -80.115 9.950 -79.825 10.675 ;
        RECT -78.285 10.565 -78.115 11.090 ;
        RECT -71.905 10.565 -71.735 11.090 ;
        RECT -70.280 10.675 -69.820 10.845 ;
        RECT -78.285 10.235 -77.735 10.565 ;
        RECT -72.285 10.235 -71.735 10.565 ;
        RECT -78.285 9.710 -78.115 10.235 ;
        RECT -71.905 9.710 -71.735 10.235 ;
        RECT -70.195 9.950 -69.905 10.675 ;
        RECT -68.365 10.565 -68.195 11.090 ;
        RECT -61.985 10.565 -61.815 11.090 ;
        RECT -60.360 10.675 -59.900 10.845 ;
        RECT -68.365 10.235 -67.815 10.565 ;
        RECT -62.365 10.235 -61.815 10.565 ;
        RECT -68.365 9.710 -68.195 10.235 ;
        RECT -61.985 9.710 -61.815 10.235 ;
        RECT -60.275 9.950 -59.985 10.675 ;
        RECT -58.445 10.565 -58.275 11.090 ;
        RECT -52.065 10.565 -51.895 11.090 ;
        RECT -50.440 10.675 -49.980 10.845 ;
        RECT -58.445 10.235 -57.895 10.565 ;
        RECT -52.445 10.235 -51.895 10.565 ;
        RECT -58.445 9.710 -58.275 10.235 ;
        RECT -52.065 9.710 -51.895 10.235 ;
        RECT -50.355 9.950 -50.065 10.675 ;
        RECT -48.525 10.565 -48.355 11.090 ;
        RECT -42.145 10.565 -41.975 11.090 ;
        RECT -40.520 10.675 -40.060 10.845 ;
        RECT -48.525 10.235 -47.975 10.565 ;
        RECT -42.525 10.235 -41.975 10.565 ;
        RECT -48.525 9.710 -48.355 10.235 ;
        RECT -42.145 9.710 -41.975 10.235 ;
        RECT -40.435 9.950 -40.145 10.675 ;
        RECT -38.605 10.565 -38.435 11.090 ;
        RECT -32.225 10.565 -32.055 11.090 ;
        RECT -30.600 10.675 -30.140 10.845 ;
        RECT -38.605 10.235 -38.055 10.565 ;
        RECT -32.605 10.235 -32.055 10.565 ;
        RECT -38.605 9.710 -38.435 10.235 ;
        RECT -32.225 9.710 -32.055 10.235 ;
        RECT -30.515 9.950 -30.225 10.675 ;
        RECT -28.685 10.565 -28.515 11.090 ;
        RECT -22.305 10.565 -22.135 11.090 ;
        RECT -20.680 10.675 -20.220 10.845 ;
        RECT -28.685 10.235 -28.135 10.565 ;
        RECT -22.685 10.235 -22.135 10.565 ;
        RECT -28.685 9.710 -28.515 10.235 ;
        RECT -22.305 9.710 -22.135 10.235 ;
        RECT -20.595 9.950 -20.305 10.675 ;
        RECT -18.765 10.565 -18.595 11.090 ;
        RECT -12.385 10.565 -12.215 11.090 ;
        RECT -10.760 10.675 -10.300 10.845 ;
        RECT -18.765 10.235 -18.215 10.565 ;
        RECT -12.765 10.235 -12.215 10.565 ;
        RECT -18.765 9.710 -18.595 10.235 ;
        RECT -12.385 9.710 -12.215 10.235 ;
        RECT -10.675 9.950 -10.385 10.675 ;
        RECT -8.845 10.565 -8.675 11.090 ;
        RECT -2.465 10.565 -2.295 11.090 ;
        RECT -0.840 10.675 -0.380 10.845 ;
        RECT -8.845 10.235 -8.295 10.565 ;
        RECT -2.845 10.235 -2.295 10.565 ;
        RECT -8.845 9.710 -8.675 10.235 ;
        RECT -2.465 9.710 -2.295 10.235 ;
        RECT -0.755 9.950 -0.465 10.675 ;
        RECT 1.075 10.565 1.245 11.090 ;
        RECT 7.455 10.565 7.625 11.090 ;
        RECT 9.080 10.675 9.540 10.845 ;
        RECT 1.075 10.235 1.625 10.565 ;
        RECT 7.075 10.235 7.625 10.565 ;
        RECT 1.075 9.710 1.245 10.235 ;
        RECT 7.455 9.710 7.625 10.235 ;
        RECT 9.165 9.950 9.455 10.675 ;
        RECT 10.995 10.565 11.165 11.090 ;
        RECT 17.375 10.565 17.545 11.090 ;
        RECT 19.000 10.675 19.460 10.845 ;
        RECT 10.995 10.235 11.545 10.565 ;
        RECT 16.995 10.235 17.545 10.565 ;
        RECT 10.995 9.710 11.165 10.235 ;
        RECT 17.375 9.710 17.545 10.235 ;
        RECT 19.085 9.950 19.375 10.675 ;
        RECT 20.915 10.565 21.085 11.090 ;
        RECT 20.915 10.235 21.465 10.565 ;
        RECT 20.915 9.710 21.085 10.235 ;
        RECT -284.940 9.195 -281.720 9.365 ;
        RECT -275.020 9.195 -271.800 9.365 ;
        RECT -265.100 9.195 -261.880 9.365 ;
        RECT -255.180 9.195 -251.960 9.365 ;
        RECT -245.260 9.195 -242.040 9.365 ;
        RECT -235.340 9.195 -232.120 9.365 ;
        RECT -225.420 9.195 -222.200 9.365 ;
        RECT -215.500 9.195 -212.280 9.365 ;
        RECT -205.580 9.195 -202.360 9.365 ;
        RECT -195.660 9.195 -192.440 9.365 ;
        RECT -185.740 9.195 -182.520 9.365 ;
        RECT -175.820 9.195 -172.600 9.365 ;
        RECT -165.900 9.195 -162.680 9.365 ;
        RECT -155.980 9.195 -152.760 9.365 ;
        RECT -146.060 9.195 -142.840 9.365 ;
        RECT -136.140 9.195 -132.920 9.365 ;
        RECT -126.220 9.195 -123.000 9.365 ;
        RECT -116.300 9.195 -113.080 9.365 ;
        RECT -106.380 9.195 -103.160 9.365 ;
        RECT -96.460 9.195 -93.240 9.365 ;
        RECT -86.540 9.195 -83.320 9.365 ;
        RECT -76.620 9.195 -73.400 9.365 ;
        RECT -66.700 9.195 -63.480 9.365 ;
        RECT -56.780 9.195 -53.560 9.365 ;
        RECT -46.860 9.195 -43.640 9.365 ;
        RECT -36.940 9.195 -33.720 9.365 ;
        RECT -27.020 9.195 -23.800 9.365 ;
        RECT -17.100 9.195 -13.880 9.365 ;
        RECT -7.180 9.195 -3.960 9.365 ;
        RECT 2.740 9.195 5.960 9.365 ;
        RECT 12.660 9.195 15.880 9.365 ;
        RECT -283.955 8.395 -283.645 9.195 ;
        RECT -283.475 8.470 -283.185 9.195 ;
        RECT -283.015 8.395 -282.705 9.195 ;
        RECT -274.035 8.395 -273.725 9.195 ;
        RECT -273.555 8.470 -273.265 9.195 ;
        RECT -273.095 8.395 -272.785 9.195 ;
        RECT -264.115 8.395 -263.805 9.195 ;
        RECT -263.635 8.470 -263.345 9.195 ;
        RECT -263.175 8.395 -262.865 9.195 ;
        RECT -254.195 8.395 -253.885 9.195 ;
        RECT -253.715 8.470 -253.425 9.195 ;
        RECT -253.255 8.395 -252.945 9.195 ;
        RECT -244.275 8.395 -243.965 9.195 ;
        RECT -243.795 8.470 -243.505 9.195 ;
        RECT -243.335 8.395 -243.025 9.195 ;
        RECT -234.355 8.395 -234.045 9.195 ;
        RECT -233.875 8.470 -233.585 9.195 ;
        RECT -233.415 8.395 -233.105 9.195 ;
        RECT -224.435 8.395 -224.125 9.195 ;
        RECT -223.955 8.470 -223.665 9.195 ;
        RECT -223.495 8.395 -223.185 9.195 ;
        RECT -214.515 8.395 -214.205 9.195 ;
        RECT -214.035 8.470 -213.745 9.195 ;
        RECT -213.575 8.395 -213.265 9.195 ;
        RECT -204.595 8.395 -204.285 9.195 ;
        RECT -204.115 8.470 -203.825 9.195 ;
        RECT -203.655 8.395 -203.345 9.195 ;
        RECT -194.675 8.395 -194.365 9.195 ;
        RECT -194.195 8.470 -193.905 9.195 ;
        RECT -193.735 8.395 -193.425 9.195 ;
        RECT -184.755 8.395 -184.445 9.195 ;
        RECT -184.275 8.470 -183.985 9.195 ;
        RECT -183.815 8.395 -183.505 9.195 ;
        RECT -174.835 8.395 -174.525 9.195 ;
        RECT -174.355 8.470 -174.065 9.195 ;
        RECT -173.895 8.395 -173.585 9.195 ;
        RECT -164.915 8.395 -164.605 9.195 ;
        RECT -164.435 8.470 -164.145 9.195 ;
        RECT -163.975 8.395 -163.665 9.195 ;
        RECT -154.995 8.395 -154.685 9.195 ;
        RECT -154.515 8.470 -154.225 9.195 ;
        RECT -154.055 8.395 -153.745 9.195 ;
        RECT -145.075 8.395 -144.765 9.195 ;
        RECT -144.595 8.470 -144.305 9.195 ;
        RECT -144.135 8.395 -143.825 9.195 ;
        RECT -135.155 8.395 -134.845 9.195 ;
        RECT -134.675 8.470 -134.385 9.195 ;
        RECT -134.215 8.395 -133.905 9.195 ;
        RECT -125.235 8.395 -124.925 9.195 ;
        RECT -124.755 8.470 -124.465 9.195 ;
        RECT -124.295 8.395 -123.985 9.195 ;
        RECT -115.315 8.395 -115.005 9.195 ;
        RECT -114.835 8.470 -114.545 9.195 ;
        RECT -114.375 8.395 -114.065 9.195 ;
        RECT -105.395 8.395 -105.085 9.195 ;
        RECT -104.915 8.470 -104.625 9.195 ;
        RECT -104.455 8.395 -104.145 9.195 ;
        RECT -95.475 8.395 -95.165 9.195 ;
        RECT -94.995 8.470 -94.705 9.195 ;
        RECT -94.535 8.395 -94.225 9.195 ;
        RECT -85.555 8.395 -85.245 9.195 ;
        RECT -85.075 8.470 -84.785 9.195 ;
        RECT -84.615 8.395 -84.305 9.195 ;
        RECT -75.635 8.395 -75.325 9.195 ;
        RECT -75.155 8.470 -74.865 9.195 ;
        RECT -74.695 8.395 -74.385 9.195 ;
        RECT -65.715 8.395 -65.405 9.195 ;
        RECT -65.235 8.470 -64.945 9.195 ;
        RECT -64.775 8.395 -64.465 9.195 ;
        RECT -55.795 8.395 -55.485 9.195 ;
        RECT -55.315 8.470 -55.025 9.195 ;
        RECT -54.855 8.395 -54.545 9.195 ;
        RECT -45.875 8.395 -45.565 9.195 ;
        RECT -45.395 8.470 -45.105 9.195 ;
        RECT -44.935 8.395 -44.625 9.195 ;
        RECT -35.955 8.395 -35.645 9.195 ;
        RECT -35.475 8.470 -35.185 9.195 ;
        RECT -35.015 8.395 -34.705 9.195 ;
        RECT -26.035 8.395 -25.725 9.195 ;
        RECT -25.555 8.470 -25.265 9.195 ;
        RECT -25.095 8.395 -24.785 9.195 ;
        RECT -16.115 8.395 -15.805 9.195 ;
        RECT -15.635 8.470 -15.345 9.195 ;
        RECT -15.175 8.395 -14.865 9.195 ;
        RECT -6.195 8.395 -5.885 9.195 ;
        RECT -5.715 8.470 -5.425 9.195 ;
        RECT -5.255 8.395 -4.945 9.195 ;
        RECT 3.725 8.395 4.035 9.195 ;
        RECT 4.205 8.470 4.495 9.195 ;
        RECT 4.665 8.395 4.975 9.195 ;
        RECT 13.645 8.395 13.955 9.195 ;
        RECT 14.125 8.470 14.415 9.195 ;
        RECT 14.585 8.395 14.895 9.195 ;
        RECT -288.915 6.645 -288.605 7.445 ;
        RECT -288.435 6.645 -288.145 7.370 ;
        RECT -287.975 6.645 -287.665 7.445 ;
        RECT -278.995 6.645 -278.685 7.445 ;
        RECT -278.515 6.645 -278.225 7.370 ;
        RECT -278.055 6.645 -277.745 7.445 ;
        RECT -269.075 6.645 -268.765 7.445 ;
        RECT -268.595 6.645 -268.305 7.370 ;
        RECT -268.135 6.645 -267.825 7.445 ;
        RECT -259.155 6.645 -258.845 7.445 ;
        RECT -258.675 6.645 -258.385 7.370 ;
        RECT -258.215 6.645 -257.905 7.445 ;
        RECT -249.235 6.645 -248.925 7.445 ;
        RECT -248.755 6.645 -248.465 7.370 ;
        RECT -248.295 6.645 -247.985 7.445 ;
        RECT -239.315 6.645 -239.005 7.445 ;
        RECT -238.835 6.645 -238.545 7.370 ;
        RECT -238.375 6.645 -238.065 7.445 ;
        RECT -229.395 6.645 -229.085 7.445 ;
        RECT -228.915 6.645 -228.625 7.370 ;
        RECT -228.455 6.645 -228.145 7.445 ;
        RECT -219.475 6.645 -219.165 7.445 ;
        RECT -218.995 6.645 -218.705 7.370 ;
        RECT -218.535 6.645 -218.225 7.445 ;
        RECT -209.555 6.645 -209.245 7.445 ;
        RECT -209.075 6.645 -208.785 7.370 ;
        RECT -208.615 6.645 -208.305 7.445 ;
        RECT -199.635 6.645 -199.325 7.445 ;
        RECT -199.155 6.645 -198.865 7.370 ;
        RECT -198.695 6.645 -198.385 7.445 ;
        RECT -189.715 6.645 -189.405 7.445 ;
        RECT -189.235 6.645 -188.945 7.370 ;
        RECT -188.775 6.645 -188.465 7.445 ;
        RECT -179.795 6.645 -179.485 7.445 ;
        RECT -179.315 6.645 -179.025 7.370 ;
        RECT -178.855 6.645 -178.545 7.445 ;
        RECT -169.875 6.645 -169.565 7.445 ;
        RECT -169.395 6.645 -169.105 7.370 ;
        RECT -168.935 6.645 -168.625 7.445 ;
        RECT -159.955 6.645 -159.645 7.445 ;
        RECT -159.475 6.645 -159.185 7.370 ;
        RECT -159.015 6.645 -158.705 7.445 ;
        RECT -150.035 6.645 -149.725 7.445 ;
        RECT -149.555 6.645 -149.265 7.370 ;
        RECT -149.095 6.645 -148.785 7.445 ;
        RECT -140.115 6.645 -139.805 7.445 ;
        RECT -139.635 6.645 -139.345 7.370 ;
        RECT -139.175 6.645 -138.865 7.445 ;
        RECT -130.195 6.645 -129.885 7.445 ;
        RECT -129.715 6.645 -129.425 7.370 ;
        RECT -129.255 6.645 -128.945 7.445 ;
        RECT -120.275 6.645 -119.965 7.445 ;
        RECT -119.795 6.645 -119.505 7.370 ;
        RECT -119.335 6.645 -119.025 7.445 ;
        RECT -110.355 6.645 -110.045 7.445 ;
        RECT -109.875 6.645 -109.585 7.370 ;
        RECT -109.415 6.645 -109.105 7.445 ;
        RECT -100.435 6.645 -100.125 7.445 ;
        RECT -99.955 6.645 -99.665 7.370 ;
        RECT -99.495 6.645 -99.185 7.445 ;
        RECT -90.515 6.645 -90.205 7.445 ;
        RECT -90.035 6.645 -89.745 7.370 ;
        RECT -89.575 6.645 -89.265 7.445 ;
        RECT -80.595 6.645 -80.285 7.445 ;
        RECT -80.115 6.645 -79.825 7.370 ;
        RECT -79.655 6.645 -79.345 7.445 ;
        RECT -70.675 6.645 -70.365 7.445 ;
        RECT -70.195 6.645 -69.905 7.370 ;
        RECT -69.735 6.645 -69.425 7.445 ;
        RECT -60.755 6.645 -60.445 7.445 ;
        RECT -60.275 6.645 -59.985 7.370 ;
        RECT -59.815 6.645 -59.505 7.445 ;
        RECT -50.835 6.645 -50.525 7.445 ;
        RECT -50.355 6.645 -50.065 7.370 ;
        RECT -49.895 6.645 -49.585 7.445 ;
        RECT -40.915 6.645 -40.605 7.445 ;
        RECT -40.435 6.645 -40.145 7.370 ;
        RECT -39.975 6.645 -39.665 7.445 ;
        RECT -30.995 6.645 -30.685 7.445 ;
        RECT -30.515 6.645 -30.225 7.370 ;
        RECT -30.055 6.645 -29.745 7.445 ;
        RECT -21.075 6.645 -20.765 7.445 ;
        RECT -20.595 6.645 -20.305 7.370 ;
        RECT -20.135 6.645 -19.825 7.445 ;
        RECT -11.155 6.645 -10.845 7.445 ;
        RECT -10.675 6.645 -10.385 7.370 ;
        RECT -10.215 6.645 -9.905 7.445 ;
        RECT -1.235 6.645 -0.925 7.445 ;
        RECT -0.755 6.645 -0.465 7.370 ;
        RECT -0.295 6.645 0.015 7.445 ;
        RECT 8.685 6.645 8.995 7.445 ;
        RECT 9.165 6.645 9.455 7.370 ;
        RECT 9.625 6.645 9.935 7.445 ;
        RECT 18.605 6.645 18.915 7.445 ;
        RECT 19.085 6.645 19.375 7.370 ;
        RECT 19.545 6.645 19.855 7.445 ;
        RECT -289.900 6.475 -286.680 6.645 ;
        RECT -279.980 6.475 -276.760 6.645 ;
        RECT -270.060 6.475 -266.840 6.645 ;
        RECT -260.140 6.475 -256.920 6.645 ;
        RECT -250.220 6.475 -247.000 6.645 ;
        RECT -240.300 6.475 -237.080 6.645 ;
        RECT -230.380 6.475 -227.160 6.645 ;
        RECT -220.460 6.475 -217.240 6.645 ;
        RECT -210.540 6.475 -207.320 6.645 ;
        RECT -200.620 6.475 -197.400 6.645 ;
        RECT -190.700 6.475 -187.480 6.645 ;
        RECT -180.780 6.475 -177.560 6.645 ;
        RECT -170.860 6.475 -167.640 6.645 ;
        RECT -160.940 6.475 -157.720 6.645 ;
        RECT -151.020 6.475 -147.800 6.645 ;
        RECT -141.100 6.475 -137.880 6.645 ;
        RECT -131.180 6.475 -127.960 6.645 ;
        RECT -121.260 6.475 -118.040 6.645 ;
        RECT -111.340 6.475 -108.120 6.645 ;
        RECT -101.420 6.475 -98.200 6.645 ;
        RECT -91.500 6.475 -88.280 6.645 ;
        RECT -81.580 6.475 -78.360 6.645 ;
        RECT -71.660 6.475 -68.440 6.645 ;
        RECT -61.740 6.475 -58.520 6.645 ;
        RECT -51.820 6.475 -48.600 6.645 ;
        RECT -41.900 6.475 -38.680 6.645 ;
        RECT -31.980 6.475 -28.760 6.645 ;
        RECT -22.060 6.475 -18.840 6.645 ;
        RECT -12.140 6.475 -8.920 6.645 ;
        RECT -2.220 6.475 1.000 6.645 ;
        RECT 7.700 6.475 10.920 6.645 ;
        RECT 17.620 6.475 20.840 6.645 ;
        RECT -285.185 5.605 -285.015 6.130 ;
        RECT -285.565 5.275 -285.015 5.605 ;
        RECT -285.185 4.750 -285.015 5.275 ;
        RECT -283.475 5.255 -283.185 5.980 ;
        RECT -281.645 5.605 -281.475 6.130 ;
        RECT -275.265 5.605 -275.095 6.130 ;
        RECT -281.645 5.275 -281.095 5.605 ;
        RECT -275.645 5.275 -275.095 5.605 ;
        RECT -283.560 5.085 -283.100 5.255 ;
        RECT -281.645 4.750 -281.475 5.275 ;
        RECT -275.265 4.750 -275.095 5.275 ;
        RECT -273.555 5.255 -273.265 5.980 ;
        RECT -271.725 5.605 -271.555 6.130 ;
        RECT -265.345 5.605 -265.175 6.130 ;
        RECT -271.725 5.275 -271.175 5.605 ;
        RECT -265.725 5.275 -265.175 5.605 ;
        RECT -273.640 5.085 -273.180 5.255 ;
        RECT -271.725 4.750 -271.555 5.275 ;
        RECT -265.345 4.750 -265.175 5.275 ;
        RECT -263.635 5.255 -263.345 5.980 ;
        RECT -261.805 5.605 -261.635 6.130 ;
        RECT -255.425 5.605 -255.255 6.130 ;
        RECT -261.805 5.275 -261.255 5.605 ;
        RECT -255.805 5.275 -255.255 5.605 ;
        RECT -263.720 5.085 -263.260 5.255 ;
        RECT -261.805 4.750 -261.635 5.275 ;
        RECT -255.425 4.750 -255.255 5.275 ;
        RECT -253.715 5.255 -253.425 5.980 ;
        RECT -251.885 5.605 -251.715 6.130 ;
        RECT -245.505 5.605 -245.335 6.130 ;
        RECT -251.885 5.275 -251.335 5.605 ;
        RECT -245.885 5.275 -245.335 5.605 ;
        RECT -253.800 5.085 -253.340 5.255 ;
        RECT -251.885 4.750 -251.715 5.275 ;
        RECT -245.505 4.750 -245.335 5.275 ;
        RECT -243.795 5.255 -243.505 5.980 ;
        RECT -241.965 5.605 -241.795 6.130 ;
        RECT -235.585 5.605 -235.415 6.130 ;
        RECT -241.965 5.275 -241.415 5.605 ;
        RECT -235.965 5.275 -235.415 5.605 ;
        RECT -243.880 5.085 -243.420 5.255 ;
        RECT -241.965 4.750 -241.795 5.275 ;
        RECT -235.585 4.750 -235.415 5.275 ;
        RECT -233.875 5.255 -233.585 5.980 ;
        RECT -232.045 5.605 -231.875 6.130 ;
        RECT -225.665 5.605 -225.495 6.130 ;
        RECT -232.045 5.275 -231.495 5.605 ;
        RECT -226.045 5.275 -225.495 5.605 ;
        RECT -233.960 5.085 -233.500 5.255 ;
        RECT -232.045 4.750 -231.875 5.275 ;
        RECT -225.665 4.750 -225.495 5.275 ;
        RECT -223.955 5.255 -223.665 5.980 ;
        RECT -222.125 5.605 -221.955 6.130 ;
        RECT -215.745 5.605 -215.575 6.130 ;
        RECT -222.125 5.275 -221.575 5.605 ;
        RECT -216.125 5.275 -215.575 5.605 ;
        RECT -224.040 5.085 -223.580 5.255 ;
        RECT -222.125 4.750 -221.955 5.275 ;
        RECT -215.745 4.750 -215.575 5.275 ;
        RECT -214.035 5.255 -213.745 5.980 ;
        RECT -212.205 5.605 -212.035 6.130 ;
        RECT -205.825 5.605 -205.655 6.130 ;
        RECT -212.205 5.275 -211.655 5.605 ;
        RECT -206.205 5.275 -205.655 5.605 ;
        RECT -214.120 5.085 -213.660 5.255 ;
        RECT -212.205 4.750 -212.035 5.275 ;
        RECT -205.825 4.750 -205.655 5.275 ;
        RECT -204.115 5.255 -203.825 5.980 ;
        RECT -202.285 5.605 -202.115 6.130 ;
        RECT -195.905 5.605 -195.735 6.130 ;
        RECT -202.285 5.275 -201.735 5.605 ;
        RECT -196.285 5.275 -195.735 5.605 ;
        RECT -204.200 5.085 -203.740 5.255 ;
        RECT -202.285 4.750 -202.115 5.275 ;
        RECT -195.905 4.750 -195.735 5.275 ;
        RECT -194.195 5.255 -193.905 5.980 ;
        RECT -192.365 5.605 -192.195 6.130 ;
        RECT -185.985 5.605 -185.815 6.130 ;
        RECT -192.365 5.275 -191.815 5.605 ;
        RECT -186.365 5.275 -185.815 5.605 ;
        RECT -194.280 5.085 -193.820 5.255 ;
        RECT -192.365 4.750 -192.195 5.275 ;
        RECT -185.985 4.750 -185.815 5.275 ;
        RECT -184.275 5.255 -183.985 5.980 ;
        RECT -182.445 5.605 -182.275 6.130 ;
        RECT -176.065 5.605 -175.895 6.130 ;
        RECT -182.445 5.275 -181.895 5.605 ;
        RECT -176.445 5.275 -175.895 5.605 ;
        RECT -184.360 5.085 -183.900 5.255 ;
        RECT -182.445 4.750 -182.275 5.275 ;
        RECT -176.065 4.750 -175.895 5.275 ;
        RECT -174.355 5.255 -174.065 5.980 ;
        RECT -172.525 5.605 -172.355 6.130 ;
        RECT -166.145 5.605 -165.975 6.130 ;
        RECT -172.525 5.275 -171.975 5.605 ;
        RECT -166.525 5.275 -165.975 5.605 ;
        RECT -174.440 5.085 -173.980 5.255 ;
        RECT -172.525 4.750 -172.355 5.275 ;
        RECT -166.145 4.750 -165.975 5.275 ;
        RECT -164.435 5.255 -164.145 5.980 ;
        RECT -162.605 5.605 -162.435 6.130 ;
        RECT -156.225 5.605 -156.055 6.130 ;
        RECT -162.605 5.275 -162.055 5.605 ;
        RECT -156.605 5.275 -156.055 5.605 ;
        RECT -164.520 5.085 -164.060 5.255 ;
        RECT -162.605 4.750 -162.435 5.275 ;
        RECT -156.225 4.750 -156.055 5.275 ;
        RECT -154.515 5.255 -154.225 5.980 ;
        RECT -152.685 5.605 -152.515 6.130 ;
        RECT -146.305 5.605 -146.135 6.130 ;
        RECT -152.685 5.275 -152.135 5.605 ;
        RECT -146.685 5.275 -146.135 5.605 ;
        RECT -154.600 5.085 -154.140 5.255 ;
        RECT -152.685 4.750 -152.515 5.275 ;
        RECT -146.305 4.750 -146.135 5.275 ;
        RECT -144.595 5.255 -144.305 5.980 ;
        RECT -142.765 5.605 -142.595 6.130 ;
        RECT -136.385 5.605 -136.215 6.130 ;
        RECT -142.765 5.275 -142.215 5.605 ;
        RECT -136.765 5.275 -136.215 5.605 ;
        RECT -144.680 5.085 -144.220 5.255 ;
        RECT -142.765 4.750 -142.595 5.275 ;
        RECT -136.385 4.750 -136.215 5.275 ;
        RECT -134.675 5.255 -134.385 5.980 ;
        RECT -132.845 5.605 -132.675 6.130 ;
        RECT -126.465 5.605 -126.295 6.130 ;
        RECT -132.845 5.275 -132.295 5.605 ;
        RECT -126.845 5.275 -126.295 5.605 ;
        RECT -134.760 5.085 -134.300 5.255 ;
        RECT -132.845 4.750 -132.675 5.275 ;
        RECT -126.465 4.750 -126.295 5.275 ;
        RECT -124.755 5.255 -124.465 5.980 ;
        RECT -122.925 5.605 -122.755 6.130 ;
        RECT -116.545 5.605 -116.375 6.130 ;
        RECT -122.925 5.275 -122.375 5.605 ;
        RECT -116.925 5.275 -116.375 5.605 ;
        RECT -124.840 5.085 -124.380 5.255 ;
        RECT -122.925 4.750 -122.755 5.275 ;
        RECT -116.545 4.750 -116.375 5.275 ;
        RECT -114.835 5.255 -114.545 5.980 ;
        RECT -113.005 5.605 -112.835 6.130 ;
        RECT -106.625 5.605 -106.455 6.130 ;
        RECT -113.005 5.275 -112.455 5.605 ;
        RECT -107.005 5.275 -106.455 5.605 ;
        RECT -114.920 5.085 -114.460 5.255 ;
        RECT -113.005 4.750 -112.835 5.275 ;
        RECT -106.625 4.750 -106.455 5.275 ;
        RECT -104.915 5.255 -104.625 5.980 ;
        RECT -103.085 5.605 -102.915 6.130 ;
        RECT -96.705 5.605 -96.535 6.130 ;
        RECT -103.085 5.275 -102.535 5.605 ;
        RECT -97.085 5.275 -96.535 5.605 ;
        RECT -105.000 5.085 -104.540 5.255 ;
        RECT -103.085 4.750 -102.915 5.275 ;
        RECT -96.705 4.750 -96.535 5.275 ;
        RECT -94.995 5.255 -94.705 5.980 ;
        RECT -93.165 5.605 -92.995 6.130 ;
        RECT -86.785 5.605 -86.615 6.130 ;
        RECT -93.165 5.275 -92.615 5.605 ;
        RECT -87.165 5.275 -86.615 5.605 ;
        RECT -95.080 5.085 -94.620 5.255 ;
        RECT -93.165 4.750 -92.995 5.275 ;
        RECT -86.785 4.750 -86.615 5.275 ;
        RECT -85.075 5.255 -84.785 5.980 ;
        RECT -83.245 5.605 -83.075 6.130 ;
        RECT -76.865 5.605 -76.695 6.130 ;
        RECT -83.245 5.275 -82.695 5.605 ;
        RECT -77.245 5.275 -76.695 5.605 ;
        RECT -85.160 5.085 -84.700 5.255 ;
        RECT -83.245 4.750 -83.075 5.275 ;
        RECT -76.865 4.750 -76.695 5.275 ;
        RECT -75.155 5.255 -74.865 5.980 ;
        RECT -73.325 5.605 -73.155 6.130 ;
        RECT -66.945 5.605 -66.775 6.130 ;
        RECT -73.325 5.275 -72.775 5.605 ;
        RECT -67.325 5.275 -66.775 5.605 ;
        RECT -75.240 5.085 -74.780 5.255 ;
        RECT -73.325 4.750 -73.155 5.275 ;
        RECT -66.945 4.750 -66.775 5.275 ;
        RECT -65.235 5.255 -64.945 5.980 ;
        RECT -63.405 5.605 -63.235 6.130 ;
        RECT -57.025 5.605 -56.855 6.130 ;
        RECT -63.405 5.275 -62.855 5.605 ;
        RECT -57.405 5.275 -56.855 5.605 ;
        RECT -65.320 5.085 -64.860 5.255 ;
        RECT -63.405 4.750 -63.235 5.275 ;
        RECT -57.025 4.750 -56.855 5.275 ;
        RECT -55.315 5.255 -55.025 5.980 ;
        RECT -53.485 5.605 -53.315 6.130 ;
        RECT -47.105 5.605 -46.935 6.130 ;
        RECT -53.485 5.275 -52.935 5.605 ;
        RECT -47.485 5.275 -46.935 5.605 ;
        RECT -55.400 5.085 -54.940 5.255 ;
        RECT -53.485 4.750 -53.315 5.275 ;
        RECT -47.105 4.750 -46.935 5.275 ;
        RECT -45.395 5.255 -45.105 5.980 ;
        RECT -43.565 5.605 -43.395 6.130 ;
        RECT -37.185 5.605 -37.015 6.130 ;
        RECT -43.565 5.275 -43.015 5.605 ;
        RECT -37.565 5.275 -37.015 5.605 ;
        RECT -45.480 5.085 -45.020 5.255 ;
        RECT -43.565 4.750 -43.395 5.275 ;
        RECT -37.185 4.750 -37.015 5.275 ;
        RECT -35.475 5.255 -35.185 5.980 ;
        RECT -33.645 5.605 -33.475 6.130 ;
        RECT -27.265 5.605 -27.095 6.130 ;
        RECT -33.645 5.275 -33.095 5.605 ;
        RECT -27.645 5.275 -27.095 5.605 ;
        RECT -35.560 5.085 -35.100 5.255 ;
        RECT -33.645 4.750 -33.475 5.275 ;
        RECT -27.265 4.750 -27.095 5.275 ;
        RECT -25.555 5.255 -25.265 5.980 ;
        RECT -23.725 5.605 -23.555 6.130 ;
        RECT -17.345 5.605 -17.175 6.130 ;
        RECT -23.725 5.275 -23.175 5.605 ;
        RECT -17.725 5.275 -17.175 5.605 ;
        RECT -25.640 5.085 -25.180 5.255 ;
        RECT -23.725 4.750 -23.555 5.275 ;
        RECT -17.345 4.750 -17.175 5.275 ;
        RECT -15.635 5.255 -15.345 5.980 ;
        RECT -13.805 5.605 -13.635 6.130 ;
        RECT -7.425 5.605 -7.255 6.130 ;
        RECT -13.805 5.275 -13.255 5.605 ;
        RECT -7.805 5.275 -7.255 5.605 ;
        RECT -15.720 5.085 -15.260 5.255 ;
        RECT -13.805 4.750 -13.635 5.275 ;
        RECT -7.425 4.750 -7.255 5.275 ;
        RECT -5.715 5.255 -5.425 5.980 ;
        RECT -3.885 5.605 -3.715 6.130 ;
        RECT 2.495 5.605 2.665 6.130 ;
        RECT -3.885 5.275 -3.335 5.605 ;
        RECT 2.115 5.275 2.665 5.605 ;
        RECT -5.800 5.085 -5.340 5.255 ;
        RECT -3.885 4.750 -3.715 5.275 ;
        RECT 2.495 4.750 2.665 5.275 ;
        RECT 4.205 5.255 4.495 5.980 ;
        RECT 6.035 5.605 6.205 6.130 ;
        RECT 12.415 5.605 12.585 6.130 ;
        RECT 6.035 5.275 6.585 5.605 ;
        RECT 12.035 5.275 12.585 5.605 ;
        RECT 4.120 5.085 4.580 5.255 ;
        RECT 6.035 4.750 6.205 5.275 ;
        RECT 12.415 4.750 12.585 5.275 ;
        RECT 14.125 5.255 14.415 5.980 ;
        RECT 15.955 5.605 16.125 6.130 ;
        RECT 15.955 5.275 16.505 5.605 ;
        RECT 14.040 5.085 14.500 5.255 ;
        RECT 15.955 4.750 16.125 5.275 ;
        RECT -289.785 -78.385 -289.615 -77.860 ;
        RECT -288.160 -78.275 -287.700 -78.105 ;
        RECT -290.165 -78.715 -289.615 -78.385 ;
        RECT -289.785 -79.240 -289.615 -78.715 ;
        RECT -288.075 -79.000 -287.785 -78.275 ;
        RECT -286.245 -78.385 -286.075 -77.860 ;
        RECT -279.865 -78.385 -279.695 -77.860 ;
        RECT -278.240 -78.275 -277.780 -78.105 ;
        RECT -286.245 -78.715 -285.695 -78.385 ;
        RECT -280.245 -78.715 -279.695 -78.385 ;
        RECT -286.245 -79.240 -286.075 -78.715 ;
        RECT -279.865 -79.240 -279.695 -78.715 ;
        RECT -278.155 -79.000 -277.865 -78.275 ;
        RECT -276.325 -78.385 -276.155 -77.860 ;
        RECT -269.945 -78.385 -269.775 -77.860 ;
        RECT -268.320 -78.275 -267.860 -78.105 ;
        RECT -276.325 -78.715 -275.775 -78.385 ;
        RECT -270.325 -78.715 -269.775 -78.385 ;
        RECT -276.325 -79.240 -276.155 -78.715 ;
        RECT -269.945 -79.240 -269.775 -78.715 ;
        RECT -268.235 -79.000 -267.945 -78.275 ;
        RECT -266.405 -78.385 -266.235 -77.860 ;
        RECT -260.025 -78.385 -259.855 -77.860 ;
        RECT -258.400 -78.275 -257.940 -78.105 ;
        RECT -266.405 -78.715 -265.855 -78.385 ;
        RECT -260.405 -78.715 -259.855 -78.385 ;
        RECT -266.405 -79.240 -266.235 -78.715 ;
        RECT -260.025 -79.240 -259.855 -78.715 ;
        RECT -258.315 -79.000 -258.025 -78.275 ;
        RECT -256.485 -78.385 -256.315 -77.860 ;
        RECT -250.105 -78.385 -249.935 -77.860 ;
        RECT -248.480 -78.275 -248.020 -78.105 ;
        RECT -256.485 -78.715 -255.935 -78.385 ;
        RECT -250.485 -78.715 -249.935 -78.385 ;
        RECT -256.485 -79.240 -256.315 -78.715 ;
        RECT -250.105 -79.240 -249.935 -78.715 ;
        RECT -248.395 -79.000 -248.105 -78.275 ;
        RECT -246.565 -78.385 -246.395 -77.860 ;
        RECT -240.185 -78.385 -240.015 -77.860 ;
        RECT -238.560 -78.275 -238.100 -78.105 ;
        RECT -246.565 -78.715 -246.015 -78.385 ;
        RECT -240.565 -78.715 -240.015 -78.385 ;
        RECT -246.565 -79.240 -246.395 -78.715 ;
        RECT -240.185 -79.240 -240.015 -78.715 ;
        RECT -238.475 -79.000 -238.185 -78.275 ;
        RECT -236.645 -78.385 -236.475 -77.860 ;
        RECT -230.265 -78.385 -230.095 -77.860 ;
        RECT -228.640 -78.275 -228.180 -78.105 ;
        RECT -236.645 -78.715 -236.095 -78.385 ;
        RECT -230.645 -78.715 -230.095 -78.385 ;
        RECT -236.645 -79.240 -236.475 -78.715 ;
        RECT -230.265 -79.240 -230.095 -78.715 ;
        RECT -228.555 -79.000 -228.265 -78.275 ;
        RECT -226.725 -78.385 -226.555 -77.860 ;
        RECT -220.345 -78.385 -220.175 -77.860 ;
        RECT -218.720 -78.275 -218.260 -78.105 ;
        RECT -226.725 -78.715 -226.175 -78.385 ;
        RECT -220.725 -78.715 -220.175 -78.385 ;
        RECT -226.725 -79.240 -226.555 -78.715 ;
        RECT -220.345 -79.240 -220.175 -78.715 ;
        RECT -218.635 -79.000 -218.345 -78.275 ;
        RECT -216.805 -78.385 -216.635 -77.860 ;
        RECT -210.425 -78.385 -210.255 -77.860 ;
        RECT -208.800 -78.275 -208.340 -78.105 ;
        RECT -216.805 -78.715 -216.255 -78.385 ;
        RECT -210.805 -78.715 -210.255 -78.385 ;
        RECT -216.805 -79.240 -216.635 -78.715 ;
        RECT -210.425 -79.240 -210.255 -78.715 ;
        RECT -208.715 -79.000 -208.425 -78.275 ;
        RECT -206.885 -78.385 -206.715 -77.860 ;
        RECT -200.505 -78.385 -200.335 -77.860 ;
        RECT -198.880 -78.275 -198.420 -78.105 ;
        RECT -206.885 -78.715 -206.335 -78.385 ;
        RECT -200.885 -78.715 -200.335 -78.385 ;
        RECT -206.885 -79.240 -206.715 -78.715 ;
        RECT -200.505 -79.240 -200.335 -78.715 ;
        RECT -198.795 -79.000 -198.505 -78.275 ;
        RECT -196.965 -78.385 -196.795 -77.860 ;
        RECT -190.585 -78.385 -190.415 -77.860 ;
        RECT -188.960 -78.275 -188.500 -78.105 ;
        RECT -196.965 -78.715 -196.415 -78.385 ;
        RECT -190.965 -78.715 -190.415 -78.385 ;
        RECT -196.965 -79.240 -196.795 -78.715 ;
        RECT -190.585 -79.240 -190.415 -78.715 ;
        RECT -188.875 -79.000 -188.585 -78.275 ;
        RECT -187.045 -78.385 -186.875 -77.860 ;
        RECT -180.665 -78.385 -180.495 -77.860 ;
        RECT -179.040 -78.275 -178.580 -78.105 ;
        RECT -187.045 -78.715 -186.495 -78.385 ;
        RECT -181.045 -78.715 -180.495 -78.385 ;
        RECT -187.045 -79.240 -186.875 -78.715 ;
        RECT -180.665 -79.240 -180.495 -78.715 ;
        RECT -178.955 -79.000 -178.665 -78.275 ;
        RECT -177.125 -78.385 -176.955 -77.860 ;
        RECT -170.745 -78.385 -170.575 -77.860 ;
        RECT -169.120 -78.275 -168.660 -78.105 ;
        RECT -177.125 -78.715 -176.575 -78.385 ;
        RECT -171.125 -78.715 -170.575 -78.385 ;
        RECT -177.125 -79.240 -176.955 -78.715 ;
        RECT -170.745 -79.240 -170.575 -78.715 ;
        RECT -169.035 -79.000 -168.745 -78.275 ;
        RECT -167.205 -78.385 -167.035 -77.860 ;
        RECT -160.825 -78.385 -160.655 -77.860 ;
        RECT -159.200 -78.275 -158.740 -78.105 ;
        RECT -167.205 -78.715 -166.655 -78.385 ;
        RECT -161.205 -78.715 -160.655 -78.385 ;
        RECT -167.205 -79.240 -167.035 -78.715 ;
        RECT -160.825 -79.240 -160.655 -78.715 ;
        RECT -159.115 -79.000 -158.825 -78.275 ;
        RECT -157.285 -78.385 -157.115 -77.860 ;
        RECT -150.905 -78.385 -150.735 -77.860 ;
        RECT -149.280 -78.275 -148.820 -78.105 ;
        RECT -157.285 -78.715 -156.735 -78.385 ;
        RECT -151.285 -78.715 -150.735 -78.385 ;
        RECT -157.285 -79.240 -157.115 -78.715 ;
        RECT -150.905 -79.240 -150.735 -78.715 ;
        RECT -149.195 -79.000 -148.905 -78.275 ;
        RECT -147.365 -78.385 -147.195 -77.860 ;
        RECT -140.985 -78.385 -140.815 -77.860 ;
        RECT -139.360 -78.275 -138.900 -78.105 ;
        RECT -147.365 -78.715 -146.815 -78.385 ;
        RECT -141.365 -78.715 -140.815 -78.385 ;
        RECT -147.365 -79.240 -147.195 -78.715 ;
        RECT -140.985 -79.240 -140.815 -78.715 ;
        RECT -139.275 -79.000 -138.985 -78.275 ;
        RECT -137.445 -78.385 -137.275 -77.860 ;
        RECT -131.065 -78.385 -130.895 -77.860 ;
        RECT -129.440 -78.275 -128.980 -78.105 ;
        RECT -137.445 -78.715 -136.895 -78.385 ;
        RECT -131.445 -78.715 -130.895 -78.385 ;
        RECT -137.445 -79.240 -137.275 -78.715 ;
        RECT -131.065 -79.240 -130.895 -78.715 ;
        RECT -129.355 -79.000 -129.065 -78.275 ;
        RECT -127.525 -78.385 -127.355 -77.860 ;
        RECT -121.145 -78.385 -120.975 -77.860 ;
        RECT -119.520 -78.275 -119.060 -78.105 ;
        RECT -127.525 -78.715 -126.975 -78.385 ;
        RECT -121.525 -78.715 -120.975 -78.385 ;
        RECT -127.525 -79.240 -127.355 -78.715 ;
        RECT -121.145 -79.240 -120.975 -78.715 ;
        RECT -119.435 -79.000 -119.145 -78.275 ;
        RECT -117.605 -78.385 -117.435 -77.860 ;
        RECT -111.225 -78.385 -111.055 -77.860 ;
        RECT -109.600 -78.275 -109.140 -78.105 ;
        RECT -117.605 -78.715 -117.055 -78.385 ;
        RECT -111.605 -78.715 -111.055 -78.385 ;
        RECT -117.605 -79.240 -117.435 -78.715 ;
        RECT -111.225 -79.240 -111.055 -78.715 ;
        RECT -109.515 -79.000 -109.225 -78.275 ;
        RECT -107.685 -78.385 -107.515 -77.860 ;
        RECT -101.305 -78.385 -101.135 -77.860 ;
        RECT -99.680 -78.275 -99.220 -78.105 ;
        RECT -107.685 -78.715 -107.135 -78.385 ;
        RECT -101.685 -78.715 -101.135 -78.385 ;
        RECT -107.685 -79.240 -107.515 -78.715 ;
        RECT -101.305 -79.240 -101.135 -78.715 ;
        RECT -99.595 -79.000 -99.305 -78.275 ;
        RECT -97.765 -78.385 -97.595 -77.860 ;
        RECT -91.385 -78.385 -91.215 -77.860 ;
        RECT -89.760 -78.275 -89.300 -78.105 ;
        RECT -97.765 -78.715 -97.215 -78.385 ;
        RECT -91.765 -78.715 -91.215 -78.385 ;
        RECT -97.765 -79.240 -97.595 -78.715 ;
        RECT -91.385 -79.240 -91.215 -78.715 ;
        RECT -89.675 -79.000 -89.385 -78.275 ;
        RECT -87.845 -78.385 -87.675 -77.860 ;
        RECT -81.465 -78.385 -81.295 -77.860 ;
        RECT -79.840 -78.275 -79.380 -78.105 ;
        RECT -87.845 -78.715 -87.295 -78.385 ;
        RECT -81.845 -78.715 -81.295 -78.385 ;
        RECT -87.845 -79.240 -87.675 -78.715 ;
        RECT -81.465 -79.240 -81.295 -78.715 ;
        RECT -79.755 -79.000 -79.465 -78.275 ;
        RECT -77.925 -78.385 -77.755 -77.860 ;
        RECT -71.545 -78.385 -71.375 -77.860 ;
        RECT -69.920 -78.275 -69.460 -78.105 ;
        RECT -77.925 -78.715 -77.375 -78.385 ;
        RECT -71.925 -78.715 -71.375 -78.385 ;
        RECT -77.925 -79.240 -77.755 -78.715 ;
        RECT -71.545 -79.240 -71.375 -78.715 ;
        RECT -69.835 -79.000 -69.545 -78.275 ;
        RECT -68.005 -78.385 -67.835 -77.860 ;
        RECT -61.625 -78.385 -61.455 -77.860 ;
        RECT -60.000 -78.275 -59.540 -78.105 ;
        RECT -68.005 -78.715 -67.455 -78.385 ;
        RECT -62.005 -78.715 -61.455 -78.385 ;
        RECT -68.005 -79.240 -67.835 -78.715 ;
        RECT -61.625 -79.240 -61.455 -78.715 ;
        RECT -59.915 -79.000 -59.625 -78.275 ;
        RECT -58.085 -78.385 -57.915 -77.860 ;
        RECT -51.705 -78.385 -51.535 -77.860 ;
        RECT -50.080 -78.275 -49.620 -78.105 ;
        RECT -58.085 -78.715 -57.535 -78.385 ;
        RECT -52.085 -78.715 -51.535 -78.385 ;
        RECT -58.085 -79.240 -57.915 -78.715 ;
        RECT -51.705 -79.240 -51.535 -78.715 ;
        RECT -49.995 -79.000 -49.705 -78.275 ;
        RECT -48.165 -78.385 -47.995 -77.860 ;
        RECT -41.785 -78.385 -41.615 -77.860 ;
        RECT -40.160 -78.275 -39.700 -78.105 ;
        RECT -48.165 -78.715 -47.615 -78.385 ;
        RECT -42.165 -78.715 -41.615 -78.385 ;
        RECT -48.165 -79.240 -47.995 -78.715 ;
        RECT -41.785 -79.240 -41.615 -78.715 ;
        RECT -40.075 -79.000 -39.785 -78.275 ;
        RECT -38.245 -78.385 -38.075 -77.860 ;
        RECT -31.865 -78.385 -31.695 -77.860 ;
        RECT -30.240 -78.275 -29.780 -78.105 ;
        RECT -38.245 -78.715 -37.695 -78.385 ;
        RECT -32.245 -78.715 -31.695 -78.385 ;
        RECT -38.245 -79.240 -38.075 -78.715 ;
        RECT -31.865 -79.240 -31.695 -78.715 ;
        RECT -30.155 -79.000 -29.865 -78.275 ;
        RECT -28.325 -78.385 -28.155 -77.860 ;
        RECT -21.945 -78.385 -21.775 -77.860 ;
        RECT -20.320 -78.275 -19.860 -78.105 ;
        RECT -28.325 -78.715 -27.775 -78.385 ;
        RECT -22.325 -78.715 -21.775 -78.385 ;
        RECT -28.325 -79.240 -28.155 -78.715 ;
        RECT -21.945 -79.240 -21.775 -78.715 ;
        RECT -20.235 -79.000 -19.945 -78.275 ;
        RECT -18.405 -78.385 -18.235 -77.860 ;
        RECT -12.025 -78.385 -11.855 -77.860 ;
        RECT -10.400 -78.275 -9.940 -78.105 ;
        RECT -18.405 -78.715 -17.855 -78.385 ;
        RECT -12.405 -78.715 -11.855 -78.385 ;
        RECT -18.405 -79.240 -18.235 -78.715 ;
        RECT -12.025 -79.240 -11.855 -78.715 ;
        RECT -10.315 -79.000 -10.025 -78.275 ;
        RECT -8.485 -78.385 -8.315 -77.860 ;
        RECT -2.105 -78.385 -1.935 -77.860 ;
        RECT -0.480 -78.275 -0.020 -78.105 ;
        RECT -8.485 -78.715 -7.935 -78.385 ;
        RECT -2.485 -78.715 -1.935 -78.385 ;
        RECT -8.485 -79.240 -8.315 -78.715 ;
        RECT -2.105 -79.240 -1.935 -78.715 ;
        RECT -0.395 -79.000 -0.105 -78.275 ;
        RECT 1.435 -78.385 1.605 -77.860 ;
        RECT 7.815 -78.385 7.985 -77.860 ;
        RECT 9.440 -78.275 9.900 -78.105 ;
        RECT 1.435 -78.715 1.985 -78.385 ;
        RECT 7.435 -78.715 7.985 -78.385 ;
        RECT 1.435 -79.240 1.605 -78.715 ;
        RECT 7.815 -79.240 7.985 -78.715 ;
        RECT 9.525 -79.000 9.815 -78.275 ;
        RECT 11.355 -78.385 11.525 -77.860 ;
        RECT 17.735 -78.385 17.905 -77.860 ;
        RECT 19.360 -78.275 19.820 -78.105 ;
        RECT 11.355 -78.715 11.905 -78.385 ;
        RECT 17.355 -78.715 17.905 -78.385 ;
        RECT 11.355 -79.240 11.525 -78.715 ;
        RECT 17.735 -79.240 17.905 -78.715 ;
        RECT 19.445 -79.000 19.735 -78.275 ;
        RECT 21.275 -78.385 21.445 -77.860 ;
        RECT 21.275 -78.715 21.825 -78.385 ;
        RECT 21.275 -79.240 21.445 -78.715 ;
        RECT -284.580 -79.755 -281.360 -79.585 ;
        RECT -274.660 -79.755 -271.440 -79.585 ;
        RECT -264.740 -79.755 -261.520 -79.585 ;
        RECT -254.820 -79.755 -251.600 -79.585 ;
        RECT -244.900 -79.755 -241.680 -79.585 ;
        RECT -234.980 -79.755 -231.760 -79.585 ;
        RECT -225.060 -79.755 -221.840 -79.585 ;
        RECT -215.140 -79.755 -211.920 -79.585 ;
        RECT -205.220 -79.755 -202.000 -79.585 ;
        RECT -195.300 -79.755 -192.080 -79.585 ;
        RECT -185.380 -79.755 -182.160 -79.585 ;
        RECT -175.460 -79.755 -172.240 -79.585 ;
        RECT -165.540 -79.755 -162.320 -79.585 ;
        RECT -155.620 -79.755 -152.400 -79.585 ;
        RECT -145.700 -79.755 -142.480 -79.585 ;
        RECT -135.780 -79.755 -132.560 -79.585 ;
        RECT -125.860 -79.755 -122.640 -79.585 ;
        RECT -115.940 -79.755 -112.720 -79.585 ;
        RECT -106.020 -79.755 -102.800 -79.585 ;
        RECT -96.100 -79.755 -92.880 -79.585 ;
        RECT -86.180 -79.755 -82.960 -79.585 ;
        RECT -76.260 -79.755 -73.040 -79.585 ;
        RECT -66.340 -79.755 -63.120 -79.585 ;
        RECT -56.420 -79.755 -53.200 -79.585 ;
        RECT -46.500 -79.755 -43.280 -79.585 ;
        RECT -36.580 -79.755 -33.360 -79.585 ;
        RECT -26.660 -79.755 -23.440 -79.585 ;
        RECT -16.740 -79.755 -13.520 -79.585 ;
        RECT -6.820 -79.755 -3.600 -79.585 ;
        RECT 3.100 -79.755 6.320 -79.585 ;
        RECT 13.020 -79.755 16.240 -79.585 ;
        RECT -283.595 -80.555 -283.285 -79.755 ;
        RECT -283.115 -80.480 -282.825 -79.755 ;
        RECT -282.655 -80.555 -282.345 -79.755 ;
        RECT -273.675 -80.555 -273.365 -79.755 ;
        RECT -273.195 -80.480 -272.905 -79.755 ;
        RECT -272.735 -80.555 -272.425 -79.755 ;
        RECT -263.755 -80.555 -263.445 -79.755 ;
        RECT -263.275 -80.480 -262.985 -79.755 ;
        RECT -262.815 -80.555 -262.505 -79.755 ;
        RECT -253.835 -80.555 -253.525 -79.755 ;
        RECT -253.355 -80.480 -253.065 -79.755 ;
        RECT -252.895 -80.555 -252.585 -79.755 ;
        RECT -243.915 -80.555 -243.605 -79.755 ;
        RECT -243.435 -80.480 -243.145 -79.755 ;
        RECT -242.975 -80.555 -242.665 -79.755 ;
        RECT -233.995 -80.555 -233.685 -79.755 ;
        RECT -233.515 -80.480 -233.225 -79.755 ;
        RECT -233.055 -80.555 -232.745 -79.755 ;
        RECT -224.075 -80.555 -223.765 -79.755 ;
        RECT -223.595 -80.480 -223.305 -79.755 ;
        RECT -223.135 -80.555 -222.825 -79.755 ;
        RECT -214.155 -80.555 -213.845 -79.755 ;
        RECT -213.675 -80.480 -213.385 -79.755 ;
        RECT -213.215 -80.555 -212.905 -79.755 ;
        RECT -204.235 -80.555 -203.925 -79.755 ;
        RECT -203.755 -80.480 -203.465 -79.755 ;
        RECT -203.295 -80.555 -202.985 -79.755 ;
        RECT -194.315 -80.555 -194.005 -79.755 ;
        RECT -193.835 -80.480 -193.545 -79.755 ;
        RECT -193.375 -80.555 -193.065 -79.755 ;
        RECT -184.395 -80.555 -184.085 -79.755 ;
        RECT -183.915 -80.480 -183.625 -79.755 ;
        RECT -183.455 -80.555 -183.145 -79.755 ;
        RECT -174.475 -80.555 -174.165 -79.755 ;
        RECT -173.995 -80.480 -173.705 -79.755 ;
        RECT -173.535 -80.555 -173.225 -79.755 ;
        RECT -164.555 -80.555 -164.245 -79.755 ;
        RECT -164.075 -80.480 -163.785 -79.755 ;
        RECT -163.615 -80.555 -163.305 -79.755 ;
        RECT -154.635 -80.555 -154.325 -79.755 ;
        RECT -154.155 -80.480 -153.865 -79.755 ;
        RECT -153.695 -80.555 -153.385 -79.755 ;
        RECT -144.715 -80.555 -144.405 -79.755 ;
        RECT -144.235 -80.480 -143.945 -79.755 ;
        RECT -143.775 -80.555 -143.465 -79.755 ;
        RECT -134.795 -80.555 -134.485 -79.755 ;
        RECT -134.315 -80.480 -134.025 -79.755 ;
        RECT -133.855 -80.555 -133.545 -79.755 ;
        RECT -124.875 -80.555 -124.565 -79.755 ;
        RECT -124.395 -80.480 -124.105 -79.755 ;
        RECT -123.935 -80.555 -123.625 -79.755 ;
        RECT -114.955 -80.555 -114.645 -79.755 ;
        RECT -114.475 -80.480 -114.185 -79.755 ;
        RECT -114.015 -80.555 -113.705 -79.755 ;
        RECT -105.035 -80.555 -104.725 -79.755 ;
        RECT -104.555 -80.480 -104.265 -79.755 ;
        RECT -104.095 -80.555 -103.785 -79.755 ;
        RECT -95.115 -80.555 -94.805 -79.755 ;
        RECT -94.635 -80.480 -94.345 -79.755 ;
        RECT -94.175 -80.555 -93.865 -79.755 ;
        RECT -85.195 -80.555 -84.885 -79.755 ;
        RECT -84.715 -80.480 -84.425 -79.755 ;
        RECT -84.255 -80.555 -83.945 -79.755 ;
        RECT -75.275 -80.555 -74.965 -79.755 ;
        RECT -74.795 -80.480 -74.505 -79.755 ;
        RECT -74.335 -80.555 -74.025 -79.755 ;
        RECT -65.355 -80.555 -65.045 -79.755 ;
        RECT -64.875 -80.480 -64.585 -79.755 ;
        RECT -64.415 -80.555 -64.105 -79.755 ;
        RECT -55.435 -80.555 -55.125 -79.755 ;
        RECT -54.955 -80.480 -54.665 -79.755 ;
        RECT -54.495 -80.555 -54.185 -79.755 ;
        RECT -45.515 -80.555 -45.205 -79.755 ;
        RECT -45.035 -80.480 -44.745 -79.755 ;
        RECT -44.575 -80.555 -44.265 -79.755 ;
        RECT -35.595 -80.555 -35.285 -79.755 ;
        RECT -35.115 -80.480 -34.825 -79.755 ;
        RECT -34.655 -80.555 -34.345 -79.755 ;
        RECT -25.675 -80.555 -25.365 -79.755 ;
        RECT -25.195 -80.480 -24.905 -79.755 ;
        RECT -24.735 -80.555 -24.425 -79.755 ;
        RECT -15.755 -80.555 -15.445 -79.755 ;
        RECT -15.275 -80.480 -14.985 -79.755 ;
        RECT -14.815 -80.555 -14.505 -79.755 ;
        RECT -5.835 -80.555 -5.525 -79.755 ;
        RECT -5.355 -80.480 -5.065 -79.755 ;
        RECT -4.895 -80.555 -4.585 -79.755 ;
        RECT 4.085 -80.555 4.395 -79.755 ;
        RECT 4.565 -80.480 4.855 -79.755 ;
        RECT 5.025 -80.555 5.335 -79.755 ;
        RECT 14.005 -80.555 14.315 -79.755 ;
        RECT 14.485 -80.480 14.775 -79.755 ;
        RECT 14.945 -80.555 15.255 -79.755 ;
        RECT -288.555 -82.305 -288.245 -81.505 ;
        RECT -288.075 -82.305 -287.785 -81.580 ;
        RECT -287.615 -82.305 -287.305 -81.505 ;
        RECT -278.635 -82.305 -278.325 -81.505 ;
        RECT -278.155 -82.305 -277.865 -81.580 ;
        RECT -277.695 -82.305 -277.385 -81.505 ;
        RECT -268.715 -82.305 -268.405 -81.505 ;
        RECT -268.235 -82.305 -267.945 -81.580 ;
        RECT -267.775 -82.305 -267.465 -81.505 ;
        RECT -258.795 -82.305 -258.485 -81.505 ;
        RECT -258.315 -82.305 -258.025 -81.580 ;
        RECT -257.855 -82.305 -257.545 -81.505 ;
        RECT -248.875 -82.305 -248.565 -81.505 ;
        RECT -248.395 -82.305 -248.105 -81.580 ;
        RECT -247.935 -82.305 -247.625 -81.505 ;
        RECT -238.955 -82.305 -238.645 -81.505 ;
        RECT -238.475 -82.305 -238.185 -81.580 ;
        RECT -238.015 -82.305 -237.705 -81.505 ;
        RECT -229.035 -82.305 -228.725 -81.505 ;
        RECT -228.555 -82.305 -228.265 -81.580 ;
        RECT -228.095 -82.305 -227.785 -81.505 ;
        RECT -219.115 -82.305 -218.805 -81.505 ;
        RECT -218.635 -82.305 -218.345 -81.580 ;
        RECT -218.175 -82.305 -217.865 -81.505 ;
        RECT -209.195 -82.305 -208.885 -81.505 ;
        RECT -208.715 -82.305 -208.425 -81.580 ;
        RECT -208.255 -82.305 -207.945 -81.505 ;
        RECT -199.275 -82.305 -198.965 -81.505 ;
        RECT -198.795 -82.305 -198.505 -81.580 ;
        RECT -198.335 -82.305 -198.025 -81.505 ;
        RECT -189.355 -82.305 -189.045 -81.505 ;
        RECT -188.875 -82.305 -188.585 -81.580 ;
        RECT -188.415 -82.305 -188.105 -81.505 ;
        RECT -179.435 -82.305 -179.125 -81.505 ;
        RECT -178.955 -82.305 -178.665 -81.580 ;
        RECT -178.495 -82.305 -178.185 -81.505 ;
        RECT -169.515 -82.305 -169.205 -81.505 ;
        RECT -169.035 -82.305 -168.745 -81.580 ;
        RECT -168.575 -82.305 -168.265 -81.505 ;
        RECT -159.595 -82.305 -159.285 -81.505 ;
        RECT -159.115 -82.305 -158.825 -81.580 ;
        RECT -158.655 -82.305 -158.345 -81.505 ;
        RECT -149.675 -82.305 -149.365 -81.505 ;
        RECT -149.195 -82.305 -148.905 -81.580 ;
        RECT -148.735 -82.305 -148.425 -81.505 ;
        RECT -139.755 -82.305 -139.445 -81.505 ;
        RECT -139.275 -82.305 -138.985 -81.580 ;
        RECT -138.815 -82.305 -138.505 -81.505 ;
        RECT -129.835 -82.305 -129.525 -81.505 ;
        RECT -129.355 -82.305 -129.065 -81.580 ;
        RECT -128.895 -82.305 -128.585 -81.505 ;
        RECT -119.915 -82.305 -119.605 -81.505 ;
        RECT -119.435 -82.305 -119.145 -81.580 ;
        RECT -118.975 -82.305 -118.665 -81.505 ;
        RECT -109.995 -82.305 -109.685 -81.505 ;
        RECT -109.515 -82.305 -109.225 -81.580 ;
        RECT -109.055 -82.305 -108.745 -81.505 ;
        RECT -100.075 -82.305 -99.765 -81.505 ;
        RECT -99.595 -82.305 -99.305 -81.580 ;
        RECT -99.135 -82.305 -98.825 -81.505 ;
        RECT -90.155 -82.305 -89.845 -81.505 ;
        RECT -89.675 -82.305 -89.385 -81.580 ;
        RECT -89.215 -82.305 -88.905 -81.505 ;
        RECT -80.235 -82.305 -79.925 -81.505 ;
        RECT -79.755 -82.305 -79.465 -81.580 ;
        RECT -79.295 -82.305 -78.985 -81.505 ;
        RECT -70.315 -82.305 -70.005 -81.505 ;
        RECT -69.835 -82.305 -69.545 -81.580 ;
        RECT -69.375 -82.305 -69.065 -81.505 ;
        RECT -60.395 -82.305 -60.085 -81.505 ;
        RECT -59.915 -82.305 -59.625 -81.580 ;
        RECT -59.455 -82.305 -59.145 -81.505 ;
        RECT -50.475 -82.305 -50.165 -81.505 ;
        RECT -49.995 -82.305 -49.705 -81.580 ;
        RECT -49.535 -82.305 -49.225 -81.505 ;
        RECT -40.555 -82.305 -40.245 -81.505 ;
        RECT -40.075 -82.305 -39.785 -81.580 ;
        RECT -39.615 -82.305 -39.305 -81.505 ;
        RECT -30.635 -82.305 -30.325 -81.505 ;
        RECT -30.155 -82.305 -29.865 -81.580 ;
        RECT -29.695 -82.305 -29.385 -81.505 ;
        RECT -20.715 -82.305 -20.405 -81.505 ;
        RECT -20.235 -82.305 -19.945 -81.580 ;
        RECT -19.775 -82.305 -19.465 -81.505 ;
        RECT -10.795 -82.305 -10.485 -81.505 ;
        RECT -10.315 -82.305 -10.025 -81.580 ;
        RECT -9.855 -82.305 -9.545 -81.505 ;
        RECT -0.875 -82.305 -0.565 -81.505 ;
        RECT -0.395 -82.305 -0.105 -81.580 ;
        RECT 0.065 -82.305 0.375 -81.505 ;
        RECT 9.045 -82.305 9.355 -81.505 ;
        RECT 9.525 -82.305 9.815 -81.580 ;
        RECT 9.985 -82.305 10.295 -81.505 ;
        RECT 18.965 -82.305 19.275 -81.505 ;
        RECT 19.445 -82.305 19.735 -81.580 ;
        RECT 19.905 -82.305 20.215 -81.505 ;
        RECT -289.540 -82.475 -286.320 -82.305 ;
        RECT -279.620 -82.475 -276.400 -82.305 ;
        RECT -269.700 -82.475 -266.480 -82.305 ;
        RECT -259.780 -82.475 -256.560 -82.305 ;
        RECT -249.860 -82.475 -246.640 -82.305 ;
        RECT -239.940 -82.475 -236.720 -82.305 ;
        RECT -230.020 -82.475 -226.800 -82.305 ;
        RECT -220.100 -82.475 -216.880 -82.305 ;
        RECT -210.180 -82.475 -206.960 -82.305 ;
        RECT -200.260 -82.475 -197.040 -82.305 ;
        RECT -190.340 -82.475 -187.120 -82.305 ;
        RECT -180.420 -82.475 -177.200 -82.305 ;
        RECT -170.500 -82.475 -167.280 -82.305 ;
        RECT -160.580 -82.475 -157.360 -82.305 ;
        RECT -150.660 -82.475 -147.440 -82.305 ;
        RECT -140.740 -82.475 -137.520 -82.305 ;
        RECT -130.820 -82.475 -127.600 -82.305 ;
        RECT -120.900 -82.475 -117.680 -82.305 ;
        RECT -110.980 -82.475 -107.760 -82.305 ;
        RECT -101.060 -82.475 -97.840 -82.305 ;
        RECT -91.140 -82.475 -87.920 -82.305 ;
        RECT -81.220 -82.475 -78.000 -82.305 ;
        RECT -71.300 -82.475 -68.080 -82.305 ;
        RECT -61.380 -82.475 -58.160 -82.305 ;
        RECT -51.460 -82.475 -48.240 -82.305 ;
        RECT -41.540 -82.475 -38.320 -82.305 ;
        RECT -31.620 -82.475 -28.400 -82.305 ;
        RECT -21.700 -82.475 -18.480 -82.305 ;
        RECT -11.780 -82.475 -8.560 -82.305 ;
        RECT -1.860 -82.475 1.360 -82.305 ;
        RECT 8.060 -82.475 11.280 -82.305 ;
        RECT 17.980 -82.475 21.200 -82.305 ;
        RECT -284.825 -83.345 -284.655 -82.820 ;
        RECT -285.205 -83.675 -284.655 -83.345 ;
        RECT -284.825 -84.200 -284.655 -83.675 ;
        RECT -283.115 -83.695 -282.825 -82.970 ;
        RECT -281.285 -83.345 -281.115 -82.820 ;
        RECT -274.905 -83.345 -274.735 -82.820 ;
        RECT -281.285 -83.675 -280.735 -83.345 ;
        RECT -275.285 -83.675 -274.735 -83.345 ;
        RECT -283.200 -83.865 -282.740 -83.695 ;
        RECT -281.285 -84.200 -281.115 -83.675 ;
        RECT -274.905 -84.200 -274.735 -83.675 ;
        RECT -273.195 -83.695 -272.905 -82.970 ;
        RECT -271.365 -83.345 -271.195 -82.820 ;
        RECT -264.985 -83.345 -264.815 -82.820 ;
        RECT -271.365 -83.675 -270.815 -83.345 ;
        RECT -265.365 -83.675 -264.815 -83.345 ;
        RECT -273.280 -83.865 -272.820 -83.695 ;
        RECT -271.365 -84.200 -271.195 -83.675 ;
        RECT -264.985 -84.200 -264.815 -83.675 ;
        RECT -263.275 -83.695 -262.985 -82.970 ;
        RECT -261.445 -83.345 -261.275 -82.820 ;
        RECT -255.065 -83.345 -254.895 -82.820 ;
        RECT -261.445 -83.675 -260.895 -83.345 ;
        RECT -255.445 -83.675 -254.895 -83.345 ;
        RECT -263.360 -83.865 -262.900 -83.695 ;
        RECT -261.445 -84.200 -261.275 -83.675 ;
        RECT -255.065 -84.200 -254.895 -83.675 ;
        RECT -253.355 -83.695 -253.065 -82.970 ;
        RECT -251.525 -83.345 -251.355 -82.820 ;
        RECT -245.145 -83.345 -244.975 -82.820 ;
        RECT -251.525 -83.675 -250.975 -83.345 ;
        RECT -245.525 -83.675 -244.975 -83.345 ;
        RECT -253.440 -83.865 -252.980 -83.695 ;
        RECT -251.525 -84.200 -251.355 -83.675 ;
        RECT -245.145 -84.200 -244.975 -83.675 ;
        RECT -243.435 -83.695 -243.145 -82.970 ;
        RECT -241.605 -83.345 -241.435 -82.820 ;
        RECT -235.225 -83.345 -235.055 -82.820 ;
        RECT -241.605 -83.675 -241.055 -83.345 ;
        RECT -235.605 -83.675 -235.055 -83.345 ;
        RECT -243.520 -83.865 -243.060 -83.695 ;
        RECT -241.605 -84.200 -241.435 -83.675 ;
        RECT -235.225 -84.200 -235.055 -83.675 ;
        RECT -233.515 -83.695 -233.225 -82.970 ;
        RECT -231.685 -83.345 -231.515 -82.820 ;
        RECT -225.305 -83.345 -225.135 -82.820 ;
        RECT -231.685 -83.675 -231.135 -83.345 ;
        RECT -225.685 -83.675 -225.135 -83.345 ;
        RECT -233.600 -83.865 -233.140 -83.695 ;
        RECT -231.685 -84.200 -231.515 -83.675 ;
        RECT -225.305 -84.200 -225.135 -83.675 ;
        RECT -223.595 -83.695 -223.305 -82.970 ;
        RECT -221.765 -83.345 -221.595 -82.820 ;
        RECT -215.385 -83.345 -215.215 -82.820 ;
        RECT -221.765 -83.675 -221.215 -83.345 ;
        RECT -215.765 -83.675 -215.215 -83.345 ;
        RECT -223.680 -83.865 -223.220 -83.695 ;
        RECT -221.765 -84.200 -221.595 -83.675 ;
        RECT -215.385 -84.200 -215.215 -83.675 ;
        RECT -213.675 -83.695 -213.385 -82.970 ;
        RECT -211.845 -83.345 -211.675 -82.820 ;
        RECT -205.465 -83.345 -205.295 -82.820 ;
        RECT -211.845 -83.675 -211.295 -83.345 ;
        RECT -205.845 -83.675 -205.295 -83.345 ;
        RECT -213.760 -83.865 -213.300 -83.695 ;
        RECT -211.845 -84.200 -211.675 -83.675 ;
        RECT -205.465 -84.200 -205.295 -83.675 ;
        RECT -203.755 -83.695 -203.465 -82.970 ;
        RECT -201.925 -83.345 -201.755 -82.820 ;
        RECT -195.545 -83.345 -195.375 -82.820 ;
        RECT -201.925 -83.675 -201.375 -83.345 ;
        RECT -195.925 -83.675 -195.375 -83.345 ;
        RECT -203.840 -83.865 -203.380 -83.695 ;
        RECT -201.925 -84.200 -201.755 -83.675 ;
        RECT -195.545 -84.200 -195.375 -83.675 ;
        RECT -193.835 -83.695 -193.545 -82.970 ;
        RECT -192.005 -83.345 -191.835 -82.820 ;
        RECT -185.625 -83.345 -185.455 -82.820 ;
        RECT -192.005 -83.675 -191.455 -83.345 ;
        RECT -186.005 -83.675 -185.455 -83.345 ;
        RECT -193.920 -83.865 -193.460 -83.695 ;
        RECT -192.005 -84.200 -191.835 -83.675 ;
        RECT -185.625 -84.200 -185.455 -83.675 ;
        RECT -183.915 -83.695 -183.625 -82.970 ;
        RECT -182.085 -83.345 -181.915 -82.820 ;
        RECT -175.705 -83.345 -175.535 -82.820 ;
        RECT -182.085 -83.675 -181.535 -83.345 ;
        RECT -176.085 -83.675 -175.535 -83.345 ;
        RECT -184.000 -83.865 -183.540 -83.695 ;
        RECT -182.085 -84.200 -181.915 -83.675 ;
        RECT -175.705 -84.200 -175.535 -83.675 ;
        RECT -173.995 -83.695 -173.705 -82.970 ;
        RECT -172.165 -83.345 -171.995 -82.820 ;
        RECT -165.785 -83.345 -165.615 -82.820 ;
        RECT -172.165 -83.675 -171.615 -83.345 ;
        RECT -166.165 -83.675 -165.615 -83.345 ;
        RECT -174.080 -83.865 -173.620 -83.695 ;
        RECT -172.165 -84.200 -171.995 -83.675 ;
        RECT -165.785 -84.200 -165.615 -83.675 ;
        RECT -164.075 -83.695 -163.785 -82.970 ;
        RECT -162.245 -83.345 -162.075 -82.820 ;
        RECT -155.865 -83.345 -155.695 -82.820 ;
        RECT -162.245 -83.675 -161.695 -83.345 ;
        RECT -156.245 -83.675 -155.695 -83.345 ;
        RECT -164.160 -83.865 -163.700 -83.695 ;
        RECT -162.245 -84.200 -162.075 -83.675 ;
        RECT -155.865 -84.200 -155.695 -83.675 ;
        RECT -154.155 -83.695 -153.865 -82.970 ;
        RECT -152.325 -83.345 -152.155 -82.820 ;
        RECT -145.945 -83.345 -145.775 -82.820 ;
        RECT -152.325 -83.675 -151.775 -83.345 ;
        RECT -146.325 -83.675 -145.775 -83.345 ;
        RECT -154.240 -83.865 -153.780 -83.695 ;
        RECT -152.325 -84.200 -152.155 -83.675 ;
        RECT -145.945 -84.200 -145.775 -83.675 ;
        RECT -144.235 -83.695 -143.945 -82.970 ;
        RECT -142.405 -83.345 -142.235 -82.820 ;
        RECT -136.025 -83.345 -135.855 -82.820 ;
        RECT -142.405 -83.675 -141.855 -83.345 ;
        RECT -136.405 -83.675 -135.855 -83.345 ;
        RECT -144.320 -83.865 -143.860 -83.695 ;
        RECT -142.405 -84.200 -142.235 -83.675 ;
        RECT -136.025 -84.200 -135.855 -83.675 ;
        RECT -134.315 -83.695 -134.025 -82.970 ;
        RECT -132.485 -83.345 -132.315 -82.820 ;
        RECT -126.105 -83.345 -125.935 -82.820 ;
        RECT -132.485 -83.675 -131.935 -83.345 ;
        RECT -126.485 -83.675 -125.935 -83.345 ;
        RECT -134.400 -83.865 -133.940 -83.695 ;
        RECT -132.485 -84.200 -132.315 -83.675 ;
        RECT -126.105 -84.200 -125.935 -83.675 ;
        RECT -124.395 -83.695 -124.105 -82.970 ;
        RECT -122.565 -83.345 -122.395 -82.820 ;
        RECT -116.185 -83.345 -116.015 -82.820 ;
        RECT -122.565 -83.675 -122.015 -83.345 ;
        RECT -116.565 -83.675 -116.015 -83.345 ;
        RECT -124.480 -83.865 -124.020 -83.695 ;
        RECT -122.565 -84.200 -122.395 -83.675 ;
        RECT -116.185 -84.200 -116.015 -83.675 ;
        RECT -114.475 -83.695 -114.185 -82.970 ;
        RECT -112.645 -83.345 -112.475 -82.820 ;
        RECT -106.265 -83.345 -106.095 -82.820 ;
        RECT -112.645 -83.675 -112.095 -83.345 ;
        RECT -106.645 -83.675 -106.095 -83.345 ;
        RECT -114.560 -83.865 -114.100 -83.695 ;
        RECT -112.645 -84.200 -112.475 -83.675 ;
        RECT -106.265 -84.200 -106.095 -83.675 ;
        RECT -104.555 -83.695 -104.265 -82.970 ;
        RECT -102.725 -83.345 -102.555 -82.820 ;
        RECT -96.345 -83.345 -96.175 -82.820 ;
        RECT -102.725 -83.675 -102.175 -83.345 ;
        RECT -96.725 -83.675 -96.175 -83.345 ;
        RECT -104.640 -83.865 -104.180 -83.695 ;
        RECT -102.725 -84.200 -102.555 -83.675 ;
        RECT -96.345 -84.200 -96.175 -83.675 ;
        RECT -94.635 -83.695 -94.345 -82.970 ;
        RECT -92.805 -83.345 -92.635 -82.820 ;
        RECT -86.425 -83.345 -86.255 -82.820 ;
        RECT -92.805 -83.675 -92.255 -83.345 ;
        RECT -86.805 -83.675 -86.255 -83.345 ;
        RECT -94.720 -83.865 -94.260 -83.695 ;
        RECT -92.805 -84.200 -92.635 -83.675 ;
        RECT -86.425 -84.200 -86.255 -83.675 ;
        RECT -84.715 -83.695 -84.425 -82.970 ;
        RECT -82.885 -83.345 -82.715 -82.820 ;
        RECT -76.505 -83.345 -76.335 -82.820 ;
        RECT -82.885 -83.675 -82.335 -83.345 ;
        RECT -76.885 -83.675 -76.335 -83.345 ;
        RECT -84.800 -83.865 -84.340 -83.695 ;
        RECT -82.885 -84.200 -82.715 -83.675 ;
        RECT -76.505 -84.200 -76.335 -83.675 ;
        RECT -74.795 -83.695 -74.505 -82.970 ;
        RECT -72.965 -83.345 -72.795 -82.820 ;
        RECT -66.585 -83.345 -66.415 -82.820 ;
        RECT -72.965 -83.675 -72.415 -83.345 ;
        RECT -66.965 -83.675 -66.415 -83.345 ;
        RECT -74.880 -83.865 -74.420 -83.695 ;
        RECT -72.965 -84.200 -72.795 -83.675 ;
        RECT -66.585 -84.200 -66.415 -83.675 ;
        RECT -64.875 -83.695 -64.585 -82.970 ;
        RECT -63.045 -83.345 -62.875 -82.820 ;
        RECT -56.665 -83.345 -56.495 -82.820 ;
        RECT -63.045 -83.675 -62.495 -83.345 ;
        RECT -57.045 -83.675 -56.495 -83.345 ;
        RECT -64.960 -83.865 -64.500 -83.695 ;
        RECT -63.045 -84.200 -62.875 -83.675 ;
        RECT -56.665 -84.200 -56.495 -83.675 ;
        RECT -54.955 -83.695 -54.665 -82.970 ;
        RECT -53.125 -83.345 -52.955 -82.820 ;
        RECT -46.745 -83.345 -46.575 -82.820 ;
        RECT -53.125 -83.675 -52.575 -83.345 ;
        RECT -47.125 -83.675 -46.575 -83.345 ;
        RECT -55.040 -83.865 -54.580 -83.695 ;
        RECT -53.125 -84.200 -52.955 -83.675 ;
        RECT -46.745 -84.200 -46.575 -83.675 ;
        RECT -45.035 -83.695 -44.745 -82.970 ;
        RECT -43.205 -83.345 -43.035 -82.820 ;
        RECT -36.825 -83.345 -36.655 -82.820 ;
        RECT -43.205 -83.675 -42.655 -83.345 ;
        RECT -37.205 -83.675 -36.655 -83.345 ;
        RECT -45.120 -83.865 -44.660 -83.695 ;
        RECT -43.205 -84.200 -43.035 -83.675 ;
        RECT -36.825 -84.200 -36.655 -83.675 ;
        RECT -35.115 -83.695 -34.825 -82.970 ;
        RECT -33.285 -83.345 -33.115 -82.820 ;
        RECT -26.905 -83.345 -26.735 -82.820 ;
        RECT -33.285 -83.675 -32.735 -83.345 ;
        RECT -27.285 -83.675 -26.735 -83.345 ;
        RECT -35.200 -83.865 -34.740 -83.695 ;
        RECT -33.285 -84.200 -33.115 -83.675 ;
        RECT -26.905 -84.200 -26.735 -83.675 ;
        RECT -25.195 -83.695 -24.905 -82.970 ;
        RECT -23.365 -83.345 -23.195 -82.820 ;
        RECT -16.985 -83.345 -16.815 -82.820 ;
        RECT -23.365 -83.675 -22.815 -83.345 ;
        RECT -17.365 -83.675 -16.815 -83.345 ;
        RECT -25.280 -83.865 -24.820 -83.695 ;
        RECT -23.365 -84.200 -23.195 -83.675 ;
        RECT -16.985 -84.200 -16.815 -83.675 ;
        RECT -15.275 -83.695 -14.985 -82.970 ;
        RECT -13.445 -83.345 -13.275 -82.820 ;
        RECT -7.065 -83.345 -6.895 -82.820 ;
        RECT -13.445 -83.675 -12.895 -83.345 ;
        RECT -7.445 -83.675 -6.895 -83.345 ;
        RECT -15.360 -83.865 -14.900 -83.695 ;
        RECT -13.445 -84.200 -13.275 -83.675 ;
        RECT -7.065 -84.200 -6.895 -83.675 ;
        RECT -5.355 -83.695 -5.065 -82.970 ;
        RECT -3.525 -83.345 -3.355 -82.820 ;
        RECT 2.855 -83.345 3.025 -82.820 ;
        RECT -3.525 -83.675 -2.975 -83.345 ;
        RECT 2.475 -83.675 3.025 -83.345 ;
        RECT -5.440 -83.865 -4.980 -83.695 ;
        RECT -3.525 -84.200 -3.355 -83.675 ;
        RECT 2.855 -84.200 3.025 -83.675 ;
        RECT 4.565 -83.695 4.855 -82.970 ;
        RECT 6.395 -83.345 6.565 -82.820 ;
        RECT 12.775 -83.345 12.945 -82.820 ;
        RECT 6.395 -83.675 6.945 -83.345 ;
        RECT 12.395 -83.675 12.945 -83.345 ;
        RECT 4.480 -83.865 4.940 -83.695 ;
        RECT 6.395 -84.200 6.565 -83.675 ;
        RECT 12.775 -84.200 12.945 -83.675 ;
        RECT 14.485 -83.695 14.775 -82.970 ;
        RECT 16.315 -83.345 16.485 -82.820 ;
        RECT 16.315 -83.675 16.865 -83.345 ;
        RECT 14.400 -83.865 14.860 -83.695 ;
        RECT 16.315 -84.200 16.485 -83.675 ;
        RECT -291.545 -172.965 -291.375 -172.440 ;
        RECT -289.920 -172.855 -289.460 -172.685 ;
        RECT -291.925 -173.295 -291.375 -172.965 ;
        RECT -291.545 -173.820 -291.375 -173.295 ;
        RECT -289.835 -173.580 -289.545 -172.855 ;
        RECT -288.005 -172.965 -287.835 -172.440 ;
        RECT -281.625 -172.965 -281.455 -172.440 ;
        RECT -280.000 -172.855 -279.540 -172.685 ;
        RECT -288.005 -173.295 -287.455 -172.965 ;
        RECT -282.005 -173.295 -281.455 -172.965 ;
        RECT -288.005 -173.820 -287.835 -173.295 ;
        RECT -281.625 -173.820 -281.455 -173.295 ;
        RECT -279.915 -173.580 -279.625 -172.855 ;
        RECT -278.085 -172.965 -277.915 -172.440 ;
        RECT -271.705 -172.965 -271.535 -172.440 ;
        RECT -270.080 -172.855 -269.620 -172.685 ;
        RECT -278.085 -173.295 -277.535 -172.965 ;
        RECT -272.085 -173.295 -271.535 -172.965 ;
        RECT -278.085 -173.820 -277.915 -173.295 ;
        RECT -271.705 -173.820 -271.535 -173.295 ;
        RECT -269.995 -173.580 -269.705 -172.855 ;
        RECT -268.165 -172.965 -267.995 -172.440 ;
        RECT -261.785 -172.965 -261.615 -172.440 ;
        RECT -260.160 -172.855 -259.700 -172.685 ;
        RECT -268.165 -173.295 -267.615 -172.965 ;
        RECT -262.165 -173.295 -261.615 -172.965 ;
        RECT -268.165 -173.820 -267.995 -173.295 ;
        RECT -261.785 -173.820 -261.615 -173.295 ;
        RECT -260.075 -173.580 -259.785 -172.855 ;
        RECT -258.245 -172.965 -258.075 -172.440 ;
        RECT -251.865 -172.965 -251.695 -172.440 ;
        RECT -250.240 -172.855 -249.780 -172.685 ;
        RECT -258.245 -173.295 -257.695 -172.965 ;
        RECT -252.245 -173.295 -251.695 -172.965 ;
        RECT -258.245 -173.820 -258.075 -173.295 ;
        RECT -251.865 -173.820 -251.695 -173.295 ;
        RECT -250.155 -173.580 -249.865 -172.855 ;
        RECT -248.325 -172.965 -248.155 -172.440 ;
        RECT -241.945 -172.965 -241.775 -172.440 ;
        RECT -240.320 -172.855 -239.860 -172.685 ;
        RECT -248.325 -173.295 -247.775 -172.965 ;
        RECT -242.325 -173.295 -241.775 -172.965 ;
        RECT -248.325 -173.820 -248.155 -173.295 ;
        RECT -241.945 -173.820 -241.775 -173.295 ;
        RECT -240.235 -173.580 -239.945 -172.855 ;
        RECT -238.405 -172.965 -238.235 -172.440 ;
        RECT -232.025 -172.965 -231.855 -172.440 ;
        RECT -230.400 -172.855 -229.940 -172.685 ;
        RECT -238.405 -173.295 -237.855 -172.965 ;
        RECT -232.405 -173.295 -231.855 -172.965 ;
        RECT -238.405 -173.820 -238.235 -173.295 ;
        RECT -232.025 -173.820 -231.855 -173.295 ;
        RECT -230.315 -173.580 -230.025 -172.855 ;
        RECT -228.485 -172.965 -228.315 -172.440 ;
        RECT -222.105 -172.965 -221.935 -172.440 ;
        RECT -220.480 -172.855 -220.020 -172.685 ;
        RECT -228.485 -173.295 -227.935 -172.965 ;
        RECT -222.485 -173.295 -221.935 -172.965 ;
        RECT -228.485 -173.820 -228.315 -173.295 ;
        RECT -222.105 -173.820 -221.935 -173.295 ;
        RECT -220.395 -173.580 -220.105 -172.855 ;
        RECT -218.565 -172.965 -218.395 -172.440 ;
        RECT -212.185 -172.965 -212.015 -172.440 ;
        RECT -210.560 -172.855 -210.100 -172.685 ;
        RECT -218.565 -173.295 -218.015 -172.965 ;
        RECT -212.565 -173.295 -212.015 -172.965 ;
        RECT -218.565 -173.820 -218.395 -173.295 ;
        RECT -212.185 -173.820 -212.015 -173.295 ;
        RECT -210.475 -173.580 -210.185 -172.855 ;
        RECT -208.645 -172.965 -208.475 -172.440 ;
        RECT -202.265 -172.965 -202.095 -172.440 ;
        RECT -200.640 -172.855 -200.180 -172.685 ;
        RECT -208.645 -173.295 -208.095 -172.965 ;
        RECT -202.645 -173.295 -202.095 -172.965 ;
        RECT -208.645 -173.820 -208.475 -173.295 ;
        RECT -202.265 -173.820 -202.095 -173.295 ;
        RECT -200.555 -173.580 -200.265 -172.855 ;
        RECT -198.725 -172.965 -198.555 -172.440 ;
        RECT -192.345 -172.965 -192.175 -172.440 ;
        RECT -190.720 -172.855 -190.260 -172.685 ;
        RECT -198.725 -173.295 -198.175 -172.965 ;
        RECT -192.725 -173.295 -192.175 -172.965 ;
        RECT -198.725 -173.820 -198.555 -173.295 ;
        RECT -192.345 -173.820 -192.175 -173.295 ;
        RECT -190.635 -173.580 -190.345 -172.855 ;
        RECT -188.805 -172.965 -188.635 -172.440 ;
        RECT -182.425 -172.965 -182.255 -172.440 ;
        RECT -180.800 -172.855 -180.340 -172.685 ;
        RECT -188.805 -173.295 -188.255 -172.965 ;
        RECT -182.805 -173.295 -182.255 -172.965 ;
        RECT -188.805 -173.820 -188.635 -173.295 ;
        RECT -182.425 -173.820 -182.255 -173.295 ;
        RECT -180.715 -173.580 -180.425 -172.855 ;
        RECT -178.885 -172.965 -178.715 -172.440 ;
        RECT -172.505 -172.965 -172.335 -172.440 ;
        RECT -170.880 -172.855 -170.420 -172.685 ;
        RECT -178.885 -173.295 -178.335 -172.965 ;
        RECT -172.885 -173.295 -172.335 -172.965 ;
        RECT -178.885 -173.820 -178.715 -173.295 ;
        RECT -172.505 -173.820 -172.335 -173.295 ;
        RECT -170.795 -173.580 -170.505 -172.855 ;
        RECT -168.965 -172.965 -168.795 -172.440 ;
        RECT -162.585 -172.965 -162.415 -172.440 ;
        RECT -160.960 -172.855 -160.500 -172.685 ;
        RECT -168.965 -173.295 -168.415 -172.965 ;
        RECT -162.965 -173.295 -162.415 -172.965 ;
        RECT -168.965 -173.820 -168.795 -173.295 ;
        RECT -162.585 -173.820 -162.415 -173.295 ;
        RECT -160.875 -173.580 -160.585 -172.855 ;
        RECT -159.045 -172.965 -158.875 -172.440 ;
        RECT -152.665 -172.965 -152.495 -172.440 ;
        RECT -151.040 -172.855 -150.580 -172.685 ;
        RECT -159.045 -173.295 -158.495 -172.965 ;
        RECT -153.045 -173.295 -152.495 -172.965 ;
        RECT -159.045 -173.820 -158.875 -173.295 ;
        RECT -152.665 -173.820 -152.495 -173.295 ;
        RECT -150.955 -173.580 -150.665 -172.855 ;
        RECT -149.125 -172.965 -148.955 -172.440 ;
        RECT -142.745 -172.965 -142.575 -172.440 ;
        RECT -141.120 -172.855 -140.660 -172.685 ;
        RECT -149.125 -173.295 -148.575 -172.965 ;
        RECT -143.125 -173.295 -142.575 -172.965 ;
        RECT -149.125 -173.820 -148.955 -173.295 ;
        RECT -142.745 -173.820 -142.575 -173.295 ;
        RECT -141.035 -173.580 -140.745 -172.855 ;
        RECT -139.205 -172.965 -139.035 -172.440 ;
        RECT -132.825 -172.965 -132.655 -172.440 ;
        RECT -131.200 -172.855 -130.740 -172.685 ;
        RECT -139.205 -173.295 -138.655 -172.965 ;
        RECT -133.205 -173.295 -132.655 -172.965 ;
        RECT -139.205 -173.820 -139.035 -173.295 ;
        RECT -132.825 -173.820 -132.655 -173.295 ;
        RECT -131.115 -173.580 -130.825 -172.855 ;
        RECT -129.285 -172.965 -129.115 -172.440 ;
        RECT -122.905 -172.965 -122.735 -172.440 ;
        RECT -121.280 -172.855 -120.820 -172.685 ;
        RECT -129.285 -173.295 -128.735 -172.965 ;
        RECT -123.285 -173.295 -122.735 -172.965 ;
        RECT -129.285 -173.820 -129.115 -173.295 ;
        RECT -122.905 -173.820 -122.735 -173.295 ;
        RECT -121.195 -173.580 -120.905 -172.855 ;
        RECT -119.365 -172.965 -119.195 -172.440 ;
        RECT -112.985 -172.965 -112.815 -172.440 ;
        RECT -111.360 -172.855 -110.900 -172.685 ;
        RECT -119.365 -173.295 -118.815 -172.965 ;
        RECT -113.365 -173.295 -112.815 -172.965 ;
        RECT -119.365 -173.820 -119.195 -173.295 ;
        RECT -112.985 -173.820 -112.815 -173.295 ;
        RECT -111.275 -173.580 -110.985 -172.855 ;
        RECT -109.445 -172.965 -109.275 -172.440 ;
        RECT -103.065 -172.965 -102.895 -172.440 ;
        RECT -101.440 -172.855 -100.980 -172.685 ;
        RECT -109.445 -173.295 -108.895 -172.965 ;
        RECT -103.445 -173.295 -102.895 -172.965 ;
        RECT -109.445 -173.820 -109.275 -173.295 ;
        RECT -103.065 -173.820 -102.895 -173.295 ;
        RECT -101.355 -173.580 -101.065 -172.855 ;
        RECT -99.525 -172.965 -99.355 -172.440 ;
        RECT -93.145 -172.965 -92.975 -172.440 ;
        RECT -91.520 -172.855 -91.060 -172.685 ;
        RECT -99.525 -173.295 -98.975 -172.965 ;
        RECT -93.525 -173.295 -92.975 -172.965 ;
        RECT -99.525 -173.820 -99.355 -173.295 ;
        RECT -93.145 -173.820 -92.975 -173.295 ;
        RECT -91.435 -173.580 -91.145 -172.855 ;
        RECT -89.605 -172.965 -89.435 -172.440 ;
        RECT -83.225 -172.965 -83.055 -172.440 ;
        RECT -81.600 -172.855 -81.140 -172.685 ;
        RECT -89.605 -173.295 -89.055 -172.965 ;
        RECT -83.605 -173.295 -83.055 -172.965 ;
        RECT -89.605 -173.820 -89.435 -173.295 ;
        RECT -83.225 -173.820 -83.055 -173.295 ;
        RECT -81.515 -173.580 -81.225 -172.855 ;
        RECT -79.685 -172.965 -79.515 -172.440 ;
        RECT -73.305 -172.965 -73.135 -172.440 ;
        RECT -71.680 -172.855 -71.220 -172.685 ;
        RECT -79.685 -173.295 -79.135 -172.965 ;
        RECT -73.685 -173.295 -73.135 -172.965 ;
        RECT -79.685 -173.820 -79.515 -173.295 ;
        RECT -73.305 -173.820 -73.135 -173.295 ;
        RECT -71.595 -173.580 -71.305 -172.855 ;
        RECT -69.765 -172.965 -69.595 -172.440 ;
        RECT -63.385 -172.965 -63.215 -172.440 ;
        RECT -61.760 -172.855 -61.300 -172.685 ;
        RECT -69.765 -173.295 -69.215 -172.965 ;
        RECT -63.765 -173.295 -63.215 -172.965 ;
        RECT -69.765 -173.820 -69.595 -173.295 ;
        RECT -63.385 -173.820 -63.215 -173.295 ;
        RECT -61.675 -173.580 -61.385 -172.855 ;
        RECT -59.845 -172.965 -59.675 -172.440 ;
        RECT -53.465 -172.965 -53.295 -172.440 ;
        RECT -51.840 -172.855 -51.380 -172.685 ;
        RECT -59.845 -173.295 -59.295 -172.965 ;
        RECT -53.845 -173.295 -53.295 -172.965 ;
        RECT -59.845 -173.820 -59.675 -173.295 ;
        RECT -53.465 -173.820 -53.295 -173.295 ;
        RECT -51.755 -173.580 -51.465 -172.855 ;
        RECT -49.925 -172.965 -49.755 -172.440 ;
        RECT -43.545 -172.965 -43.375 -172.440 ;
        RECT -41.920 -172.855 -41.460 -172.685 ;
        RECT -49.925 -173.295 -49.375 -172.965 ;
        RECT -43.925 -173.295 -43.375 -172.965 ;
        RECT -49.925 -173.820 -49.755 -173.295 ;
        RECT -43.545 -173.820 -43.375 -173.295 ;
        RECT -41.835 -173.580 -41.545 -172.855 ;
        RECT -40.005 -172.965 -39.835 -172.440 ;
        RECT -33.625 -172.965 -33.455 -172.440 ;
        RECT -32.000 -172.855 -31.540 -172.685 ;
        RECT -40.005 -173.295 -39.455 -172.965 ;
        RECT -34.005 -173.295 -33.455 -172.965 ;
        RECT -40.005 -173.820 -39.835 -173.295 ;
        RECT -33.625 -173.820 -33.455 -173.295 ;
        RECT -31.915 -173.580 -31.625 -172.855 ;
        RECT -30.085 -172.965 -29.915 -172.440 ;
        RECT -23.705 -172.965 -23.535 -172.440 ;
        RECT -22.080 -172.855 -21.620 -172.685 ;
        RECT -30.085 -173.295 -29.535 -172.965 ;
        RECT -24.085 -173.295 -23.535 -172.965 ;
        RECT -30.085 -173.820 -29.915 -173.295 ;
        RECT -23.705 -173.820 -23.535 -173.295 ;
        RECT -21.995 -173.580 -21.705 -172.855 ;
        RECT -20.165 -172.965 -19.995 -172.440 ;
        RECT -13.785 -172.965 -13.615 -172.440 ;
        RECT -12.160 -172.855 -11.700 -172.685 ;
        RECT -20.165 -173.295 -19.615 -172.965 ;
        RECT -14.165 -173.295 -13.615 -172.965 ;
        RECT -20.165 -173.820 -19.995 -173.295 ;
        RECT -13.785 -173.820 -13.615 -173.295 ;
        RECT -12.075 -173.580 -11.785 -172.855 ;
        RECT -10.245 -172.965 -10.075 -172.440 ;
        RECT -3.865 -172.965 -3.695 -172.440 ;
        RECT -2.240 -172.855 -1.780 -172.685 ;
        RECT -10.245 -173.295 -9.695 -172.965 ;
        RECT -4.245 -173.295 -3.695 -172.965 ;
        RECT -10.245 -173.820 -10.075 -173.295 ;
        RECT -3.865 -173.820 -3.695 -173.295 ;
        RECT -2.155 -173.580 -1.865 -172.855 ;
        RECT -0.325 -172.965 -0.155 -172.440 ;
        RECT 6.055 -172.965 6.225 -172.440 ;
        RECT 7.680 -172.855 8.140 -172.685 ;
        RECT -0.325 -173.295 0.225 -172.965 ;
        RECT 5.675 -173.295 6.225 -172.965 ;
        RECT -0.325 -173.820 -0.155 -173.295 ;
        RECT 6.055 -173.820 6.225 -173.295 ;
        RECT 7.765 -173.580 8.055 -172.855 ;
        RECT 9.595 -172.965 9.765 -172.440 ;
        RECT 15.975 -172.965 16.145 -172.440 ;
        RECT 17.600 -172.855 18.060 -172.685 ;
        RECT 9.595 -173.295 10.145 -172.965 ;
        RECT 15.595 -173.295 16.145 -172.965 ;
        RECT 9.595 -173.820 9.765 -173.295 ;
        RECT 15.975 -173.820 16.145 -173.295 ;
        RECT 17.685 -173.580 17.975 -172.855 ;
        RECT 19.515 -172.965 19.685 -172.440 ;
        RECT 19.515 -173.295 20.065 -172.965 ;
        RECT 19.515 -173.820 19.685 -173.295 ;
        RECT -286.340 -174.335 -283.120 -174.165 ;
        RECT -276.420 -174.335 -273.200 -174.165 ;
        RECT -266.500 -174.335 -263.280 -174.165 ;
        RECT -256.580 -174.335 -253.360 -174.165 ;
        RECT -246.660 -174.335 -243.440 -174.165 ;
        RECT -236.740 -174.335 -233.520 -174.165 ;
        RECT -226.820 -174.335 -223.600 -174.165 ;
        RECT -216.900 -174.335 -213.680 -174.165 ;
        RECT -206.980 -174.335 -203.760 -174.165 ;
        RECT -197.060 -174.335 -193.840 -174.165 ;
        RECT -187.140 -174.335 -183.920 -174.165 ;
        RECT -177.220 -174.335 -174.000 -174.165 ;
        RECT -167.300 -174.335 -164.080 -174.165 ;
        RECT -157.380 -174.335 -154.160 -174.165 ;
        RECT -147.460 -174.335 -144.240 -174.165 ;
        RECT -137.540 -174.335 -134.320 -174.165 ;
        RECT -127.620 -174.335 -124.400 -174.165 ;
        RECT -117.700 -174.335 -114.480 -174.165 ;
        RECT -107.780 -174.335 -104.560 -174.165 ;
        RECT -97.860 -174.335 -94.640 -174.165 ;
        RECT -87.940 -174.335 -84.720 -174.165 ;
        RECT -78.020 -174.335 -74.800 -174.165 ;
        RECT -68.100 -174.335 -64.880 -174.165 ;
        RECT -58.180 -174.335 -54.960 -174.165 ;
        RECT -48.260 -174.335 -45.040 -174.165 ;
        RECT -38.340 -174.335 -35.120 -174.165 ;
        RECT -28.420 -174.335 -25.200 -174.165 ;
        RECT -18.500 -174.335 -15.280 -174.165 ;
        RECT -8.580 -174.335 -5.360 -174.165 ;
        RECT 1.340 -174.335 4.560 -174.165 ;
        RECT 11.260 -174.335 14.480 -174.165 ;
        RECT -285.355 -175.135 -285.045 -174.335 ;
        RECT -284.875 -175.060 -284.585 -174.335 ;
        RECT -284.415 -175.135 -284.105 -174.335 ;
        RECT -275.435 -175.135 -275.125 -174.335 ;
        RECT -274.955 -175.060 -274.665 -174.335 ;
        RECT -274.495 -175.135 -274.185 -174.335 ;
        RECT -265.515 -175.135 -265.205 -174.335 ;
        RECT -265.035 -175.060 -264.745 -174.335 ;
        RECT -264.575 -175.135 -264.265 -174.335 ;
        RECT -255.595 -175.135 -255.285 -174.335 ;
        RECT -255.115 -175.060 -254.825 -174.335 ;
        RECT -254.655 -175.135 -254.345 -174.335 ;
        RECT -245.675 -175.135 -245.365 -174.335 ;
        RECT -245.195 -175.060 -244.905 -174.335 ;
        RECT -244.735 -175.135 -244.425 -174.335 ;
        RECT -235.755 -175.135 -235.445 -174.335 ;
        RECT -235.275 -175.060 -234.985 -174.335 ;
        RECT -234.815 -175.135 -234.505 -174.335 ;
        RECT -225.835 -175.135 -225.525 -174.335 ;
        RECT -225.355 -175.060 -225.065 -174.335 ;
        RECT -224.895 -175.135 -224.585 -174.335 ;
        RECT -215.915 -175.135 -215.605 -174.335 ;
        RECT -215.435 -175.060 -215.145 -174.335 ;
        RECT -214.975 -175.135 -214.665 -174.335 ;
        RECT -205.995 -175.135 -205.685 -174.335 ;
        RECT -205.515 -175.060 -205.225 -174.335 ;
        RECT -205.055 -175.135 -204.745 -174.335 ;
        RECT -196.075 -175.135 -195.765 -174.335 ;
        RECT -195.595 -175.060 -195.305 -174.335 ;
        RECT -195.135 -175.135 -194.825 -174.335 ;
        RECT -186.155 -175.135 -185.845 -174.335 ;
        RECT -185.675 -175.060 -185.385 -174.335 ;
        RECT -185.215 -175.135 -184.905 -174.335 ;
        RECT -176.235 -175.135 -175.925 -174.335 ;
        RECT -175.755 -175.060 -175.465 -174.335 ;
        RECT -175.295 -175.135 -174.985 -174.335 ;
        RECT -166.315 -175.135 -166.005 -174.335 ;
        RECT -165.835 -175.060 -165.545 -174.335 ;
        RECT -165.375 -175.135 -165.065 -174.335 ;
        RECT -156.395 -175.135 -156.085 -174.335 ;
        RECT -155.915 -175.060 -155.625 -174.335 ;
        RECT -155.455 -175.135 -155.145 -174.335 ;
        RECT -146.475 -175.135 -146.165 -174.335 ;
        RECT -145.995 -175.060 -145.705 -174.335 ;
        RECT -145.535 -175.135 -145.225 -174.335 ;
        RECT -136.555 -175.135 -136.245 -174.335 ;
        RECT -136.075 -175.060 -135.785 -174.335 ;
        RECT -135.615 -175.135 -135.305 -174.335 ;
        RECT -126.635 -175.135 -126.325 -174.335 ;
        RECT -126.155 -175.060 -125.865 -174.335 ;
        RECT -125.695 -175.135 -125.385 -174.335 ;
        RECT -116.715 -175.135 -116.405 -174.335 ;
        RECT -116.235 -175.060 -115.945 -174.335 ;
        RECT -115.775 -175.135 -115.465 -174.335 ;
        RECT -106.795 -175.135 -106.485 -174.335 ;
        RECT -106.315 -175.060 -106.025 -174.335 ;
        RECT -105.855 -175.135 -105.545 -174.335 ;
        RECT -96.875 -175.135 -96.565 -174.335 ;
        RECT -96.395 -175.060 -96.105 -174.335 ;
        RECT -95.935 -175.135 -95.625 -174.335 ;
        RECT -86.955 -175.135 -86.645 -174.335 ;
        RECT -86.475 -175.060 -86.185 -174.335 ;
        RECT -86.015 -175.135 -85.705 -174.335 ;
        RECT -77.035 -175.135 -76.725 -174.335 ;
        RECT -76.555 -175.060 -76.265 -174.335 ;
        RECT -76.095 -175.135 -75.785 -174.335 ;
        RECT -67.115 -175.135 -66.805 -174.335 ;
        RECT -66.635 -175.060 -66.345 -174.335 ;
        RECT -66.175 -175.135 -65.865 -174.335 ;
        RECT -57.195 -175.135 -56.885 -174.335 ;
        RECT -56.715 -175.060 -56.425 -174.335 ;
        RECT -56.255 -175.135 -55.945 -174.335 ;
        RECT -47.275 -175.135 -46.965 -174.335 ;
        RECT -46.795 -175.060 -46.505 -174.335 ;
        RECT -46.335 -175.135 -46.025 -174.335 ;
        RECT -37.355 -175.135 -37.045 -174.335 ;
        RECT -36.875 -175.060 -36.585 -174.335 ;
        RECT -36.415 -175.135 -36.105 -174.335 ;
        RECT -27.435 -175.135 -27.125 -174.335 ;
        RECT -26.955 -175.060 -26.665 -174.335 ;
        RECT -26.495 -175.135 -26.185 -174.335 ;
        RECT -17.515 -175.135 -17.205 -174.335 ;
        RECT -17.035 -175.060 -16.745 -174.335 ;
        RECT -16.575 -175.135 -16.265 -174.335 ;
        RECT -7.595 -175.135 -7.285 -174.335 ;
        RECT -7.115 -175.060 -6.825 -174.335 ;
        RECT -6.655 -175.135 -6.345 -174.335 ;
        RECT 2.325 -175.135 2.635 -174.335 ;
        RECT 2.805 -175.060 3.095 -174.335 ;
        RECT 3.265 -175.135 3.575 -174.335 ;
        RECT 12.245 -175.135 12.555 -174.335 ;
        RECT 12.725 -175.060 13.015 -174.335 ;
        RECT 13.185 -175.135 13.495 -174.335 ;
        RECT -290.315 -176.885 -290.005 -176.085 ;
        RECT -289.835 -176.885 -289.545 -176.160 ;
        RECT -289.375 -176.885 -289.065 -176.085 ;
        RECT -280.395 -176.885 -280.085 -176.085 ;
        RECT -279.915 -176.885 -279.625 -176.160 ;
        RECT -279.455 -176.885 -279.145 -176.085 ;
        RECT -270.475 -176.885 -270.165 -176.085 ;
        RECT -269.995 -176.885 -269.705 -176.160 ;
        RECT -269.535 -176.885 -269.225 -176.085 ;
        RECT -260.555 -176.885 -260.245 -176.085 ;
        RECT -260.075 -176.885 -259.785 -176.160 ;
        RECT -259.615 -176.885 -259.305 -176.085 ;
        RECT -250.635 -176.885 -250.325 -176.085 ;
        RECT -250.155 -176.885 -249.865 -176.160 ;
        RECT -249.695 -176.885 -249.385 -176.085 ;
        RECT -240.715 -176.885 -240.405 -176.085 ;
        RECT -240.235 -176.885 -239.945 -176.160 ;
        RECT -239.775 -176.885 -239.465 -176.085 ;
        RECT -230.795 -176.885 -230.485 -176.085 ;
        RECT -230.315 -176.885 -230.025 -176.160 ;
        RECT -229.855 -176.885 -229.545 -176.085 ;
        RECT -220.875 -176.885 -220.565 -176.085 ;
        RECT -220.395 -176.885 -220.105 -176.160 ;
        RECT -219.935 -176.885 -219.625 -176.085 ;
        RECT -210.955 -176.885 -210.645 -176.085 ;
        RECT -210.475 -176.885 -210.185 -176.160 ;
        RECT -210.015 -176.885 -209.705 -176.085 ;
        RECT -201.035 -176.885 -200.725 -176.085 ;
        RECT -200.555 -176.885 -200.265 -176.160 ;
        RECT -200.095 -176.885 -199.785 -176.085 ;
        RECT -191.115 -176.885 -190.805 -176.085 ;
        RECT -190.635 -176.885 -190.345 -176.160 ;
        RECT -190.175 -176.885 -189.865 -176.085 ;
        RECT -181.195 -176.885 -180.885 -176.085 ;
        RECT -180.715 -176.885 -180.425 -176.160 ;
        RECT -180.255 -176.885 -179.945 -176.085 ;
        RECT -171.275 -176.885 -170.965 -176.085 ;
        RECT -170.795 -176.885 -170.505 -176.160 ;
        RECT -170.335 -176.885 -170.025 -176.085 ;
        RECT -161.355 -176.885 -161.045 -176.085 ;
        RECT -160.875 -176.885 -160.585 -176.160 ;
        RECT -160.415 -176.885 -160.105 -176.085 ;
        RECT -151.435 -176.885 -151.125 -176.085 ;
        RECT -150.955 -176.885 -150.665 -176.160 ;
        RECT -150.495 -176.885 -150.185 -176.085 ;
        RECT -141.515 -176.885 -141.205 -176.085 ;
        RECT -141.035 -176.885 -140.745 -176.160 ;
        RECT -140.575 -176.885 -140.265 -176.085 ;
        RECT -131.595 -176.885 -131.285 -176.085 ;
        RECT -131.115 -176.885 -130.825 -176.160 ;
        RECT -130.655 -176.885 -130.345 -176.085 ;
        RECT -121.675 -176.885 -121.365 -176.085 ;
        RECT -121.195 -176.885 -120.905 -176.160 ;
        RECT -120.735 -176.885 -120.425 -176.085 ;
        RECT -111.755 -176.885 -111.445 -176.085 ;
        RECT -111.275 -176.885 -110.985 -176.160 ;
        RECT -110.815 -176.885 -110.505 -176.085 ;
        RECT -101.835 -176.885 -101.525 -176.085 ;
        RECT -101.355 -176.885 -101.065 -176.160 ;
        RECT -100.895 -176.885 -100.585 -176.085 ;
        RECT -91.915 -176.885 -91.605 -176.085 ;
        RECT -91.435 -176.885 -91.145 -176.160 ;
        RECT -90.975 -176.885 -90.665 -176.085 ;
        RECT -81.995 -176.885 -81.685 -176.085 ;
        RECT -81.515 -176.885 -81.225 -176.160 ;
        RECT -81.055 -176.885 -80.745 -176.085 ;
        RECT -72.075 -176.885 -71.765 -176.085 ;
        RECT -71.595 -176.885 -71.305 -176.160 ;
        RECT -71.135 -176.885 -70.825 -176.085 ;
        RECT -62.155 -176.885 -61.845 -176.085 ;
        RECT -61.675 -176.885 -61.385 -176.160 ;
        RECT -61.215 -176.885 -60.905 -176.085 ;
        RECT -52.235 -176.885 -51.925 -176.085 ;
        RECT -51.755 -176.885 -51.465 -176.160 ;
        RECT -51.295 -176.885 -50.985 -176.085 ;
        RECT -42.315 -176.885 -42.005 -176.085 ;
        RECT -41.835 -176.885 -41.545 -176.160 ;
        RECT -41.375 -176.885 -41.065 -176.085 ;
        RECT -32.395 -176.885 -32.085 -176.085 ;
        RECT -31.915 -176.885 -31.625 -176.160 ;
        RECT -31.455 -176.885 -31.145 -176.085 ;
        RECT -22.475 -176.885 -22.165 -176.085 ;
        RECT -21.995 -176.885 -21.705 -176.160 ;
        RECT -21.535 -176.885 -21.225 -176.085 ;
        RECT -12.555 -176.885 -12.245 -176.085 ;
        RECT -12.075 -176.885 -11.785 -176.160 ;
        RECT -11.615 -176.885 -11.305 -176.085 ;
        RECT -2.635 -176.885 -2.325 -176.085 ;
        RECT -2.155 -176.885 -1.865 -176.160 ;
        RECT -1.695 -176.885 -1.385 -176.085 ;
        RECT 7.285 -176.885 7.595 -176.085 ;
        RECT 7.765 -176.885 8.055 -176.160 ;
        RECT 8.225 -176.885 8.535 -176.085 ;
        RECT 17.205 -176.885 17.515 -176.085 ;
        RECT 17.685 -176.885 17.975 -176.160 ;
        RECT 18.145 -176.885 18.455 -176.085 ;
        RECT -291.300 -177.055 -288.080 -176.885 ;
        RECT -281.380 -177.055 -278.160 -176.885 ;
        RECT -271.460 -177.055 -268.240 -176.885 ;
        RECT -261.540 -177.055 -258.320 -176.885 ;
        RECT -251.620 -177.055 -248.400 -176.885 ;
        RECT -241.700 -177.055 -238.480 -176.885 ;
        RECT -231.780 -177.055 -228.560 -176.885 ;
        RECT -221.860 -177.055 -218.640 -176.885 ;
        RECT -211.940 -177.055 -208.720 -176.885 ;
        RECT -202.020 -177.055 -198.800 -176.885 ;
        RECT -192.100 -177.055 -188.880 -176.885 ;
        RECT -182.180 -177.055 -178.960 -176.885 ;
        RECT -172.260 -177.055 -169.040 -176.885 ;
        RECT -162.340 -177.055 -159.120 -176.885 ;
        RECT -152.420 -177.055 -149.200 -176.885 ;
        RECT -142.500 -177.055 -139.280 -176.885 ;
        RECT -132.580 -177.055 -129.360 -176.885 ;
        RECT -122.660 -177.055 -119.440 -176.885 ;
        RECT -112.740 -177.055 -109.520 -176.885 ;
        RECT -102.820 -177.055 -99.600 -176.885 ;
        RECT -92.900 -177.055 -89.680 -176.885 ;
        RECT -82.980 -177.055 -79.760 -176.885 ;
        RECT -73.060 -177.055 -69.840 -176.885 ;
        RECT -63.140 -177.055 -59.920 -176.885 ;
        RECT -53.220 -177.055 -50.000 -176.885 ;
        RECT -43.300 -177.055 -40.080 -176.885 ;
        RECT -33.380 -177.055 -30.160 -176.885 ;
        RECT -23.460 -177.055 -20.240 -176.885 ;
        RECT -13.540 -177.055 -10.320 -176.885 ;
        RECT -3.620 -177.055 -0.400 -176.885 ;
        RECT 6.300 -177.055 9.520 -176.885 ;
        RECT 16.220 -177.055 19.440 -176.885 ;
        RECT -286.585 -177.925 -286.415 -177.400 ;
        RECT -286.965 -178.255 -286.415 -177.925 ;
        RECT -286.585 -178.780 -286.415 -178.255 ;
        RECT -284.875 -178.275 -284.585 -177.550 ;
        RECT -283.045 -177.925 -282.875 -177.400 ;
        RECT -276.665 -177.925 -276.495 -177.400 ;
        RECT -283.045 -178.255 -282.495 -177.925 ;
        RECT -277.045 -178.255 -276.495 -177.925 ;
        RECT -284.960 -178.445 -284.500 -178.275 ;
        RECT -283.045 -178.780 -282.875 -178.255 ;
        RECT -276.665 -178.780 -276.495 -178.255 ;
        RECT -274.955 -178.275 -274.665 -177.550 ;
        RECT -273.125 -177.925 -272.955 -177.400 ;
        RECT -266.745 -177.925 -266.575 -177.400 ;
        RECT -273.125 -178.255 -272.575 -177.925 ;
        RECT -267.125 -178.255 -266.575 -177.925 ;
        RECT -275.040 -178.445 -274.580 -178.275 ;
        RECT -273.125 -178.780 -272.955 -178.255 ;
        RECT -266.745 -178.780 -266.575 -178.255 ;
        RECT -265.035 -178.275 -264.745 -177.550 ;
        RECT -263.205 -177.925 -263.035 -177.400 ;
        RECT -256.825 -177.925 -256.655 -177.400 ;
        RECT -263.205 -178.255 -262.655 -177.925 ;
        RECT -257.205 -178.255 -256.655 -177.925 ;
        RECT -265.120 -178.445 -264.660 -178.275 ;
        RECT -263.205 -178.780 -263.035 -178.255 ;
        RECT -256.825 -178.780 -256.655 -178.255 ;
        RECT -255.115 -178.275 -254.825 -177.550 ;
        RECT -253.285 -177.925 -253.115 -177.400 ;
        RECT -246.905 -177.925 -246.735 -177.400 ;
        RECT -253.285 -178.255 -252.735 -177.925 ;
        RECT -247.285 -178.255 -246.735 -177.925 ;
        RECT -255.200 -178.445 -254.740 -178.275 ;
        RECT -253.285 -178.780 -253.115 -178.255 ;
        RECT -246.905 -178.780 -246.735 -178.255 ;
        RECT -245.195 -178.275 -244.905 -177.550 ;
        RECT -243.365 -177.925 -243.195 -177.400 ;
        RECT -236.985 -177.925 -236.815 -177.400 ;
        RECT -243.365 -178.255 -242.815 -177.925 ;
        RECT -237.365 -178.255 -236.815 -177.925 ;
        RECT -245.280 -178.445 -244.820 -178.275 ;
        RECT -243.365 -178.780 -243.195 -178.255 ;
        RECT -236.985 -178.780 -236.815 -178.255 ;
        RECT -235.275 -178.275 -234.985 -177.550 ;
        RECT -233.445 -177.925 -233.275 -177.400 ;
        RECT -227.065 -177.925 -226.895 -177.400 ;
        RECT -233.445 -178.255 -232.895 -177.925 ;
        RECT -227.445 -178.255 -226.895 -177.925 ;
        RECT -235.360 -178.445 -234.900 -178.275 ;
        RECT -233.445 -178.780 -233.275 -178.255 ;
        RECT -227.065 -178.780 -226.895 -178.255 ;
        RECT -225.355 -178.275 -225.065 -177.550 ;
        RECT -223.525 -177.925 -223.355 -177.400 ;
        RECT -217.145 -177.925 -216.975 -177.400 ;
        RECT -223.525 -178.255 -222.975 -177.925 ;
        RECT -217.525 -178.255 -216.975 -177.925 ;
        RECT -225.440 -178.445 -224.980 -178.275 ;
        RECT -223.525 -178.780 -223.355 -178.255 ;
        RECT -217.145 -178.780 -216.975 -178.255 ;
        RECT -215.435 -178.275 -215.145 -177.550 ;
        RECT -213.605 -177.925 -213.435 -177.400 ;
        RECT -207.225 -177.925 -207.055 -177.400 ;
        RECT -213.605 -178.255 -213.055 -177.925 ;
        RECT -207.605 -178.255 -207.055 -177.925 ;
        RECT -215.520 -178.445 -215.060 -178.275 ;
        RECT -213.605 -178.780 -213.435 -178.255 ;
        RECT -207.225 -178.780 -207.055 -178.255 ;
        RECT -205.515 -178.275 -205.225 -177.550 ;
        RECT -203.685 -177.925 -203.515 -177.400 ;
        RECT -197.305 -177.925 -197.135 -177.400 ;
        RECT -203.685 -178.255 -203.135 -177.925 ;
        RECT -197.685 -178.255 -197.135 -177.925 ;
        RECT -205.600 -178.445 -205.140 -178.275 ;
        RECT -203.685 -178.780 -203.515 -178.255 ;
        RECT -197.305 -178.780 -197.135 -178.255 ;
        RECT -195.595 -178.275 -195.305 -177.550 ;
        RECT -193.765 -177.925 -193.595 -177.400 ;
        RECT -187.385 -177.925 -187.215 -177.400 ;
        RECT -193.765 -178.255 -193.215 -177.925 ;
        RECT -187.765 -178.255 -187.215 -177.925 ;
        RECT -195.680 -178.445 -195.220 -178.275 ;
        RECT -193.765 -178.780 -193.595 -178.255 ;
        RECT -187.385 -178.780 -187.215 -178.255 ;
        RECT -185.675 -178.275 -185.385 -177.550 ;
        RECT -183.845 -177.925 -183.675 -177.400 ;
        RECT -177.465 -177.925 -177.295 -177.400 ;
        RECT -183.845 -178.255 -183.295 -177.925 ;
        RECT -177.845 -178.255 -177.295 -177.925 ;
        RECT -185.760 -178.445 -185.300 -178.275 ;
        RECT -183.845 -178.780 -183.675 -178.255 ;
        RECT -177.465 -178.780 -177.295 -178.255 ;
        RECT -175.755 -178.275 -175.465 -177.550 ;
        RECT -173.925 -177.925 -173.755 -177.400 ;
        RECT -167.545 -177.925 -167.375 -177.400 ;
        RECT -173.925 -178.255 -173.375 -177.925 ;
        RECT -167.925 -178.255 -167.375 -177.925 ;
        RECT -175.840 -178.445 -175.380 -178.275 ;
        RECT -173.925 -178.780 -173.755 -178.255 ;
        RECT -167.545 -178.780 -167.375 -178.255 ;
        RECT -165.835 -178.275 -165.545 -177.550 ;
        RECT -164.005 -177.925 -163.835 -177.400 ;
        RECT -157.625 -177.925 -157.455 -177.400 ;
        RECT -164.005 -178.255 -163.455 -177.925 ;
        RECT -158.005 -178.255 -157.455 -177.925 ;
        RECT -165.920 -178.445 -165.460 -178.275 ;
        RECT -164.005 -178.780 -163.835 -178.255 ;
        RECT -157.625 -178.780 -157.455 -178.255 ;
        RECT -155.915 -178.275 -155.625 -177.550 ;
        RECT -154.085 -177.925 -153.915 -177.400 ;
        RECT -147.705 -177.925 -147.535 -177.400 ;
        RECT -154.085 -178.255 -153.535 -177.925 ;
        RECT -148.085 -178.255 -147.535 -177.925 ;
        RECT -156.000 -178.445 -155.540 -178.275 ;
        RECT -154.085 -178.780 -153.915 -178.255 ;
        RECT -147.705 -178.780 -147.535 -178.255 ;
        RECT -145.995 -178.275 -145.705 -177.550 ;
        RECT -144.165 -177.925 -143.995 -177.400 ;
        RECT -137.785 -177.925 -137.615 -177.400 ;
        RECT -144.165 -178.255 -143.615 -177.925 ;
        RECT -138.165 -178.255 -137.615 -177.925 ;
        RECT -146.080 -178.445 -145.620 -178.275 ;
        RECT -144.165 -178.780 -143.995 -178.255 ;
        RECT -137.785 -178.780 -137.615 -178.255 ;
        RECT -136.075 -178.275 -135.785 -177.550 ;
        RECT -134.245 -177.925 -134.075 -177.400 ;
        RECT -127.865 -177.925 -127.695 -177.400 ;
        RECT -134.245 -178.255 -133.695 -177.925 ;
        RECT -128.245 -178.255 -127.695 -177.925 ;
        RECT -136.160 -178.445 -135.700 -178.275 ;
        RECT -134.245 -178.780 -134.075 -178.255 ;
        RECT -127.865 -178.780 -127.695 -178.255 ;
        RECT -126.155 -178.275 -125.865 -177.550 ;
        RECT -124.325 -177.925 -124.155 -177.400 ;
        RECT -117.945 -177.925 -117.775 -177.400 ;
        RECT -124.325 -178.255 -123.775 -177.925 ;
        RECT -118.325 -178.255 -117.775 -177.925 ;
        RECT -126.240 -178.445 -125.780 -178.275 ;
        RECT -124.325 -178.780 -124.155 -178.255 ;
        RECT -117.945 -178.780 -117.775 -178.255 ;
        RECT -116.235 -178.275 -115.945 -177.550 ;
        RECT -114.405 -177.925 -114.235 -177.400 ;
        RECT -108.025 -177.925 -107.855 -177.400 ;
        RECT -114.405 -178.255 -113.855 -177.925 ;
        RECT -108.405 -178.255 -107.855 -177.925 ;
        RECT -116.320 -178.445 -115.860 -178.275 ;
        RECT -114.405 -178.780 -114.235 -178.255 ;
        RECT -108.025 -178.780 -107.855 -178.255 ;
        RECT -106.315 -178.275 -106.025 -177.550 ;
        RECT -104.485 -177.925 -104.315 -177.400 ;
        RECT -98.105 -177.925 -97.935 -177.400 ;
        RECT -104.485 -178.255 -103.935 -177.925 ;
        RECT -98.485 -178.255 -97.935 -177.925 ;
        RECT -106.400 -178.445 -105.940 -178.275 ;
        RECT -104.485 -178.780 -104.315 -178.255 ;
        RECT -98.105 -178.780 -97.935 -178.255 ;
        RECT -96.395 -178.275 -96.105 -177.550 ;
        RECT -94.565 -177.925 -94.395 -177.400 ;
        RECT -88.185 -177.925 -88.015 -177.400 ;
        RECT -94.565 -178.255 -94.015 -177.925 ;
        RECT -88.565 -178.255 -88.015 -177.925 ;
        RECT -96.480 -178.445 -96.020 -178.275 ;
        RECT -94.565 -178.780 -94.395 -178.255 ;
        RECT -88.185 -178.780 -88.015 -178.255 ;
        RECT -86.475 -178.275 -86.185 -177.550 ;
        RECT -84.645 -177.925 -84.475 -177.400 ;
        RECT -78.265 -177.925 -78.095 -177.400 ;
        RECT -84.645 -178.255 -84.095 -177.925 ;
        RECT -78.645 -178.255 -78.095 -177.925 ;
        RECT -86.560 -178.445 -86.100 -178.275 ;
        RECT -84.645 -178.780 -84.475 -178.255 ;
        RECT -78.265 -178.780 -78.095 -178.255 ;
        RECT -76.555 -178.275 -76.265 -177.550 ;
        RECT -74.725 -177.925 -74.555 -177.400 ;
        RECT -68.345 -177.925 -68.175 -177.400 ;
        RECT -74.725 -178.255 -74.175 -177.925 ;
        RECT -68.725 -178.255 -68.175 -177.925 ;
        RECT -76.640 -178.445 -76.180 -178.275 ;
        RECT -74.725 -178.780 -74.555 -178.255 ;
        RECT -68.345 -178.780 -68.175 -178.255 ;
        RECT -66.635 -178.275 -66.345 -177.550 ;
        RECT -64.805 -177.925 -64.635 -177.400 ;
        RECT -58.425 -177.925 -58.255 -177.400 ;
        RECT -64.805 -178.255 -64.255 -177.925 ;
        RECT -58.805 -178.255 -58.255 -177.925 ;
        RECT -66.720 -178.445 -66.260 -178.275 ;
        RECT -64.805 -178.780 -64.635 -178.255 ;
        RECT -58.425 -178.780 -58.255 -178.255 ;
        RECT -56.715 -178.275 -56.425 -177.550 ;
        RECT -54.885 -177.925 -54.715 -177.400 ;
        RECT -48.505 -177.925 -48.335 -177.400 ;
        RECT -54.885 -178.255 -54.335 -177.925 ;
        RECT -48.885 -178.255 -48.335 -177.925 ;
        RECT -56.800 -178.445 -56.340 -178.275 ;
        RECT -54.885 -178.780 -54.715 -178.255 ;
        RECT -48.505 -178.780 -48.335 -178.255 ;
        RECT -46.795 -178.275 -46.505 -177.550 ;
        RECT -44.965 -177.925 -44.795 -177.400 ;
        RECT -38.585 -177.925 -38.415 -177.400 ;
        RECT -44.965 -178.255 -44.415 -177.925 ;
        RECT -38.965 -178.255 -38.415 -177.925 ;
        RECT -46.880 -178.445 -46.420 -178.275 ;
        RECT -44.965 -178.780 -44.795 -178.255 ;
        RECT -38.585 -178.780 -38.415 -178.255 ;
        RECT -36.875 -178.275 -36.585 -177.550 ;
        RECT -35.045 -177.925 -34.875 -177.400 ;
        RECT -28.665 -177.925 -28.495 -177.400 ;
        RECT -35.045 -178.255 -34.495 -177.925 ;
        RECT -29.045 -178.255 -28.495 -177.925 ;
        RECT -36.960 -178.445 -36.500 -178.275 ;
        RECT -35.045 -178.780 -34.875 -178.255 ;
        RECT -28.665 -178.780 -28.495 -178.255 ;
        RECT -26.955 -178.275 -26.665 -177.550 ;
        RECT -25.125 -177.925 -24.955 -177.400 ;
        RECT -18.745 -177.925 -18.575 -177.400 ;
        RECT -25.125 -178.255 -24.575 -177.925 ;
        RECT -19.125 -178.255 -18.575 -177.925 ;
        RECT -27.040 -178.445 -26.580 -178.275 ;
        RECT -25.125 -178.780 -24.955 -178.255 ;
        RECT -18.745 -178.780 -18.575 -178.255 ;
        RECT -17.035 -178.275 -16.745 -177.550 ;
        RECT -15.205 -177.925 -15.035 -177.400 ;
        RECT -8.825 -177.925 -8.655 -177.400 ;
        RECT -15.205 -178.255 -14.655 -177.925 ;
        RECT -9.205 -178.255 -8.655 -177.925 ;
        RECT -17.120 -178.445 -16.660 -178.275 ;
        RECT -15.205 -178.780 -15.035 -178.255 ;
        RECT -8.825 -178.780 -8.655 -178.255 ;
        RECT -7.115 -178.275 -6.825 -177.550 ;
        RECT -5.285 -177.925 -5.115 -177.400 ;
        RECT 1.095 -177.925 1.265 -177.400 ;
        RECT -5.285 -178.255 -4.735 -177.925 ;
        RECT 0.715 -178.255 1.265 -177.925 ;
        RECT -7.200 -178.445 -6.740 -178.275 ;
        RECT -5.285 -178.780 -5.115 -178.255 ;
        RECT 1.095 -178.780 1.265 -178.255 ;
        RECT 2.805 -178.275 3.095 -177.550 ;
        RECT 4.635 -177.925 4.805 -177.400 ;
        RECT 11.015 -177.925 11.185 -177.400 ;
        RECT 4.635 -178.255 5.185 -177.925 ;
        RECT 10.635 -178.255 11.185 -177.925 ;
        RECT 2.720 -178.445 3.180 -178.275 ;
        RECT 4.635 -178.780 4.805 -178.255 ;
        RECT 11.015 -178.780 11.185 -178.255 ;
        RECT 12.725 -178.275 13.015 -177.550 ;
        RECT 14.555 -177.925 14.725 -177.400 ;
        RECT 14.555 -178.255 15.105 -177.925 ;
        RECT 12.640 -178.445 13.100 -178.275 ;
        RECT 14.555 -178.780 14.725 -178.255 ;
      LAYER mcon ;
        RECT -288.125 94.825 -287.955 94.995 ;
        RECT -286.355 94.725 -286.185 94.895 ;
        RECT -284.585 94.825 -284.415 94.995 ;
        RECT -288.125 94.365 -287.955 94.535 ;
        RECT -288.125 93.905 -287.955 94.075 ;
        RECT -278.205 94.825 -278.035 94.995 ;
        RECT -276.435 94.725 -276.265 94.895 ;
        RECT -274.665 94.825 -274.495 94.995 ;
        RECT -284.585 94.365 -284.415 94.535 ;
        RECT -278.205 94.365 -278.035 94.535 ;
        RECT -284.585 93.905 -284.415 94.075 ;
        RECT -278.205 93.905 -278.035 94.075 ;
        RECT -268.285 94.825 -268.115 94.995 ;
        RECT -266.515 94.725 -266.345 94.895 ;
        RECT -264.745 94.825 -264.575 94.995 ;
        RECT -274.665 94.365 -274.495 94.535 ;
        RECT -268.285 94.365 -268.115 94.535 ;
        RECT -274.665 93.905 -274.495 94.075 ;
        RECT -268.285 93.905 -268.115 94.075 ;
        RECT -258.365 94.825 -258.195 94.995 ;
        RECT -256.595 94.725 -256.425 94.895 ;
        RECT -254.825 94.825 -254.655 94.995 ;
        RECT -264.745 94.365 -264.575 94.535 ;
        RECT -258.365 94.365 -258.195 94.535 ;
        RECT -264.745 93.905 -264.575 94.075 ;
        RECT -258.365 93.905 -258.195 94.075 ;
        RECT -248.445 94.825 -248.275 94.995 ;
        RECT -246.675 94.725 -246.505 94.895 ;
        RECT -244.905 94.825 -244.735 94.995 ;
        RECT -254.825 94.365 -254.655 94.535 ;
        RECT -248.445 94.365 -248.275 94.535 ;
        RECT -254.825 93.905 -254.655 94.075 ;
        RECT -248.445 93.905 -248.275 94.075 ;
        RECT -238.525 94.825 -238.355 94.995 ;
        RECT -236.755 94.725 -236.585 94.895 ;
        RECT -234.985 94.825 -234.815 94.995 ;
        RECT -244.905 94.365 -244.735 94.535 ;
        RECT -238.525 94.365 -238.355 94.535 ;
        RECT -244.905 93.905 -244.735 94.075 ;
        RECT -238.525 93.905 -238.355 94.075 ;
        RECT -228.605 94.825 -228.435 94.995 ;
        RECT -226.835 94.725 -226.665 94.895 ;
        RECT -225.065 94.825 -224.895 94.995 ;
        RECT -234.985 94.365 -234.815 94.535 ;
        RECT -228.605 94.365 -228.435 94.535 ;
        RECT -234.985 93.905 -234.815 94.075 ;
        RECT -228.605 93.905 -228.435 94.075 ;
        RECT -218.685 94.825 -218.515 94.995 ;
        RECT -216.915 94.725 -216.745 94.895 ;
        RECT -215.145 94.825 -214.975 94.995 ;
        RECT -225.065 94.365 -224.895 94.535 ;
        RECT -218.685 94.365 -218.515 94.535 ;
        RECT -225.065 93.905 -224.895 94.075 ;
        RECT -218.685 93.905 -218.515 94.075 ;
        RECT -208.765 94.825 -208.595 94.995 ;
        RECT -206.995 94.725 -206.825 94.895 ;
        RECT -205.225 94.825 -205.055 94.995 ;
        RECT -215.145 94.365 -214.975 94.535 ;
        RECT -208.765 94.365 -208.595 94.535 ;
        RECT -215.145 93.905 -214.975 94.075 ;
        RECT -208.765 93.905 -208.595 94.075 ;
        RECT -198.845 94.825 -198.675 94.995 ;
        RECT -197.075 94.725 -196.905 94.895 ;
        RECT -195.305 94.825 -195.135 94.995 ;
        RECT -205.225 94.365 -205.055 94.535 ;
        RECT -198.845 94.365 -198.675 94.535 ;
        RECT -205.225 93.905 -205.055 94.075 ;
        RECT -198.845 93.905 -198.675 94.075 ;
        RECT -188.925 94.825 -188.755 94.995 ;
        RECT -187.155 94.725 -186.985 94.895 ;
        RECT -185.385 94.825 -185.215 94.995 ;
        RECT -195.305 94.365 -195.135 94.535 ;
        RECT -188.925 94.365 -188.755 94.535 ;
        RECT -195.305 93.905 -195.135 94.075 ;
        RECT -188.925 93.905 -188.755 94.075 ;
        RECT -179.005 94.825 -178.835 94.995 ;
        RECT -177.235 94.725 -177.065 94.895 ;
        RECT -175.465 94.825 -175.295 94.995 ;
        RECT -185.385 94.365 -185.215 94.535 ;
        RECT -179.005 94.365 -178.835 94.535 ;
        RECT -185.385 93.905 -185.215 94.075 ;
        RECT -179.005 93.905 -178.835 94.075 ;
        RECT -169.085 94.825 -168.915 94.995 ;
        RECT -167.315 94.725 -167.145 94.895 ;
        RECT -165.545 94.825 -165.375 94.995 ;
        RECT -175.465 94.365 -175.295 94.535 ;
        RECT -169.085 94.365 -168.915 94.535 ;
        RECT -175.465 93.905 -175.295 94.075 ;
        RECT -169.085 93.905 -168.915 94.075 ;
        RECT -159.165 94.825 -158.995 94.995 ;
        RECT -157.395 94.725 -157.225 94.895 ;
        RECT -155.625 94.825 -155.455 94.995 ;
        RECT -165.545 94.365 -165.375 94.535 ;
        RECT -159.165 94.365 -158.995 94.535 ;
        RECT -165.545 93.905 -165.375 94.075 ;
        RECT -159.165 93.905 -158.995 94.075 ;
        RECT -149.245 94.825 -149.075 94.995 ;
        RECT -147.475 94.725 -147.305 94.895 ;
        RECT -145.705 94.825 -145.535 94.995 ;
        RECT -155.625 94.365 -155.455 94.535 ;
        RECT -149.245 94.365 -149.075 94.535 ;
        RECT -155.625 93.905 -155.455 94.075 ;
        RECT -149.245 93.905 -149.075 94.075 ;
        RECT -139.325 94.825 -139.155 94.995 ;
        RECT -137.555 94.725 -137.385 94.895 ;
        RECT -135.785 94.825 -135.615 94.995 ;
        RECT -145.705 94.365 -145.535 94.535 ;
        RECT -139.325 94.365 -139.155 94.535 ;
        RECT -145.705 93.905 -145.535 94.075 ;
        RECT -139.325 93.905 -139.155 94.075 ;
        RECT -129.405 94.825 -129.235 94.995 ;
        RECT -127.635 94.725 -127.465 94.895 ;
        RECT -125.865 94.825 -125.695 94.995 ;
        RECT -135.785 94.365 -135.615 94.535 ;
        RECT -129.405 94.365 -129.235 94.535 ;
        RECT -135.785 93.905 -135.615 94.075 ;
        RECT -129.405 93.905 -129.235 94.075 ;
        RECT -119.485 94.825 -119.315 94.995 ;
        RECT -117.715 94.725 -117.545 94.895 ;
        RECT -115.945 94.825 -115.775 94.995 ;
        RECT -125.865 94.365 -125.695 94.535 ;
        RECT -119.485 94.365 -119.315 94.535 ;
        RECT -125.865 93.905 -125.695 94.075 ;
        RECT -119.485 93.905 -119.315 94.075 ;
        RECT -109.565 94.825 -109.395 94.995 ;
        RECT -107.795 94.725 -107.625 94.895 ;
        RECT -106.025 94.825 -105.855 94.995 ;
        RECT -115.945 94.365 -115.775 94.535 ;
        RECT -109.565 94.365 -109.395 94.535 ;
        RECT -115.945 93.905 -115.775 94.075 ;
        RECT -109.565 93.905 -109.395 94.075 ;
        RECT -99.645 94.825 -99.475 94.995 ;
        RECT -97.875 94.725 -97.705 94.895 ;
        RECT -96.105 94.825 -95.935 94.995 ;
        RECT -106.025 94.365 -105.855 94.535 ;
        RECT -99.645 94.365 -99.475 94.535 ;
        RECT -106.025 93.905 -105.855 94.075 ;
        RECT -99.645 93.905 -99.475 94.075 ;
        RECT -89.725 94.825 -89.555 94.995 ;
        RECT -87.955 94.725 -87.785 94.895 ;
        RECT -86.185 94.825 -86.015 94.995 ;
        RECT -96.105 94.365 -95.935 94.535 ;
        RECT -89.725 94.365 -89.555 94.535 ;
        RECT -96.105 93.905 -95.935 94.075 ;
        RECT -89.725 93.905 -89.555 94.075 ;
        RECT -79.805 94.825 -79.635 94.995 ;
        RECT -78.035 94.725 -77.865 94.895 ;
        RECT -76.265 94.825 -76.095 94.995 ;
        RECT -86.185 94.365 -86.015 94.535 ;
        RECT -79.805 94.365 -79.635 94.535 ;
        RECT -86.185 93.905 -86.015 94.075 ;
        RECT -79.805 93.905 -79.635 94.075 ;
        RECT -69.885 94.825 -69.715 94.995 ;
        RECT -68.115 94.725 -67.945 94.895 ;
        RECT -66.345 94.825 -66.175 94.995 ;
        RECT -76.265 94.365 -76.095 94.535 ;
        RECT -69.885 94.365 -69.715 94.535 ;
        RECT -76.265 93.905 -76.095 94.075 ;
        RECT -69.885 93.905 -69.715 94.075 ;
        RECT -59.965 94.825 -59.795 94.995 ;
        RECT -58.195 94.725 -58.025 94.895 ;
        RECT -56.425 94.825 -56.255 94.995 ;
        RECT -66.345 94.365 -66.175 94.535 ;
        RECT -59.965 94.365 -59.795 94.535 ;
        RECT -66.345 93.905 -66.175 94.075 ;
        RECT -59.965 93.905 -59.795 94.075 ;
        RECT -50.045 94.825 -49.875 94.995 ;
        RECT -48.275 94.725 -48.105 94.895 ;
        RECT -46.505 94.825 -46.335 94.995 ;
        RECT -56.425 94.365 -56.255 94.535 ;
        RECT -50.045 94.365 -49.875 94.535 ;
        RECT -56.425 93.905 -56.255 94.075 ;
        RECT -50.045 93.905 -49.875 94.075 ;
        RECT -40.125 94.825 -39.955 94.995 ;
        RECT -38.355 94.725 -38.185 94.895 ;
        RECT -36.585 94.825 -36.415 94.995 ;
        RECT -46.505 94.365 -46.335 94.535 ;
        RECT -40.125 94.365 -39.955 94.535 ;
        RECT -46.505 93.905 -46.335 94.075 ;
        RECT -40.125 93.905 -39.955 94.075 ;
        RECT -30.205 94.825 -30.035 94.995 ;
        RECT -28.435 94.725 -28.265 94.895 ;
        RECT -26.665 94.825 -26.495 94.995 ;
        RECT -36.585 94.365 -36.415 94.535 ;
        RECT -30.205 94.365 -30.035 94.535 ;
        RECT -36.585 93.905 -36.415 94.075 ;
        RECT -30.205 93.905 -30.035 94.075 ;
        RECT -20.285 94.825 -20.115 94.995 ;
        RECT -18.515 94.725 -18.345 94.895 ;
        RECT -16.745 94.825 -16.575 94.995 ;
        RECT -26.665 94.365 -26.495 94.535 ;
        RECT -20.285 94.365 -20.115 94.535 ;
        RECT -26.665 93.905 -26.495 94.075 ;
        RECT -20.285 93.905 -20.115 94.075 ;
        RECT -10.365 94.825 -10.195 94.995 ;
        RECT -8.595 94.725 -8.425 94.895 ;
        RECT -6.825 94.825 -6.655 94.995 ;
        RECT -16.745 94.365 -16.575 94.535 ;
        RECT -10.365 94.365 -10.195 94.535 ;
        RECT -16.745 93.905 -16.575 94.075 ;
        RECT -10.365 93.905 -10.195 94.075 ;
        RECT -0.445 94.825 -0.275 94.995 ;
        RECT 1.325 94.725 1.495 94.895 ;
        RECT 3.095 94.825 3.265 94.995 ;
        RECT -6.825 94.365 -6.655 94.535 ;
        RECT -0.445 94.365 -0.275 94.535 ;
        RECT -6.825 93.905 -6.655 94.075 ;
        RECT -0.445 93.905 -0.275 94.075 ;
        RECT 9.475 94.825 9.645 94.995 ;
        RECT 11.245 94.725 11.415 94.895 ;
        RECT 13.015 94.825 13.185 94.995 ;
        RECT 3.095 94.365 3.265 94.535 ;
        RECT 9.475 94.365 9.645 94.535 ;
        RECT 3.095 93.905 3.265 94.075 ;
        RECT 9.475 93.905 9.645 94.075 ;
        RECT 19.395 94.825 19.565 94.995 ;
        RECT 21.165 94.725 21.335 94.895 ;
        RECT 22.935 94.825 23.105 94.995 ;
        RECT 13.015 94.365 13.185 94.535 ;
        RECT 19.395 94.365 19.565 94.535 ;
        RECT 13.015 93.905 13.185 94.075 ;
        RECT 19.395 93.905 19.565 94.075 ;
        RECT 22.935 94.365 23.105 94.535 ;
        RECT 22.935 93.905 23.105 94.075 ;
        RECT -282.775 93.245 -282.605 93.415 ;
        RECT -282.315 93.245 -282.145 93.415 ;
        RECT -281.855 93.245 -281.685 93.415 ;
        RECT -281.395 93.245 -281.225 93.415 ;
        RECT -280.935 93.245 -280.765 93.415 ;
        RECT -280.475 93.245 -280.305 93.415 ;
        RECT -280.015 93.245 -279.845 93.415 ;
        RECT -272.855 93.245 -272.685 93.415 ;
        RECT -272.395 93.245 -272.225 93.415 ;
        RECT -271.935 93.245 -271.765 93.415 ;
        RECT -271.475 93.245 -271.305 93.415 ;
        RECT -271.015 93.245 -270.845 93.415 ;
        RECT -270.555 93.245 -270.385 93.415 ;
        RECT -270.095 93.245 -269.925 93.415 ;
        RECT -262.935 93.245 -262.765 93.415 ;
        RECT -262.475 93.245 -262.305 93.415 ;
        RECT -262.015 93.245 -261.845 93.415 ;
        RECT -261.555 93.245 -261.385 93.415 ;
        RECT -261.095 93.245 -260.925 93.415 ;
        RECT -260.635 93.245 -260.465 93.415 ;
        RECT -260.175 93.245 -260.005 93.415 ;
        RECT -253.015 93.245 -252.845 93.415 ;
        RECT -252.555 93.245 -252.385 93.415 ;
        RECT -252.095 93.245 -251.925 93.415 ;
        RECT -251.635 93.245 -251.465 93.415 ;
        RECT -251.175 93.245 -251.005 93.415 ;
        RECT -250.715 93.245 -250.545 93.415 ;
        RECT -250.255 93.245 -250.085 93.415 ;
        RECT -243.095 93.245 -242.925 93.415 ;
        RECT -242.635 93.245 -242.465 93.415 ;
        RECT -242.175 93.245 -242.005 93.415 ;
        RECT -241.715 93.245 -241.545 93.415 ;
        RECT -241.255 93.245 -241.085 93.415 ;
        RECT -240.795 93.245 -240.625 93.415 ;
        RECT -240.335 93.245 -240.165 93.415 ;
        RECT -233.175 93.245 -233.005 93.415 ;
        RECT -232.715 93.245 -232.545 93.415 ;
        RECT -232.255 93.245 -232.085 93.415 ;
        RECT -231.795 93.245 -231.625 93.415 ;
        RECT -231.335 93.245 -231.165 93.415 ;
        RECT -230.875 93.245 -230.705 93.415 ;
        RECT -230.415 93.245 -230.245 93.415 ;
        RECT -223.255 93.245 -223.085 93.415 ;
        RECT -222.795 93.245 -222.625 93.415 ;
        RECT -222.335 93.245 -222.165 93.415 ;
        RECT -221.875 93.245 -221.705 93.415 ;
        RECT -221.415 93.245 -221.245 93.415 ;
        RECT -220.955 93.245 -220.785 93.415 ;
        RECT -220.495 93.245 -220.325 93.415 ;
        RECT -213.335 93.245 -213.165 93.415 ;
        RECT -212.875 93.245 -212.705 93.415 ;
        RECT -212.415 93.245 -212.245 93.415 ;
        RECT -211.955 93.245 -211.785 93.415 ;
        RECT -211.495 93.245 -211.325 93.415 ;
        RECT -211.035 93.245 -210.865 93.415 ;
        RECT -210.575 93.245 -210.405 93.415 ;
        RECT -203.415 93.245 -203.245 93.415 ;
        RECT -202.955 93.245 -202.785 93.415 ;
        RECT -202.495 93.245 -202.325 93.415 ;
        RECT -202.035 93.245 -201.865 93.415 ;
        RECT -201.575 93.245 -201.405 93.415 ;
        RECT -201.115 93.245 -200.945 93.415 ;
        RECT -200.655 93.245 -200.485 93.415 ;
        RECT -193.495 93.245 -193.325 93.415 ;
        RECT -193.035 93.245 -192.865 93.415 ;
        RECT -192.575 93.245 -192.405 93.415 ;
        RECT -192.115 93.245 -191.945 93.415 ;
        RECT -191.655 93.245 -191.485 93.415 ;
        RECT -191.195 93.245 -191.025 93.415 ;
        RECT -190.735 93.245 -190.565 93.415 ;
        RECT -183.575 93.245 -183.405 93.415 ;
        RECT -183.115 93.245 -182.945 93.415 ;
        RECT -182.655 93.245 -182.485 93.415 ;
        RECT -182.195 93.245 -182.025 93.415 ;
        RECT -181.735 93.245 -181.565 93.415 ;
        RECT -181.275 93.245 -181.105 93.415 ;
        RECT -180.815 93.245 -180.645 93.415 ;
        RECT -173.655 93.245 -173.485 93.415 ;
        RECT -173.195 93.245 -173.025 93.415 ;
        RECT -172.735 93.245 -172.565 93.415 ;
        RECT -172.275 93.245 -172.105 93.415 ;
        RECT -171.815 93.245 -171.645 93.415 ;
        RECT -171.355 93.245 -171.185 93.415 ;
        RECT -170.895 93.245 -170.725 93.415 ;
        RECT -163.735 93.245 -163.565 93.415 ;
        RECT -163.275 93.245 -163.105 93.415 ;
        RECT -162.815 93.245 -162.645 93.415 ;
        RECT -162.355 93.245 -162.185 93.415 ;
        RECT -161.895 93.245 -161.725 93.415 ;
        RECT -161.435 93.245 -161.265 93.415 ;
        RECT -160.975 93.245 -160.805 93.415 ;
        RECT -153.815 93.245 -153.645 93.415 ;
        RECT -153.355 93.245 -153.185 93.415 ;
        RECT -152.895 93.245 -152.725 93.415 ;
        RECT -152.435 93.245 -152.265 93.415 ;
        RECT -151.975 93.245 -151.805 93.415 ;
        RECT -151.515 93.245 -151.345 93.415 ;
        RECT -151.055 93.245 -150.885 93.415 ;
        RECT -143.895 93.245 -143.725 93.415 ;
        RECT -143.435 93.245 -143.265 93.415 ;
        RECT -142.975 93.245 -142.805 93.415 ;
        RECT -142.515 93.245 -142.345 93.415 ;
        RECT -142.055 93.245 -141.885 93.415 ;
        RECT -141.595 93.245 -141.425 93.415 ;
        RECT -141.135 93.245 -140.965 93.415 ;
        RECT -133.975 93.245 -133.805 93.415 ;
        RECT -133.515 93.245 -133.345 93.415 ;
        RECT -133.055 93.245 -132.885 93.415 ;
        RECT -132.595 93.245 -132.425 93.415 ;
        RECT -132.135 93.245 -131.965 93.415 ;
        RECT -131.675 93.245 -131.505 93.415 ;
        RECT -131.215 93.245 -131.045 93.415 ;
        RECT -124.055 93.245 -123.885 93.415 ;
        RECT -123.595 93.245 -123.425 93.415 ;
        RECT -123.135 93.245 -122.965 93.415 ;
        RECT -122.675 93.245 -122.505 93.415 ;
        RECT -122.215 93.245 -122.045 93.415 ;
        RECT -121.755 93.245 -121.585 93.415 ;
        RECT -121.295 93.245 -121.125 93.415 ;
        RECT -114.135 93.245 -113.965 93.415 ;
        RECT -113.675 93.245 -113.505 93.415 ;
        RECT -113.215 93.245 -113.045 93.415 ;
        RECT -112.755 93.245 -112.585 93.415 ;
        RECT -112.295 93.245 -112.125 93.415 ;
        RECT -111.835 93.245 -111.665 93.415 ;
        RECT -111.375 93.245 -111.205 93.415 ;
        RECT -104.215 93.245 -104.045 93.415 ;
        RECT -103.755 93.245 -103.585 93.415 ;
        RECT -103.295 93.245 -103.125 93.415 ;
        RECT -102.835 93.245 -102.665 93.415 ;
        RECT -102.375 93.245 -102.205 93.415 ;
        RECT -101.915 93.245 -101.745 93.415 ;
        RECT -101.455 93.245 -101.285 93.415 ;
        RECT -94.295 93.245 -94.125 93.415 ;
        RECT -93.835 93.245 -93.665 93.415 ;
        RECT -93.375 93.245 -93.205 93.415 ;
        RECT -92.915 93.245 -92.745 93.415 ;
        RECT -92.455 93.245 -92.285 93.415 ;
        RECT -91.995 93.245 -91.825 93.415 ;
        RECT -91.535 93.245 -91.365 93.415 ;
        RECT -84.375 93.245 -84.205 93.415 ;
        RECT -83.915 93.245 -83.745 93.415 ;
        RECT -83.455 93.245 -83.285 93.415 ;
        RECT -82.995 93.245 -82.825 93.415 ;
        RECT -82.535 93.245 -82.365 93.415 ;
        RECT -82.075 93.245 -81.905 93.415 ;
        RECT -81.615 93.245 -81.445 93.415 ;
        RECT -74.455 93.245 -74.285 93.415 ;
        RECT -73.995 93.245 -73.825 93.415 ;
        RECT -73.535 93.245 -73.365 93.415 ;
        RECT -73.075 93.245 -72.905 93.415 ;
        RECT -72.615 93.245 -72.445 93.415 ;
        RECT -72.155 93.245 -71.985 93.415 ;
        RECT -71.695 93.245 -71.525 93.415 ;
        RECT -64.535 93.245 -64.365 93.415 ;
        RECT -64.075 93.245 -63.905 93.415 ;
        RECT -63.615 93.245 -63.445 93.415 ;
        RECT -63.155 93.245 -62.985 93.415 ;
        RECT -62.695 93.245 -62.525 93.415 ;
        RECT -62.235 93.245 -62.065 93.415 ;
        RECT -61.775 93.245 -61.605 93.415 ;
        RECT -54.615 93.245 -54.445 93.415 ;
        RECT -54.155 93.245 -53.985 93.415 ;
        RECT -53.695 93.245 -53.525 93.415 ;
        RECT -53.235 93.245 -53.065 93.415 ;
        RECT -52.775 93.245 -52.605 93.415 ;
        RECT -52.315 93.245 -52.145 93.415 ;
        RECT -51.855 93.245 -51.685 93.415 ;
        RECT -44.695 93.245 -44.525 93.415 ;
        RECT -44.235 93.245 -44.065 93.415 ;
        RECT -43.775 93.245 -43.605 93.415 ;
        RECT -43.315 93.245 -43.145 93.415 ;
        RECT -42.855 93.245 -42.685 93.415 ;
        RECT -42.395 93.245 -42.225 93.415 ;
        RECT -41.935 93.245 -41.765 93.415 ;
        RECT -34.775 93.245 -34.605 93.415 ;
        RECT -34.315 93.245 -34.145 93.415 ;
        RECT -33.855 93.245 -33.685 93.415 ;
        RECT -33.395 93.245 -33.225 93.415 ;
        RECT -32.935 93.245 -32.765 93.415 ;
        RECT -32.475 93.245 -32.305 93.415 ;
        RECT -32.015 93.245 -31.845 93.415 ;
        RECT -24.855 93.245 -24.685 93.415 ;
        RECT -24.395 93.245 -24.225 93.415 ;
        RECT -23.935 93.245 -23.765 93.415 ;
        RECT -23.475 93.245 -23.305 93.415 ;
        RECT -23.015 93.245 -22.845 93.415 ;
        RECT -22.555 93.245 -22.385 93.415 ;
        RECT -22.095 93.245 -21.925 93.415 ;
        RECT -14.935 93.245 -14.765 93.415 ;
        RECT -14.475 93.245 -14.305 93.415 ;
        RECT -14.015 93.245 -13.845 93.415 ;
        RECT -13.555 93.245 -13.385 93.415 ;
        RECT -13.095 93.245 -12.925 93.415 ;
        RECT -12.635 93.245 -12.465 93.415 ;
        RECT -12.175 93.245 -12.005 93.415 ;
        RECT -5.015 93.245 -4.845 93.415 ;
        RECT -4.555 93.245 -4.385 93.415 ;
        RECT -4.095 93.245 -3.925 93.415 ;
        RECT -3.635 93.245 -3.465 93.415 ;
        RECT -3.175 93.245 -3.005 93.415 ;
        RECT -2.715 93.245 -2.545 93.415 ;
        RECT -2.255 93.245 -2.085 93.415 ;
        RECT 4.905 93.245 5.075 93.415 ;
        RECT 5.365 93.245 5.535 93.415 ;
        RECT 5.825 93.245 5.995 93.415 ;
        RECT 6.285 93.245 6.455 93.415 ;
        RECT 6.745 93.245 6.915 93.415 ;
        RECT 7.205 93.245 7.375 93.415 ;
        RECT 7.665 93.245 7.835 93.415 ;
        RECT 14.825 93.245 14.995 93.415 ;
        RECT 15.285 93.245 15.455 93.415 ;
        RECT 15.745 93.245 15.915 93.415 ;
        RECT 16.205 93.245 16.375 93.415 ;
        RECT 16.665 93.245 16.835 93.415 ;
        RECT 17.125 93.245 17.295 93.415 ;
        RECT 17.585 93.245 17.755 93.415 ;
        RECT -287.735 90.525 -287.565 90.695 ;
        RECT -287.275 90.525 -287.105 90.695 ;
        RECT -286.815 90.525 -286.645 90.695 ;
        RECT -286.355 90.525 -286.185 90.695 ;
        RECT -285.895 90.525 -285.725 90.695 ;
        RECT -285.435 90.525 -285.265 90.695 ;
        RECT -284.975 90.525 -284.805 90.695 ;
        RECT -277.815 90.525 -277.645 90.695 ;
        RECT -277.355 90.525 -277.185 90.695 ;
        RECT -276.895 90.525 -276.725 90.695 ;
        RECT -276.435 90.525 -276.265 90.695 ;
        RECT -275.975 90.525 -275.805 90.695 ;
        RECT -275.515 90.525 -275.345 90.695 ;
        RECT -275.055 90.525 -274.885 90.695 ;
        RECT -267.895 90.525 -267.725 90.695 ;
        RECT -267.435 90.525 -267.265 90.695 ;
        RECT -266.975 90.525 -266.805 90.695 ;
        RECT -266.515 90.525 -266.345 90.695 ;
        RECT -266.055 90.525 -265.885 90.695 ;
        RECT -265.595 90.525 -265.425 90.695 ;
        RECT -265.135 90.525 -264.965 90.695 ;
        RECT -257.975 90.525 -257.805 90.695 ;
        RECT -257.515 90.525 -257.345 90.695 ;
        RECT -257.055 90.525 -256.885 90.695 ;
        RECT -256.595 90.525 -256.425 90.695 ;
        RECT -256.135 90.525 -255.965 90.695 ;
        RECT -255.675 90.525 -255.505 90.695 ;
        RECT -255.215 90.525 -255.045 90.695 ;
        RECT -248.055 90.525 -247.885 90.695 ;
        RECT -247.595 90.525 -247.425 90.695 ;
        RECT -247.135 90.525 -246.965 90.695 ;
        RECT -246.675 90.525 -246.505 90.695 ;
        RECT -246.215 90.525 -246.045 90.695 ;
        RECT -245.755 90.525 -245.585 90.695 ;
        RECT -245.295 90.525 -245.125 90.695 ;
        RECT -238.135 90.525 -237.965 90.695 ;
        RECT -237.675 90.525 -237.505 90.695 ;
        RECT -237.215 90.525 -237.045 90.695 ;
        RECT -236.755 90.525 -236.585 90.695 ;
        RECT -236.295 90.525 -236.125 90.695 ;
        RECT -235.835 90.525 -235.665 90.695 ;
        RECT -235.375 90.525 -235.205 90.695 ;
        RECT -228.215 90.525 -228.045 90.695 ;
        RECT -227.755 90.525 -227.585 90.695 ;
        RECT -227.295 90.525 -227.125 90.695 ;
        RECT -226.835 90.525 -226.665 90.695 ;
        RECT -226.375 90.525 -226.205 90.695 ;
        RECT -225.915 90.525 -225.745 90.695 ;
        RECT -225.455 90.525 -225.285 90.695 ;
        RECT -218.295 90.525 -218.125 90.695 ;
        RECT -217.835 90.525 -217.665 90.695 ;
        RECT -217.375 90.525 -217.205 90.695 ;
        RECT -216.915 90.525 -216.745 90.695 ;
        RECT -216.455 90.525 -216.285 90.695 ;
        RECT -215.995 90.525 -215.825 90.695 ;
        RECT -215.535 90.525 -215.365 90.695 ;
        RECT -208.375 90.525 -208.205 90.695 ;
        RECT -207.915 90.525 -207.745 90.695 ;
        RECT -207.455 90.525 -207.285 90.695 ;
        RECT -206.995 90.525 -206.825 90.695 ;
        RECT -206.535 90.525 -206.365 90.695 ;
        RECT -206.075 90.525 -205.905 90.695 ;
        RECT -205.615 90.525 -205.445 90.695 ;
        RECT -198.455 90.525 -198.285 90.695 ;
        RECT -197.995 90.525 -197.825 90.695 ;
        RECT -197.535 90.525 -197.365 90.695 ;
        RECT -197.075 90.525 -196.905 90.695 ;
        RECT -196.615 90.525 -196.445 90.695 ;
        RECT -196.155 90.525 -195.985 90.695 ;
        RECT -195.695 90.525 -195.525 90.695 ;
        RECT -188.535 90.525 -188.365 90.695 ;
        RECT -188.075 90.525 -187.905 90.695 ;
        RECT -187.615 90.525 -187.445 90.695 ;
        RECT -187.155 90.525 -186.985 90.695 ;
        RECT -186.695 90.525 -186.525 90.695 ;
        RECT -186.235 90.525 -186.065 90.695 ;
        RECT -185.775 90.525 -185.605 90.695 ;
        RECT -178.615 90.525 -178.445 90.695 ;
        RECT -178.155 90.525 -177.985 90.695 ;
        RECT -177.695 90.525 -177.525 90.695 ;
        RECT -177.235 90.525 -177.065 90.695 ;
        RECT -176.775 90.525 -176.605 90.695 ;
        RECT -176.315 90.525 -176.145 90.695 ;
        RECT -175.855 90.525 -175.685 90.695 ;
        RECT -168.695 90.525 -168.525 90.695 ;
        RECT -168.235 90.525 -168.065 90.695 ;
        RECT -167.775 90.525 -167.605 90.695 ;
        RECT -167.315 90.525 -167.145 90.695 ;
        RECT -166.855 90.525 -166.685 90.695 ;
        RECT -166.395 90.525 -166.225 90.695 ;
        RECT -165.935 90.525 -165.765 90.695 ;
        RECT -158.775 90.525 -158.605 90.695 ;
        RECT -158.315 90.525 -158.145 90.695 ;
        RECT -157.855 90.525 -157.685 90.695 ;
        RECT -157.395 90.525 -157.225 90.695 ;
        RECT -156.935 90.525 -156.765 90.695 ;
        RECT -156.475 90.525 -156.305 90.695 ;
        RECT -156.015 90.525 -155.845 90.695 ;
        RECT -148.855 90.525 -148.685 90.695 ;
        RECT -148.395 90.525 -148.225 90.695 ;
        RECT -147.935 90.525 -147.765 90.695 ;
        RECT -147.475 90.525 -147.305 90.695 ;
        RECT -147.015 90.525 -146.845 90.695 ;
        RECT -146.555 90.525 -146.385 90.695 ;
        RECT -146.095 90.525 -145.925 90.695 ;
        RECT -138.935 90.525 -138.765 90.695 ;
        RECT -138.475 90.525 -138.305 90.695 ;
        RECT -138.015 90.525 -137.845 90.695 ;
        RECT -137.555 90.525 -137.385 90.695 ;
        RECT -137.095 90.525 -136.925 90.695 ;
        RECT -136.635 90.525 -136.465 90.695 ;
        RECT -136.175 90.525 -136.005 90.695 ;
        RECT -129.015 90.525 -128.845 90.695 ;
        RECT -128.555 90.525 -128.385 90.695 ;
        RECT -128.095 90.525 -127.925 90.695 ;
        RECT -127.635 90.525 -127.465 90.695 ;
        RECT -127.175 90.525 -127.005 90.695 ;
        RECT -126.715 90.525 -126.545 90.695 ;
        RECT -126.255 90.525 -126.085 90.695 ;
        RECT -119.095 90.525 -118.925 90.695 ;
        RECT -118.635 90.525 -118.465 90.695 ;
        RECT -118.175 90.525 -118.005 90.695 ;
        RECT -117.715 90.525 -117.545 90.695 ;
        RECT -117.255 90.525 -117.085 90.695 ;
        RECT -116.795 90.525 -116.625 90.695 ;
        RECT -116.335 90.525 -116.165 90.695 ;
        RECT -109.175 90.525 -109.005 90.695 ;
        RECT -108.715 90.525 -108.545 90.695 ;
        RECT -108.255 90.525 -108.085 90.695 ;
        RECT -107.795 90.525 -107.625 90.695 ;
        RECT -107.335 90.525 -107.165 90.695 ;
        RECT -106.875 90.525 -106.705 90.695 ;
        RECT -106.415 90.525 -106.245 90.695 ;
        RECT -99.255 90.525 -99.085 90.695 ;
        RECT -98.795 90.525 -98.625 90.695 ;
        RECT -98.335 90.525 -98.165 90.695 ;
        RECT -97.875 90.525 -97.705 90.695 ;
        RECT -97.415 90.525 -97.245 90.695 ;
        RECT -96.955 90.525 -96.785 90.695 ;
        RECT -96.495 90.525 -96.325 90.695 ;
        RECT -89.335 90.525 -89.165 90.695 ;
        RECT -88.875 90.525 -88.705 90.695 ;
        RECT -88.415 90.525 -88.245 90.695 ;
        RECT -87.955 90.525 -87.785 90.695 ;
        RECT -87.495 90.525 -87.325 90.695 ;
        RECT -87.035 90.525 -86.865 90.695 ;
        RECT -86.575 90.525 -86.405 90.695 ;
        RECT -79.415 90.525 -79.245 90.695 ;
        RECT -78.955 90.525 -78.785 90.695 ;
        RECT -78.495 90.525 -78.325 90.695 ;
        RECT -78.035 90.525 -77.865 90.695 ;
        RECT -77.575 90.525 -77.405 90.695 ;
        RECT -77.115 90.525 -76.945 90.695 ;
        RECT -76.655 90.525 -76.485 90.695 ;
        RECT -69.495 90.525 -69.325 90.695 ;
        RECT -69.035 90.525 -68.865 90.695 ;
        RECT -68.575 90.525 -68.405 90.695 ;
        RECT -68.115 90.525 -67.945 90.695 ;
        RECT -67.655 90.525 -67.485 90.695 ;
        RECT -67.195 90.525 -67.025 90.695 ;
        RECT -66.735 90.525 -66.565 90.695 ;
        RECT -59.575 90.525 -59.405 90.695 ;
        RECT -59.115 90.525 -58.945 90.695 ;
        RECT -58.655 90.525 -58.485 90.695 ;
        RECT -58.195 90.525 -58.025 90.695 ;
        RECT -57.735 90.525 -57.565 90.695 ;
        RECT -57.275 90.525 -57.105 90.695 ;
        RECT -56.815 90.525 -56.645 90.695 ;
        RECT -49.655 90.525 -49.485 90.695 ;
        RECT -49.195 90.525 -49.025 90.695 ;
        RECT -48.735 90.525 -48.565 90.695 ;
        RECT -48.275 90.525 -48.105 90.695 ;
        RECT -47.815 90.525 -47.645 90.695 ;
        RECT -47.355 90.525 -47.185 90.695 ;
        RECT -46.895 90.525 -46.725 90.695 ;
        RECT -39.735 90.525 -39.565 90.695 ;
        RECT -39.275 90.525 -39.105 90.695 ;
        RECT -38.815 90.525 -38.645 90.695 ;
        RECT -38.355 90.525 -38.185 90.695 ;
        RECT -37.895 90.525 -37.725 90.695 ;
        RECT -37.435 90.525 -37.265 90.695 ;
        RECT -36.975 90.525 -36.805 90.695 ;
        RECT -29.815 90.525 -29.645 90.695 ;
        RECT -29.355 90.525 -29.185 90.695 ;
        RECT -28.895 90.525 -28.725 90.695 ;
        RECT -28.435 90.525 -28.265 90.695 ;
        RECT -27.975 90.525 -27.805 90.695 ;
        RECT -27.515 90.525 -27.345 90.695 ;
        RECT -27.055 90.525 -26.885 90.695 ;
        RECT -19.895 90.525 -19.725 90.695 ;
        RECT -19.435 90.525 -19.265 90.695 ;
        RECT -18.975 90.525 -18.805 90.695 ;
        RECT -18.515 90.525 -18.345 90.695 ;
        RECT -18.055 90.525 -17.885 90.695 ;
        RECT -17.595 90.525 -17.425 90.695 ;
        RECT -17.135 90.525 -16.965 90.695 ;
        RECT -9.975 90.525 -9.805 90.695 ;
        RECT -9.515 90.525 -9.345 90.695 ;
        RECT -9.055 90.525 -8.885 90.695 ;
        RECT -8.595 90.525 -8.425 90.695 ;
        RECT -8.135 90.525 -7.965 90.695 ;
        RECT -7.675 90.525 -7.505 90.695 ;
        RECT -7.215 90.525 -7.045 90.695 ;
        RECT -0.055 90.525 0.115 90.695 ;
        RECT 0.405 90.525 0.575 90.695 ;
        RECT 0.865 90.525 1.035 90.695 ;
        RECT 1.325 90.525 1.495 90.695 ;
        RECT 1.785 90.525 1.955 90.695 ;
        RECT 2.245 90.525 2.415 90.695 ;
        RECT 2.705 90.525 2.875 90.695 ;
        RECT 9.865 90.525 10.035 90.695 ;
        RECT 10.325 90.525 10.495 90.695 ;
        RECT 10.785 90.525 10.955 90.695 ;
        RECT 11.245 90.525 11.415 90.695 ;
        RECT 11.705 90.525 11.875 90.695 ;
        RECT 12.165 90.525 12.335 90.695 ;
        RECT 12.625 90.525 12.795 90.695 ;
        RECT 19.785 90.525 19.955 90.695 ;
        RECT 20.245 90.525 20.415 90.695 ;
        RECT 20.705 90.525 20.875 90.695 ;
        RECT 21.165 90.525 21.335 90.695 ;
        RECT 21.625 90.525 21.795 90.695 ;
        RECT 22.085 90.525 22.255 90.695 ;
        RECT 22.545 90.525 22.715 90.695 ;
        RECT -283.165 89.865 -282.995 90.035 ;
        RECT -283.165 89.405 -282.995 89.575 ;
        RECT -279.625 89.865 -279.455 90.035 ;
        RECT -273.245 89.865 -273.075 90.035 ;
        RECT -279.625 89.405 -279.455 89.575 ;
        RECT -273.245 89.405 -273.075 89.575 ;
        RECT -281.395 89.135 -281.225 89.305 ;
        RECT -283.165 88.945 -282.995 89.115 ;
        RECT -279.625 88.945 -279.455 89.115 ;
        RECT -269.705 89.865 -269.535 90.035 ;
        RECT -263.325 89.865 -263.155 90.035 ;
        RECT -269.705 89.405 -269.535 89.575 ;
        RECT -263.325 89.405 -263.155 89.575 ;
        RECT -271.475 89.135 -271.305 89.305 ;
        RECT -273.245 88.945 -273.075 89.115 ;
        RECT -269.705 88.945 -269.535 89.115 ;
        RECT -259.785 89.865 -259.615 90.035 ;
        RECT -253.405 89.865 -253.235 90.035 ;
        RECT -259.785 89.405 -259.615 89.575 ;
        RECT -253.405 89.405 -253.235 89.575 ;
        RECT -261.555 89.135 -261.385 89.305 ;
        RECT -263.325 88.945 -263.155 89.115 ;
        RECT -259.785 88.945 -259.615 89.115 ;
        RECT -249.865 89.865 -249.695 90.035 ;
        RECT -243.485 89.865 -243.315 90.035 ;
        RECT -249.865 89.405 -249.695 89.575 ;
        RECT -243.485 89.405 -243.315 89.575 ;
        RECT -251.635 89.135 -251.465 89.305 ;
        RECT -253.405 88.945 -253.235 89.115 ;
        RECT -249.865 88.945 -249.695 89.115 ;
        RECT -239.945 89.865 -239.775 90.035 ;
        RECT -233.565 89.865 -233.395 90.035 ;
        RECT -239.945 89.405 -239.775 89.575 ;
        RECT -233.565 89.405 -233.395 89.575 ;
        RECT -241.715 89.135 -241.545 89.305 ;
        RECT -243.485 88.945 -243.315 89.115 ;
        RECT -239.945 88.945 -239.775 89.115 ;
        RECT -230.025 89.865 -229.855 90.035 ;
        RECT -223.645 89.865 -223.475 90.035 ;
        RECT -230.025 89.405 -229.855 89.575 ;
        RECT -223.645 89.405 -223.475 89.575 ;
        RECT -231.795 89.135 -231.625 89.305 ;
        RECT -233.565 88.945 -233.395 89.115 ;
        RECT -230.025 88.945 -229.855 89.115 ;
        RECT -220.105 89.865 -219.935 90.035 ;
        RECT -213.725 89.865 -213.555 90.035 ;
        RECT -220.105 89.405 -219.935 89.575 ;
        RECT -213.725 89.405 -213.555 89.575 ;
        RECT -221.875 89.135 -221.705 89.305 ;
        RECT -223.645 88.945 -223.475 89.115 ;
        RECT -220.105 88.945 -219.935 89.115 ;
        RECT -210.185 89.865 -210.015 90.035 ;
        RECT -203.805 89.865 -203.635 90.035 ;
        RECT -210.185 89.405 -210.015 89.575 ;
        RECT -203.805 89.405 -203.635 89.575 ;
        RECT -211.955 89.135 -211.785 89.305 ;
        RECT -213.725 88.945 -213.555 89.115 ;
        RECT -210.185 88.945 -210.015 89.115 ;
        RECT -200.265 89.865 -200.095 90.035 ;
        RECT -193.885 89.865 -193.715 90.035 ;
        RECT -200.265 89.405 -200.095 89.575 ;
        RECT -193.885 89.405 -193.715 89.575 ;
        RECT -202.035 89.135 -201.865 89.305 ;
        RECT -203.805 88.945 -203.635 89.115 ;
        RECT -200.265 88.945 -200.095 89.115 ;
        RECT -190.345 89.865 -190.175 90.035 ;
        RECT -183.965 89.865 -183.795 90.035 ;
        RECT -190.345 89.405 -190.175 89.575 ;
        RECT -183.965 89.405 -183.795 89.575 ;
        RECT -192.115 89.135 -191.945 89.305 ;
        RECT -193.885 88.945 -193.715 89.115 ;
        RECT -190.345 88.945 -190.175 89.115 ;
        RECT -180.425 89.865 -180.255 90.035 ;
        RECT -174.045 89.865 -173.875 90.035 ;
        RECT -180.425 89.405 -180.255 89.575 ;
        RECT -174.045 89.405 -173.875 89.575 ;
        RECT -182.195 89.135 -182.025 89.305 ;
        RECT -183.965 88.945 -183.795 89.115 ;
        RECT -180.425 88.945 -180.255 89.115 ;
        RECT -170.505 89.865 -170.335 90.035 ;
        RECT -164.125 89.865 -163.955 90.035 ;
        RECT -170.505 89.405 -170.335 89.575 ;
        RECT -164.125 89.405 -163.955 89.575 ;
        RECT -172.275 89.135 -172.105 89.305 ;
        RECT -174.045 88.945 -173.875 89.115 ;
        RECT -170.505 88.945 -170.335 89.115 ;
        RECT -160.585 89.865 -160.415 90.035 ;
        RECT -154.205 89.865 -154.035 90.035 ;
        RECT -160.585 89.405 -160.415 89.575 ;
        RECT -154.205 89.405 -154.035 89.575 ;
        RECT -162.355 89.135 -162.185 89.305 ;
        RECT -164.125 88.945 -163.955 89.115 ;
        RECT -160.585 88.945 -160.415 89.115 ;
        RECT -150.665 89.865 -150.495 90.035 ;
        RECT -144.285 89.865 -144.115 90.035 ;
        RECT -150.665 89.405 -150.495 89.575 ;
        RECT -144.285 89.405 -144.115 89.575 ;
        RECT -152.435 89.135 -152.265 89.305 ;
        RECT -154.205 88.945 -154.035 89.115 ;
        RECT -150.665 88.945 -150.495 89.115 ;
        RECT -140.745 89.865 -140.575 90.035 ;
        RECT -134.365 89.865 -134.195 90.035 ;
        RECT -140.745 89.405 -140.575 89.575 ;
        RECT -134.365 89.405 -134.195 89.575 ;
        RECT -142.515 89.135 -142.345 89.305 ;
        RECT -144.285 88.945 -144.115 89.115 ;
        RECT -140.745 88.945 -140.575 89.115 ;
        RECT -130.825 89.865 -130.655 90.035 ;
        RECT -124.445 89.865 -124.275 90.035 ;
        RECT -130.825 89.405 -130.655 89.575 ;
        RECT -124.445 89.405 -124.275 89.575 ;
        RECT -132.595 89.135 -132.425 89.305 ;
        RECT -134.365 88.945 -134.195 89.115 ;
        RECT -130.825 88.945 -130.655 89.115 ;
        RECT -120.905 89.865 -120.735 90.035 ;
        RECT -114.525 89.865 -114.355 90.035 ;
        RECT -120.905 89.405 -120.735 89.575 ;
        RECT -114.525 89.405 -114.355 89.575 ;
        RECT -122.675 89.135 -122.505 89.305 ;
        RECT -124.445 88.945 -124.275 89.115 ;
        RECT -120.905 88.945 -120.735 89.115 ;
        RECT -110.985 89.865 -110.815 90.035 ;
        RECT -104.605 89.865 -104.435 90.035 ;
        RECT -110.985 89.405 -110.815 89.575 ;
        RECT -104.605 89.405 -104.435 89.575 ;
        RECT -112.755 89.135 -112.585 89.305 ;
        RECT -114.525 88.945 -114.355 89.115 ;
        RECT -110.985 88.945 -110.815 89.115 ;
        RECT -101.065 89.865 -100.895 90.035 ;
        RECT -94.685 89.865 -94.515 90.035 ;
        RECT -101.065 89.405 -100.895 89.575 ;
        RECT -94.685 89.405 -94.515 89.575 ;
        RECT -102.835 89.135 -102.665 89.305 ;
        RECT -104.605 88.945 -104.435 89.115 ;
        RECT -101.065 88.945 -100.895 89.115 ;
        RECT -91.145 89.865 -90.975 90.035 ;
        RECT -84.765 89.865 -84.595 90.035 ;
        RECT -91.145 89.405 -90.975 89.575 ;
        RECT -84.765 89.405 -84.595 89.575 ;
        RECT -92.915 89.135 -92.745 89.305 ;
        RECT -94.685 88.945 -94.515 89.115 ;
        RECT -91.145 88.945 -90.975 89.115 ;
        RECT -81.225 89.865 -81.055 90.035 ;
        RECT -74.845 89.865 -74.675 90.035 ;
        RECT -81.225 89.405 -81.055 89.575 ;
        RECT -74.845 89.405 -74.675 89.575 ;
        RECT -82.995 89.135 -82.825 89.305 ;
        RECT -84.765 88.945 -84.595 89.115 ;
        RECT -81.225 88.945 -81.055 89.115 ;
        RECT -71.305 89.865 -71.135 90.035 ;
        RECT -64.925 89.865 -64.755 90.035 ;
        RECT -71.305 89.405 -71.135 89.575 ;
        RECT -64.925 89.405 -64.755 89.575 ;
        RECT -73.075 89.135 -72.905 89.305 ;
        RECT -74.845 88.945 -74.675 89.115 ;
        RECT -71.305 88.945 -71.135 89.115 ;
        RECT -61.385 89.865 -61.215 90.035 ;
        RECT -55.005 89.865 -54.835 90.035 ;
        RECT -61.385 89.405 -61.215 89.575 ;
        RECT -55.005 89.405 -54.835 89.575 ;
        RECT -63.155 89.135 -62.985 89.305 ;
        RECT -64.925 88.945 -64.755 89.115 ;
        RECT -61.385 88.945 -61.215 89.115 ;
        RECT -51.465 89.865 -51.295 90.035 ;
        RECT -45.085 89.865 -44.915 90.035 ;
        RECT -51.465 89.405 -51.295 89.575 ;
        RECT -45.085 89.405 -44.915 89.575 ;
        RECT -53.235 89.135 -53.065 89.305 ;
        RECT -55.005 88.945 -54.835 89.115 ;
        RECT -51.465 88.945 -51.295 89.115 ;
        RECT -41.545 89.865 -41.375 90.035 ;
        RECT -35.165 89.865 -34.995 90.035 ;
        RECT -41.545 89.405 -41.375 89.575 ;
        RECT -35.165 89.405 -34.995 89.575 ;
        RECT -43.315 89.135 -43.145 89.305 ;
        RECT -45.085 88.945 -44.915 89.115 ;
        RECT -41.545 88.945 -41.375 89.115 ;
        RECT -31.625 89.865 -31.455 90.035 ;
        RECT -25.245 89.865 -25.075 90.035 ;
        RECT -31.625 89.405 -31.455 89.575 ;
        RECT -25.245 89.405 -25.075 89.575 ;
        RECT -33.395 89.135 -33.225 89.305 ;
        RECT -35.165 88.945 -34.995 89.115 ;
        RECT -31.625 88.945 -31.455 89.115 ;
        RECT -21.705 89.865 -21.535 90.035 ;
        RECT -15.325 89.865 -15.155 90.035 ;
        RECT -21.705 89.405 -21.535 89.575 ;
        RECT -15.325 89.405 -15.155 89.575 ;
        RECT -23.475 89.135 -23.305 89.305 ;
        RECT -25.245 88.945 -25.075 89.115 ;
        RECT -21.705 88.945 -21.535 89.115 ;
        RECT -11.785 89.865 -11.615 90.035 ;
        RECT -5.405 89.865 -5.235 90.035 ;
        RECT -11.785 89.405 -11.615 89.575 ;
        RECT -5.405 89.405 -5.235 89.575 ;
        RECT -13.555 89.135 -13.385 89.305 ;
        RECT -15.325 88.945 -15.155 89.115 ;
        RECT -11.785 88.945 -11.615 89.115 ;
        RECT -1.865 89.865 -1.695 90.035 ;
        RECT 4.515 89.865 4.685 90.035 ;
        RECT -1.865 89.405 -1.695 89.575 ;
        RECT 4.515 89.405 4.685 89.575 ;
        RECT -3.635 89.135 -3.465 89.305 ;
        RECT -5.405 88.945 -5.235 89.115 ;
        RECT -1.865 88.945 -1.695 89.115 ;
        RECT 8.055 89.865 8.225 90.035 ;
        RECT 14.435 89.865 14.605 90.035 ;
        RECT 8.055 89.405 8.225 89.575 ;
        RECT 14.435 89.405 14.605 89.575 ;
        RECT 6.285 89.135 6.455 89.305 ;
        RECT 4.515 88.945 4.685 89.115 ;
        RECT 8.055 88.945 8.225 89.115 ;
        RECT 17.975 89.865 18.145 90.035 ;
        RECT 17.975 89.405 18.145 89.575 ;
        RECT 16.205 89.135 16.375 89.305 ;
        RECT 14.435 88.945 14.605 89.115 ;
        RECT 17.975 88.945 18.145 89.115 ;
        RECT -290.145 10.775 -289.975 10.945 ;
        RECT -288.375 10.675 -288.205 10.845 ;
        RECT -286.605 10.775 -286.435 10.945 ;
        RECT -290.145 10.315 -289.975 10.485 ;
        RECT -290.145 9.855 -289.975 10.025 ;
        RECT -280.225 10.775 -280.055 10.945 ;
        RECT -278.455 10.675 -278.285 10.845 ;
        RECT -276.685 10.775 -276.515 10.945 ;
        RECT -286.605 10.315 -286.435 10.485 ;
        RECT -280.225 10.315 -280.055 10.485 ;
        RECT -286.605 9.855 -286.435 10.025 ;
        RECT -280.225 9.855 -280.055 10.025 ;
        RECT -270.305 10.775 -270.135 10.945 ;
        RECT -268.535 10.675 -268.365 10.845 ;
        RECT -266.765 10.775 -266.595 10.945 ;
        RECT -276.685 10.315 -276.515 10.485 ;
        RECT -270.305 10.315 -270.135 10.485 ;
        RECT -276.685 9.855 -276.515 10.025 ;
        RECT -270.305 9.855 -270.135 10.025 ;
        RECT -260.385 10.775 -260.215 10.945 ;
        RECT -258.615 10.675 -258.445 10.845 ;
        RECT -256.845 10.775 -256.675 10.945 ;
        RECT -266.765 10.315 -266.595 10.485 ;
        RECT -260.385 10.315 -260.215 10.485 ;
        RECT -266.765 9.855 -266.595 10.025 ;
        RECT -260.385 9.855 -260.215 10.025 ;
        RECT -250.465 10.775 -250.295 10.945 ;
        RECT -248.695 10.675 -248.525 10.845 ;
        RECT -246.925 10.775 -246.755 10.945 ;
        RECT -256.845 10.315 -256.675 10.485 ;
        RECT -250.465 10.315 -250.295 10.485 ;
        RECT -256.845 9.855 -256.675 10.025 ;
        RECT -250.465 9.855 -250.295 10.025 ;
        RECT -240.545 10.775 -240.375 10.945 ;
        RECT -238.775 10.675 -238.605 10.845 ;
        RECT -237.005 10.775 -236.835 10.945 ;
        RECT -246.925 10.315 -246.755 10.485 ;
        RECT -240.545 10.315 -240.375 10.485 ;
        RECT -246.925 9.855 -246.755 10.025 ;
        RECT -240.545 9.855 -240.375 10.025 ;
        RECT -230.625 10.775 -230.455 10.945 ;
        RECT -228.855 10.675 -228.685 10.845 ;
        RECT -227.085 10.775 -226.915 10.945 ;
        RECT -237.005 10.315 -236.835 10.485 ;
        RECT -230.625 10.315 -230.455 10.485 ;
        RECT -237.005 9.855 -236.835 10.025 ;
        RECT -230.625 9.855 -230.455 10.025 ;
        RECT -220.705 10.775 -220.535 10.945 ;
        RECT -218.935 10.675 -218.765 10.845 ;
        RECT -217.165 10.775 -216.995 10.945 ;
        RECT -227.085 10.315 -226.915 10.485 ;
        RECT -220.705 10.315 -220.535 10.485 ;
        RECT -227.085 9.855 -226.915 10.025 ;
        RECT -220.705 9.855 -220.535 10.025 ;
        RECT -210.785 10.775 -210.615 10.945 ;
        RECT -209.015 10.675 -208.845 10.845 ;
        RECT -207.245 10.775 -207.075 10.945 ;
        RECT -217.165 10.315 -216.995 10.485 ;
        RECT -210.785 10.315 -210.615 10.485 ;
        RECT -217.165 9.855 -216.995 10.025 ;
        RECT -210.785 9.855 -210.615 10.025 ;
        RECT -200.865 10.775 -200.695 10.945 ;
        RECT -199.095 10.675 -198.925 10.845 ;
        RECT -197.325 10.775 -197.155 10.945 ;
        RECT -207.245 10.315 -207.075 10.485 ;
        RECT -200.865 10.315 -200.695 10.485 ;
        RECT -207.245 9.855 -207.075 10.025 ;
        RECT -200.865 9.855 -200.695 10.025 ;
        RECT -190.945 10.775 -190.775 10.945 ;
        RECT -189.175 10.675 -189.005 10.845 ;
        RECT -187.405 10.775 -187.235 10.945 ;
        RECT -197.325 10.315 -197.155 10.485 ;
        RECT -190.945 10.315 -190.775 10.485 ;
        RECT -197.325 9.855 -197.155 10.025 ;
        RECT -190.945 9.855 -190.775 10.025 ;
        RECT -181.025 10.775 -180.855 10.945 ;
        RECT -179.255 10.675 -179.085 10.845 ;
        RECT -177.485 10.775 -177.315 10.945 ;
        RECT -187.405 10.315 -187.235 10.485 ;
        RECT -181.025 10.315 -180.855 10.485 ;
        RECT -187.405 9.855 -187.235 10.025 ;
        RECT -181.025 9.855 -180.855 10.025 ;
        RECT -171.105 10.775 -170.935 10.945 ;
        RECT -169.335 10.675 -169.165 10.845 ;
        RECT -167.565 10.775 -167.395 10.945 ;
        RECT -177.485 10.315 -177.315 10.485 ;
        RECT -171.105 10.315 -170.935 10.485 ;
        RECT -177.485 9.855 -177.315 10.025 ;
        RECT -171.105 9.855 -170.935 10.025 ;
        RECT -161.185 10.775 -161.015 10.945 ;
        RECT -159.415 10.675 -159.245 10.845 ;
        RECT -157.645 10.775 -157.475 10.945 ;
        RECT -167.565 10.315 -167.395 10.485 ;
        RECT -161.185 10.315 -161.015 10.485 ;
        RECT -167.565 9.855 -167.395 10.025 ;
        RECT -161.185 9.855 -161.015 10.025 ;
        RECT -151.265 10.775 -151.095 10.945 ;
        RECT -149.495 10.675 -149.325 10.845 ;
        RECT -147.725 10.775 -147.555 10.945 ;
        RECT -157.645 10.315 -157.475 10.485 ;
        RECT -151.265 10.315 -151.095 10.485 ;
        RECT -157.645 9.855 -157.475 10.025 ;
        RECT -151.265 9.855 -151.095 10.025 ;
        RECT -141.345 10.775 -141.175 10.945 ;
        RECT -139.575 10.675 -139.405 10.845 ;
        RECT -137.805 10.775 -137.635 10.945 ;
        RECT -147.725 10.315 -147.555 10.485 ;
        RECT -141.345 10.315 -141.175 10.485 ;
        RECT -147.725 9.855 -147.555 10.025 ;
        RECT -141.345 9.855 -141.175 10.025 ;
        RECT -131.425 10.775 -131.255 10.945 ;
        RECT -129.655 10.675 -129.485 10.845 ;
        RECT -127.885 10.775 -127.715 10.945 ;
        RECT -137.805 10.315 -137.635 10.485 ;
        RECT -131.425 10.315 -131.255 10.485 ;
        RECT -137.805 9.855 -137.635 10.025 ;
        RECT -131.425 9.855 -131.255 10.025 ;
        RECT -121.505 10.775 -121.335 10.945 ;
        RECT -119.735 10.675 -119.565 10.845 ;
        RECT -117.965 10.775 -117.795 10.945 ;
        RECT -127.885 10.315 -127.715 10.485 ;
        RECT -121.505 10.315 -121.335 10.485 ;
        RECT -127.885 9.855 -127.715 10.025 ;
        RECT -121.505 9.855 -121.335 10.025 ;
        RECT -111.585 10.775 -111.415 10.945 ;
        RECT -109.815 10.675 -109.645 10.845 ;
        RECT -108.045 10.775 -107.875 10.945 ;
        RECT -117.965 10.315 -117.795 10.485 ;
        RECT -111.585 10.315 -111.415 10.485 ;
        RECT -117.965 9.855 -117.795 10.025 ;
        RECT -111.585 9.855 -111.415 10.025 ;
        RECT -101.665 10.775 -101.495 10.945 ;
        RECT -99.895 10.675 -99.725 10.845 ;
        RECT -98.125 10.775 -97.955 10.945 ;
        RECT -108.045 10.315 -107.875 10.485 ;
        RECT -101.665 10.315 -101.495 10.485 ;
        RECT -108.045 9.855 -107.875 10.025 ;
        RECT -101.665 9.855 -101.495 10.025 ;
        RECT -91.745 10.775 -91.575 10.945 ;
        RECT -89.975 10.675 -89.805 10.845 ;
        RECT -88.205 10.775 -88.035 10.945 ;
        RECT -98.125 10.315 -97.955 10.485 ;
        RECT -91.745 10.315 -91.575 10.485 ;
        RECT -98.125 9.855 -97.955 10.025 ;
        RECT -91.745 9.855 -91.575 10.025 ;
        RECT -81.825 10.775 -81.655 10.945 ;
        RECT -80.055 10.675 -79.885 10.845 ;
        RECT -78.285 10.775 -78.115 10.945 ;
        RECT -88.205 10.315 -88.035 10.485 ;
        RECT -81.825 10.315 -81.655 10.485 ;
        RECT -88.205 9.855 -88.035 10.025 ;
        RECT -81.825 9.855 -81.655 10.025 ;
        RECT -71.905 10.775 -71.735 10.945 ;
        RECT -70.135 10.675 -69.965 10.845 ;
        RECT -68.365 10.775 -68.195 10.945 ;
        RECT -78.285 10.315 -78.115 10.485 ;
        RECT -71.905 10.315 -71.735 10.485 ;
        RECT -78.285 9.855 -78.115 10.025 ;
        RECT -71.905 9.855 -71.735 10.025 ;
        RECT -61.985 10.775 -61.815 10.945 ;
        RECT -60.215 10.675 -60.045 10.845 ;
        RECT -58.445 10.775 -58.275 10.945 ;
        RECT -68.365 10.315 -68.195 10.485 ;
        RECT -61.985 10.315 -61.815 10.485 ;
        RECT -68.365 9.855 -68.195 10.025 ;
        RECT -61.985 9.855 -61.815 10.025 ;
        RECT -52.065 10.775 -51.895 10.945 ;
        RECT -50.295 10.675 -50.125 10.845 ;
        RECT -48.525 10.775 -48.355 10.945 ;
        RECT -58.445 10.315 -58.275 10.485 ;
        RECT -52.065 10.315 -51.895 10.485 ;
        RECT -58.445 9.855 -58.275 10.025 ;
        RECT -52.065 9.855 -51.895 10.025 ;
        RECT -42.145 10.775 -41.975 10.945 ;
        RECT -40.375 10.675 -40.205 10.845 ;
        RECT -38.605 10.775 -38.435 10.945 ;
        RECT -48.525 10.315 -48.355 10.485 ;
        RECT -42.145 10.315 -41.975 10.485 ;
        RECT -48.525 9.855 -48.355 10.025 ;
        RECT -42.145 9.855 -41.975 10.025 ;
        RECT -32.225 10.775 -32.055 10.945 ;
        RECT -30.455 10.675 -30.285 10.845 ;
        RECT -28.685 10.775 -28.515 10.945 ;
        RECT -38.605 10.315 -38.435 10.485 ;
        RECT -32.225 10.315 -32.055 10.485 ;
        RECT -38.605 9.855 -38.435 10.025 ;
        RECT -32.225 9.855 -32.055 10.025 ;
        RECT -22.305 10.775 -22.135 10.945 ;
        RECT -20.535 10.675 -20.365 10.845 ;
        RECT -18.765 10.775 -18.595 10.945 ;
        RECT -28.685 10.315 -28.515 10.485 ;
        RECT -22.305 10.315 -22.135 10.485 ;
        RECT -28.685 9.855 -28.515 10.025 ;
        RECT -22.305 9.855 -22.135 10.025 ;
        RECT -12.385 10.775 -12.215 10.945 ;
        RECT -10.615 10.675 -10.445 10.845 ;
        RECT -8.845 10.775 -8.675 10.945 ;
        RECT -18.765 10.315 -18.595 10.485 ;
        RECT -12.385 10.315 -12.215 10.485 ;
        RECT -18.765 9.855 -18.595 10.025 ;
        RECT -12.385 9.855 -12.215 10.025 ;
        RECT -2.465 10.775 -2.295 10.945 ;
        RECT -0.695 10.675 -0.525 10.845 ;
        RECT 1.075 10.775 1.245 10.945 ;
        RECT -8.845 10.315 -8.675 10.485 ;
        RECT -2.465 10.315 -2.295 10.485 ;
        RECT -8.845 9.855 -8.675 10.025 ;
        RECT -2.465 9.855 -2.295 10.025 ;
        RECT 7.455 10.775 7.625 10.945 ;
        RECT 9.225 10.675 9.395 10.845 ;
        RECT 10.995 10.775 11.165 10.945 ;
        RECT 1.075 10.315 1.245 10.485 ;
        RECT 7.455 10.315 7.625 10.485 ;
        RECT 1.075 9.855 1.245 10.025 ;
        RECT 7.455 9.855 7.625 10.025 ;
        RECT 17.375 10.775 17.545 10.945 ;
        RECT 19.145 10.675 19.315 10.845 ;
        RECT 20.915 10.775 21.085 10.945 ;
        RECT 10.995 10.315 11.165 10.485 ;
        RECT 17.375 10.315 17.545 10.485 ;
        RECT 10.995 9.855 11.165 10.025 ;
        RECT 17.375 9.855 17.545 10.025 ;
        RECT 20.915 10.315 21.085 10.485 ;
        RECT 20.915 9.855 21.085 10.025 ;
        RECT -284.795 9.195 -284.625 9.365 ;
        RECT -284.335 9.195 -284.165 9.365 ;
        RECT -283.875 9.195 -283.705 9.365 ;
        RECT -283.415 9.195 -283.245 9.365 ;
        RECT -282.955 9.195 -282.785 9.365 ;
        RECT -282.495 9.195 -282.325 9.365 ;
        RECT -282.035 9.195 -281.865 9.365 ;
        RECT -274.875 9.195 -274.705 9.365 ;
        RECT -274.415 9.195 -274.245 9.365 ;
        RECT -273.955 9.195 -273.785 9.365 ;
        RECT -273.495 9.195 -273.325 9.365 ;
        RECT -273.035 9.195 -272.865 9.365 ;
        RECT -272.575 9.195 -272.405 9.365 ;
        RECT -272.115 9.195 -271.945 9.365 ;
        RECT -264.955 9.195 -264.785 9.365 ;
        RECT -264.495 9.195 -264.325 9.365 ;
        RECT -264.035 9.195 -263.865 9.365 ;
        RECT -263.575 9.195 -263.405 9.365 ;
        RECT -263.115 9.195 -262.945 9.365 ;
        RECT -262.655 9.195 -262.485 9.365 ;
        RECT -262.195 9.195 -262.025 9.365 ;
        RECT -255.035 9.195 -254.865 9.365 ;
        RECT -254.575 9.195 -254.405 9.365 ;
        RECT -254.115 9.195 -253.945 9.365 ;
        RECT -253.655 9.195 -253.485 9.365 ;
        RECT -253.195 9.195 -253.025 9.365 ;
        RECT -252.735 9.195 -252.565 9.365 ;
        RECT -252.275 9.195 -252.105 9.365 ;
        RECT -245.115 9.195 -244.945 9.365 ;
        RECT -244.655 9.195 -244.485 9.365 ;
        RECT -244.195 9.195 -244.025 9.365 ;
        RECT -243.735 9.195 -243.565 9.365 ;
        RECT -243.275 9.195 -243.105 9.365 ;
        RECT -242.815 9.195 -242.645 9.365 ;
        RECT -242.355 9.195 -242.185 9.365 ;
        RECT -235.195 9.195 -235.025 9.365 ;
        RECT -234.735 9.195 -234.565 9.365 ;
        RECT -234.275 9.195 -234.105 9.365 ;
        RECT -233.815 9.195 -233.645 9.365 ;
        RECT -233.355 9.195 -233.185 9.365 ;
        RECT -232.895 9.195 -232.725 9.365 ;
        RECT -232.435 9.195 -232.265 9.365 ;
        RECT -225.275 9.195 -225.105 9.365 ;
        RECT -224.815 9.195 -224.645 9.365 ;
        RECT -224.355 9.195 -224.185 9.365 ;
        RECT -223.895 9.195 -223.725 9.365 ;
        RECT -223.435 9.195 -223.265 9.365 ;
        RECT -222.975 9.195 -222.805 9.365 ;
        RECT -222.515 9.195 -222.345 9.365 ;
        RECT -215.355 9.195 -215.185 9.365 ;
        RECT -214.895 9.195 -214.725 9.365 ;
        RECT -214.435 9.195 -214.265 9.365 ;
        RECT -213.975 9.195 -213.805 9.365 ;
        RECT -213.515 9.195 -213.345 9.365 ;
        RECT -213.055 9.195 -212.885 9.365 ;
        RECT -212.595 9.195 -212.425 9.365 ;
        RECT -205.435 9.195 -205.265 9.365 ;
        RECT -204.975 9.195 -204.805 9.365 ;
        RECT -204.515 9.195 -204.345 9.365 ;
        RECT -204.055 9.195 -203.885 9.365 ;
        RECT -203.595 9.195 -203.425 9.365 ;
        RECT -203.135 9.195 -202.965 9.365 ;
        RECT -202.675 9.195 -202.505 9.365 ;
        RECT -195.515 9.195 -195.345 9.365 ;
        RECT -195.055 9.195 -194.885 9.365 ;
        RECT -194.595 9.195 -194.425 9.365 ;
        RECT -194.135 9.195 -193.965 9.365 ;
        RECT -193.675 9.195 -193.505 9.365 ;
        RECT -193.215 9.195 -193.045 9.365 ;
        RECT -192.755 9.195 -192.585 9.365 ;
        RECT -185.595 9.195 -185.425 9.365 ;
        RECT -185.135 9.195 -184.965 9.365 ;
        RECT -184.675 9.195 -184.505 9.365 ;
        RECT -184.215 9.195 -184.045 9.365 ;
        RECT -183.755 9.195 -183.585 9.365 ;
        RECT -183.295 9.195 -183.125 9.365 ;
        RECT -182.835 9.195 -182.665 9.365 ;
        RECT -175.675 9.195 -175.505 9.365 ;
        RECT -175.215 9.195 -175.045 9.365 ;
        RECT -174.755 9.195 -174.585 9.365 ;
        RECT -174.295 9.195 -174.125 9.365 ;
        RECT -173.835 9.195 -173.665 9.365 ;
        RECT -173.375 9.195 -173.205 9.365 ;
        RECT -172.915 9.195 -172.745 9.365 ;
        RECT -165.755 9.195 -165.585 9.365 ;
        RECT -165.295 9.195 -165.125 9.365 ;
        RECT -164.835 9.195 -164.665 9.365 ;
        RECT -164.375 9.195 -164.205 9.365 ;
        RECT -163.915 9.195 -163.745 9.365 ;
        RECT -163.455 9.195 -163.285 9.365 ;
        RECT -162.995 9.195 -162.825 9.365 ;
        RECT -155.835 9.195 -155.665 9.365 ;
        RECT -155.375 9.195 -155.205 9.365 ;
        RECT -154.915 9.195 -154.745 9.365 ;
        RECT -154.455 9.195 -154.285 9.365 ;
        RECT -153.995 9.195 -153.825 9.365 ;
        RECT -153.535 9.195 -153.365 9.365 ;
        RECT -153.075 9.195 -152.905 9.365 ;
        RECT -145.915 9.195 -145.745 9.365 ;
        RECT -145.455 9.195 -145.285 9.365 ;
        RECT -144.995 9.195 -144.825 9.365 ;
        RECT -144.535 9.195 -144.365 9.365 ;
        RECT -144.075 9.195 -143.905 9.365 ;
        RECT -143.615 9.195 -143.445 9.365 ;
        RECT -143.155 9.195 -142.985 9.365 ;
        RECT -135.995 9.195 -135.825 9.365 ;
        RECT -135.535 9.195 -135.365 9.365 ;
        RECT -135.075 9.195 -134.905 9.365 ;
        RECT -134.615 9.195 -134.445 9.365 ;
        RECT -134.155 9.195 -133.985 9.365 ;
        RECT -133.695 9.195 -133.525 9.365 ;
        RECT -133.235 9.195 -133.065 9.365 ;
        RECT -126.075 9.195 -125.905 9.365 ;
        RECT -125.615 9.195 -125.445 9.365 ;
        RECT -125.155 9.195 -124.985 9.365 ;
        RECT -124.695 9.195 -124.525 9.365 ;
        RECT -124.235 9.195 -124.065 9.365 ;
        RECT -123.775 9.195 -123.605 9.365 ;
        RECT -123.315 9.195 -123.145 9.365 ;
        RECT -116.155 9.195 -115.985 9.365 ;
        RECT -115.695 9.195 -115.525 9.365 ;
        RECT -115.235 9.195 -115.065 9.365 ;
        RECT -114.775 9.195 -114.605 9.365 ;
        RECT -114.315 9.195 -114.145 9.365 ;
        RECT -113.855 9.195 -113.685 9.365 ;
        RECT -113.395 9.195 -113.225 9.365 ;
        RECT -106.235 9.195 -106.065 9.365 ;
        RECT -105.775 9.195 -105.605 9.365 ;
        RECT -105.315 9.195 -105.145 9.365 ;
        RECT -104.855 9.195 -104.685 9.365 ;
        RECT -104.395 9.195 -104.225 9.365 ;
        RECT -103.935 9.195 -103.765 9.365 ;
        RECT -103.475 9.195 -103.305 9.365 ;
        RECT -96.315 9.195 -96.145 9.365 ;
        RECT -95.855 9.195 -95.685 9.365 ;
        RECT -95.395 9.195 -95.225 9.365 ;
        RECT -94.935 9.195 -94.765 9.365 ;
        RECT -94.475 9.195 -94.305 9.365 ;
        RECT -94.015 9.195 -93.845 9.365 ;
        RECT -93.555 9.195 -93.385 9.365 ;
        RECT -86.395 9.195 -86.225 9.365 ;
        RECT -85.935 9.195 -85.765 9.365 ;
        RECT -85.475 9.195 -85.305 9.365 ;
        RECT -85.015 9.195 -84.845 9.365 ;
        RECT -84.555 9.195 -84.385 9.365 ;
        RECT -84.095 9.195 -83.925 9.365 ;
        RECT -83.635 9.195 -83.465 9.365 ;
        RECT -76.475 9.195 -76.305 9.365 ;
        RECT -76.015 9.195 -75.845 9.365 ;
        RECT -75.555 9.195 -75.385 9.365 ;
        RECT -75.095 9.195 -74.925 9.365 ;
        RECT -74.635 9.195 -74.465 9.365 ;
        RECT -74.175 9.195 -74.005 9.365 ;
        RECT -73.715 9.195 -73.545 9.365 ;
        RECT -66.555 9.195 -66.385 9.365 ;
        RECT -66.095 9.195 -65.925 9.365 ;
        RECT -65.635 9.195 -65.465 9.365 ;
        RECT -65.175 9.195 -65.005 9.365 ;
        RECT -64.715 9.195 -64.545 9.365 ;
        RECT -64.255 9.195 -64.085 9.365 ;
        RECT -63.795 9.195 -63.625 9.365 ;
        RECT -56.635 9.195 -56.465 9.365 ;
        RECT -56.175 9.195 -56.005 9.365 ;
        RECT -55.715 9.195 -55.545 9.365 ;
        RECT -55.255 9.195 -55.085 9.365 ;
        RECT -54.795 9.195 -54.625 9.365 ;
        RECT -54.335 9.195 -54.165 9.365 ;
        RECT -53.875 9.195 -53.705 9.365 ;
        RECT -46.715 9.195 -46.545 9.365 ;
        RECT -46.255 9.195 -46.085 9.365 ;
        RECT -45.795 9.195 -45.625 9.365 ;
        RECT -45.335 9.195 -45.165 9.365 ;
        RECT -44.875 9.195 -44.705 9.365 ;
        RECT -44.415 9.195 -44.245 9.365 ;
        RECT -43.955 9.195 -43.785 9.365 ;
        RECT -36.795 9.195 -36.625 9.365 ;
        RECT -36.335 9.195 -36.165 9.365 ;
        RECT -35.875 9.195 -35.705 9.365 ;
        RECT -35.415 9.195 -35.245 9.365 ;
        RECT -34.955 9.195 -34.785 9.365 ;
        RECT -34.495 9.195 -34.325 9.365 ;
        RECT -34.035 9.195 -33.865 9.365 ;
        RECT -26.875 9.195 -26.705 9.365 ;
        RECT -26.415 9.195 -26.245 9.365 ;
        RECT -25.955 9.195 -25.785 9.365 ;
        RECT -25.495 9.195 -25.325 9.365 ;
        RECT -25.035 9.195 -24.865 9.365 ;
        RECT -24.575 9.195 -24.405 9.365 ;
        RECT -24.115 9.195 -23.945 9.365 ;
        RECT -16.955 9.195 -16.785 9.365 ;
        RECT -16.495 9.195 -16.325 9.365 ;
        RECT -16.035 9.195 -15.865 9.365 ;
        RECT -15.575 9.195 -15.405 9.365 ;
        RECT -15.115 9.195 -14.945 9.365 ;
        RECT -14.655 9.195 -14.485 9.365 ;
        RECT -14.195 9.195 -14.025 9.365 ;
        RECT -7.035 9.195 -6.865 9.365 ;
        RECT -6.575 9.195 -6.405 9.365 ;
        RECT -6.115 9.195 -5.945 9.365 ;
        RECT -5.655 9.195 -5.485 9.365 ;
        RECT -5.195 9.195 -5.025 9.365 ;
        RECT -4.735 9.195 -4.565 9.365 ;
        RECT -4.275 9.195 -4.105 9.365 ;
        RECT 2.885 9.195 3.055 9.365 ;
        RECT 3.345 9.195 3.515 9.365 ;
        RECT 3.805 9.195 3.975 9.365 ;
        RECT 4.265 9.195 4.435 9.365 ;
        RECT 4.725 9.195 4.895 9.365 ;
        RECT 5.185 9.195 5.355 9.365 ;
        RECT 5.645 9.195 5.815 9.365 ;
        RECT 12.805 9.195 12.975 9.365 ;
        RECT 13.265 9.195 13.435 9.365 ;
        RECT 13.725 9.195 13.895 9.365 ;
        RECT 14.185 9.195 14.355 9.365 ;
        RECT 14.645 9.195 14.815 9.365 ;
        RECT 15.105 9.195 15.275 9.365 ;
        RECT 15.565 9.195 15.735 9.365 ;
        RECT -289.755 6.475 -289.585 6.645 ;
        RECT -289.295 6.475 -289.125 6.645 ;
        RECT -288.835 6.475 -288.665 6.645 ;
        RECT -288.375 6.475 -288.205 6.645 ;
        RECT -287.915 6.475 -287.745 6.645 ;
        RECT -287.455 6.475 -287.285 6.645 ;
        RECT -286.995 6.475 -286.825 6.645 ;
        RECT -279.835 6.475 -279.665 6.645 ;
        RECT -279.375 6.475 -279.205 6.645 ;
        RECT -278.915 6.475 -278.745 6.645 ;
        RECT -278.455 6.475 -278.285 6.645 ;
        RECT -277.995 6.475 -277.825 6.645 ;
        RECT -277.535 6.475 -277.365 6.645 ;
        RECT -277.075 6.475 -276.905 6.645 ;
        RECT -269.915 6.475 -269.745 6.645 ;
        RECT -269.455 6.475 -269.285 6.645 ;
        RECT -268.995 6.475 -268.825 6.645 ;
        RECT -268.535 6.475 -268.365 6.645 ;
        RECT -268.075 6.475 -267.905 6.645 ;
        RECT -267.615 6.475 -267.445 6.645 ;
        RECT -267.155 6.475 -266.985 6.645 ;
        RECT -259.995 6.475 -259.825 6.645 ;
        RECT -259.535 6.475 -259.365 6.645 ;
        RECT -259.075 6.475 -258.905 6.645 ;
        RECT -258.615 6.475 -258.445 6.645 ;
        RECT -258.155 6.475 -257.985 6.645 ;
        RECT -257.695 6.475 -257.525 6.645 ;
        RECT -257.235 6.475 -257.065 6.645 ;
        RECT -250.075 6.475 -249.905 6.645 ;
        RECT -249.615 6.475 -249.445 6.645 ;
        RECT -249.155 6.475 -248.985 6.645 ;
        RECT -248.695 6.475 -248.525 6.645 ;
        RECT -248.235 6.475 -248.065 6.645 ;
        RECT -247.775 6.475 -247.605 6.645 ;
        RECT -247.315 6.475 -247.145 6.645 ;
        RECT -240.155 6.475 -239.985 6.645 ;
        RECT -239.695 6.475 -239.525 6.645 ;
        RECT -239.235 6.475 -239.065 6.645 ;
        RECT -238.775 6.475 -238.605 6.645 ;
        RECT -238.315 6.475 -238.145 6.645 ;
        RECT -237.855 6.475 -237.685 6.645 ;
        RECT -237.395 6.475 -237.225 6.645 ;
        RECT -230.235 6.475 -230.065 6.645 ;
        RECT -229.775 6.475 -229.605 6.645 ;
        RECT -229.315 6.475 -229.145 6.645 ;
        RECT -228.855 6.475 -228.685 6.645 ;
        RECT -228.395 6.475 -228.225 6.645 ;
        RECT -227.935 6.475 -227.765 6.645 ;
        RECT -227.475 6.475 -227.305 6.645 ;
        RECT -220.315 6.475 -220.145 6.645 ;
        RECT -219.855 6.475 -219.685 6.645 ;
        RECT -219.395 6.475 -219.225 6.645 ;
        RECT -218.935 6.475 -218.765 6.645 ;
        RECT -218.475 6.475 -218.305 6.645 ;
        RECT -218.015 6.475 -217.845 6.645 ;
        RECT -217.555 6.475 -217.385 6.645 ;
        RECT -210.395 6.475 -210.225 6.645 ;
        RECT -209.935 6.475 -209.765 6.645 ;
        RECT -209.475 6.475 -209.305 6.645 ;
        RECT -209.015 6.475 -208.845 6.645 ;
        RECT -208.555 6.475 -208.385 6.645 ;
        RECT -208.095 6.475 -207.925 6.645 ;
        RECT -207.635 6.475 -207.465 6.645 ;
        RECT -200.475 6.475 -200.305 6.645 ;
        RECT -200.015 6.475 -199.845 6.645 ;
        RECT -199.555 6.475 -199.385 6.645 ;
        RECT -199.095 6.475 -198.925 6.645 ;
        RECT -198.635 6.475 -198.465 6.645 ;
        RECT -198.175 6.475 -198.005 6.645 ;
        RECT -197.715 6.475 -197.545 6.645 ;
        RECT -190.555 6.475 -190.385 6.645 ;
        RECT -190.095 6.475 -189.925 6.645 ;
        RECT -189.635 6.475 -189.465 6.645 ;
        RECT -189.175 6.475 -189.005 6.645 ;
        RECT -188.715 6.475 -188.545 6.645 ;
        RECT -188.255 6.475 -188.085 6.645 ;
        RECT -187.795 6.475 -187.625 6.645 ;
        RECT -180.635 6.475 -180.465 6.645 ;
        RECT -180.175 6.475 -180.005 6.645 ;
        RECT -179.715 6.475 -179.545 6.645 ;
        RECT -179.255 6.475 -179.085 6.645 ;
        RECT -178.795 6.475 -178.625 6.645 ;
        RECT -178.335 6.475 -178.165 6.645 ;
        RECT -177.875 6.475 -177.705 6.645 ;
        RECT -170.715 6.475 -170.545 6.645 ;
        RECT -170.255 6.475 -170.085 6.645 ;
        RECT -169.795 6.475 -169.625 6.645 ;
        RECT -169.335 6.475 -169.165 6.645 ;
        RECT -168.875 6.475 -168.705 6.645 ;
        RECT -168.415 6.475 -168.245 6.645 ;
        RECT -167.955 6.475 -167.785 6.645 ;
        RECT -160.795 6.475 -160.625 6.645 ;
        RECT -160.335 6.475 -160.165 6.645 ;
        RECT -159.875 6.475 -159.705 6.645 ;
        RECT -159.415 6.475 -159.245 6.645 ;
        RECT -158.955 6.475 -158.785 6.645 ;
        RECT -158.495 6.475 -158.325 6.645 ;
        RECT -158.035 6.475 -157.865 6.645 ;
        RECT -150.875 6.475 -150.705 6.645 ;
        RECT -150.415 6.475 -150.245 6.645 ;
        RECT -149.955 6.475 -149.785 6.645 ;
        RECT -149.495 6.475 -149.325 6.645 ;
        RECT -149.035 6.475 -148.865 6.645 ;
        RECT -148.575 6.475 -148.405 6.645 ;
        RECT -148.115 6.475 -147.945 6.645 ;
        RECT -140.955 6.475 -140.785 6.645 ;
        RECT -140.495 6.475 -140.325 6.645 ;
        RECT -140.035 6.475 -139.865 6.645 ;
        RECT -139.575 6.475 -139.405 6.645 ;
        RECT -139.115 6.475 -138.945 6.645 ;
        RECT -138.655 6.475 -138.485 6.645 ;
        RECT -138.195 6.475 -138.025 6.645 ;
        RECT -131.035 6.475 -130.865 6.645 ;
        RECT -130.575 6.475 -130.405 6.645 ;
        RECT -130.115 6.475 -129.945 6.645 ;
        RECT -129.655 6.475 -129.485 6.645 ;
        RECT -129.195 6.475 -129.025 6.645 ;
        RECT -128.735 6.475 -128.565 6.645 ;
        RECT -128.275 6.475 -128.105 6.645 ;
        RECT -121.115 6.475 -120.945 6.645 ;
        RECT -120.655 6.475 -120.485 6.645 ;
        RECT -120.195 6.475 -120.025 6.645 ;
        RECT -119.735 6.475 -119.565 6.645 ;
        RECT -119.275 6.475 -119.105 6.645 ;
        RECT -118.815 6.475 -118.645 6.645 ;
        RECT -118.355 6.475 -118.185 6.645 ;
        RECT -111.195 6.475 -111.025 6.645 ;
        RECT -110.735 6.475 -110.565 6.645 ;
        RECT -110.275 6.475 -110.105 6.645 ;
        RECT -109.815 6.475 -109.645 6.645 ;
        RECT -109.355 6.475 -109.185 6.645 ;
        RECT -108.895 6.475 -108.725 6.645 ;
        RECT -108.435 6.475 -108.265 6.645 ;
        RECT -101.275 6.475 -101.105 6.645 ;
        RECT -100.815 6.475 -100.645 6.645 ;
        RECT -100.355 6.475 -100.185 6.645 ;
        RECT -99.895 6.475 -99.725 6.645 ;
        RECT -99.435 6.475 -99.265 6.645 ;
        RECT -98.975 6.475 -98.805 6.645 ;
        RECT -98.515 6.475 -98.345 6.645 ;
        RECT -91.355 6.475 -91.185 6.645 ;
        RECT -90.895 6.475 -90.725 6.645 ;
        RECT -90.435 6.475 -90.265 6.645 ;
        RECT -89.975 6.475 -89.805 6.645 ;
        RECT -89.515 6.475 -89.345 6.645 ;
        RECT -89.055 6.475 -88.885 6.645 ;
        RECT -88.595 6.475 -88.425 6.645 ;
        RECT -81.435 6.475 -81.265 6.645 ;
        RECT -80.975 6.475 -80.805 6.645 ;
        RECT -80.515 6.475 -80.345 6.645 ;
        RECT -80.055 6.475 -79.885 6.645 ;
        RECT -79.595 6.475 -79.425 6.645 ;
        RECT -79.135 6.475 -78.965 6.645 ;
        RECT -78.675 6.475 -78.505 6.645 ;
        RECT -71.515 6.475 -71.345 6.645 ;
        RECT -71.055 6.475 -70.885 6.645 ;
        RECT -70.595 6.475 -70.425 6.645 ;
        RECT -70.135 6.475 -69.965 6.645 ;
        RECT -69.675 6.475 -69.505 6.645 ;
        RECT -69.215 6.475 -69.045 6.645 ;
        RECT -68.755 6.475 -68.585 6.645 ;
        RECT -61.595 6.475 -61.425 6.645 ;
        RECT -61.135 6.475 -60.965 6.645 ;
        RECT -60.675 6.475 -60.505 6.645 ;
        RECT -60.215 6.475 -60.045 6.645 ;
        RECT -59.755 6.475 -59.585 6.645 ;
        RECT -59.295 6.475 -59.125 6.645 ;
        RECT -58.835 6.475 -58.665 6.645 ;
        RECT -51.675 6.475 -51.505 6.645 ;
        RECT -51.215 6.475 -51.045 6.645 ;
        RECT -50.755 6.475 -50.585 6.645 ;
        RECT -50.295 6.475 -50.125 6.645 ;
        RECT -49.835 6.475 -49.665 6.645 ;
        RECT -49.375 6.475 -49.205 6.645 ;
        RECT -48.915 6.475 -48.745 6.645 ;
        RECT -41.755 6.475 -41.585 6.645 ;
        RECT -41.295 6.475 -41.125 6.645 ;
        RECT -40.835 6.475 -40.665 6.645 ;
        RECT -40.375 6.475 -40.205 6.645 ;
        RECT -39.915 6.475 -39.745 6.645 ;
        RECT -39.455 6.475 -39.285 6.645 ;
        RECT -38.995 6.475 -38.825 6.645 ;
        RECT -31.835 6.475 -31.665 6.645 ;
        RECT -31.375 6.475 -31.205 6.645 ;
        RECT -30.915 6.475 -30.745 6.645 ;
        RECT -30.455 6.475 -30.285 6.645 ;
        RECT -29.995 6.475 -29.825 6.645 ;
        RECT -29.535 6.475 -29.365 6.645 ;
        RECT -29.075 6.475 -28.905 6.645 ;
        RECT -21.915 6.475 -21.745 6.645 ;
        RECT -21.455 6.475 -21.285 6.645 ;
        RECT -20.995 6.475 -20.825 6.645 ;
        RECT -20.535 6.475 -20.365 6.645 ;
        RECT -20.075 6.475 -19.905 6.645 ;
        RECT -19.615 6.475 -19.445 6.645 ;
        RECT -19.155 6.475 -18.985 6.645 ;
        RECT -11.995 6.475 -11.825 6.645 ;
        RECT -11.535 6.475 -11.365 6.645 ;
        RECT -11.075 6.475 -10.905 6.645 ;
        RECT -10.615 6.475 -10.445 6.645 ;
        RECT -10.155 6.475 -9.985 6.645 ;
        RECT -9.695 6.475 -9.525 6.645 ;
        RECT -9.235 6.475 -9.065 6.645 ;
        RECT -2.075 6.475 -1.905 6.645 ;
        RECT -1.615 6.475 -1.445 6.645 ;
        RECT -1.155 6.475 -0.985 6.645 ;
        RECT -0.695 6.475 -0.525 6.645 ;
        RECT -0.235 6.475 -0.065 6.645 ;
        RECT 0.225 6.475 0.395 6.645 ;
        RECT 0.685 6.475 0.855 6.645 ;
        RECT 7.845 6.475 8.015 6.645 ;
        RECT 8.305 6.475 8.475 6.645 ;
        RECT 8.765 6.475 8.935 6.645 ;
        RECT 9.225 6.475 9.395 6.645 ;
        RECT 9.685 6.475 9.855 6.645 ;
        RECT 10.145 6.475 10.315 6.645 ;
        RECT 10.605 6.475 10.775 6.645 ;
        RECT 17.765 6.475 17.935 6.645 ;
        RECT 18.225 6.475 18.395 6.645 ;
        RECT 18.685 6.475 18.855 6.645 ;
        RECT 19.145 6.475 19.315 6.645 ;
        RECT 19.605 6.475 19.775 6.645 ;
        RECT 20.065 6.475 20.235 6.645 ;
        RECT 20.525 6.475 20.695 6.645 ;
        RECT -285.185 5.815 -285.015 5.985 ;
        RECT -285.185 5.355 -285.015 5.525 ;
        RECT -281.645 5.815 -281.475 5.985 ;
        RECT -275.265 5.815 -275.095 5.985 ;
        RECT -281.645 5.355 -281.475 5.525 ;
        RECT -275.265 5.355 -275.095 5.525 ;
        RECT -283.415 5.085 -283.245 5.255 ;
        RECT -285.185 4.895 -285.015 5.065 ;
        RECT -281.645 4.895 -281.475 5.065 ;
        RECT -271.725 5.815 -271.555 5.985 ;
        RECT -265.345 5.815 -265.175 5.985 ;
        RECT -271.725 5.355 -271.555 5.525 ;
        RECT -265.345 5.355 -265.175 5.525 ;
        RECT -273.495 5.085 -273.325 5.255 ;
        RECT -275.265 4.895 -275.095 5.065 ;
        RECT -271.725 4.895 -271.555 5.065 ;
        RECT -261.805 5.815 -261.635 5.985 ;
        RECT -255.425 5.815 -255.255 5.985 ;
        RECT -261.805 5.355 -261.635 5.525 ;
        RECT -255.425 5.355 -255.255 5.525 ;
        RECT -263.575 5.085 -263.405 5.255 ;
        RECT -265.345 4.895 -265.175 5.065 ;
        RECT -261.805 4.895 -261.635 5.065 ;
        RECT -251.885 5.815 -251.715 5.985 ;
        RECT -245.505 5.815 -245.335 5.985 ;
        RECT -251.885 5.355 -251.715 5.525 ;
        RECT -245.505 5.355 -245.335 5.525 ;
        RECT -253.655 5.085 -253.485 5.255 ;
        RECT -255.425 4.895 -255.255 5.065 ;
        RECT -251.885 4.895 -251.715 5.065 ;
        RECT -241.965 5.815 -241.795 5.985 ;
        RECT -235.585 5.815 -235.415 5.985 ;
        RECT -241.965 5.355 -241.795 5.525 ;
        RECT -235.585 5.355 -235.415 5.525 ;
        RECT -243.735 5.085 -243.565 5.255 ;
        RECT -245.505 4.895 -245.335 5.065 ;
        RECT -241.965 4.895 -241.795 5.065 ;
        RECT -232.045 5.815 -231.875 5.985 ;
        RECT -225.665 5.815 -225.495 5.985 ;
        RECT -232.045 5.355 -231.875 5.525 ;
        RECT -225.665 5.355 -225.495 5.525 ;
        RECT -233.815 5.085 -233.645 5.255 ;
        RECT -235.585 4.895 -235.415 5.065 ;
        RECT -232.045 4.895 -231.875 5.065 ;
        RECT -222.125 5.815 -221.955 5.985 ;
        RECT -215.745 5.815 -215.575 5.985 ;
        RECT -222.125 5.355 -221.955 5.525 ;
        RECT -215.745 5.355 -215.575 5.525 ;
        RECT -223.895 5.085 -223.725 5.255 ;
        RECT -225.665 4.895 -225.495 5.065 ;
        RECT -222.125 4.895 -221.955 5.065 ;
        RECT -212.205 5.815 -212.035 5.985 ;
        RECT -205.825 5.815 -205.655 5.985 ;
        RECT -212.205 5.355 -212.035 5.525 ;
        RECT -205.825 5.355 -205.655 5.525 ;
        RECT -213.975 5.085 -213.805 5.255 ;
        RECT -215.745 4.895 -215.575 5.065 ;
        RECT -212.205 4.895 -212.035 5.065 ;
        RECT -202.285 5.815 -202.115 5.985 ;
        RECT -195.905 5.815 -195.735 5.985 ;
        RECT -202.285 5.355 -202.115 5.525 ;
        RECT -195.905 5.355 -195.735 5.525 ;
        RECT -204.055 5.085 -203.885 5.255 ;
        RECT -205.825 4.895 -205.655 5.065 ;
        RECT -202.285 4.895 -202.115 5.065 ;
        RECT -192.365 5.815 -192.195 5.985 ;
        RECT -185.985 5.815 -185.815 5.985 ;
        RECT -192.365 5.355 -192.195 5.525 ;
        RECT -185.985 5.355 -185.815 5.525 ;
        RECT -194.135 5.085 -193.965 5.255 ;
        RECT -195.905 4.895 -195.735 5.065 ;
        RECT -192.365 4.895 -192.195 5.065 ;
        RECT -182.445 5.815 -182.275 5.985 ;
        RECT -176.065 5.815 -175.895 5.985 ;
        RECT -182.445 5.355 -182.275 5.525 ;
        RECT -176.065 5.355 -175.895 5.525 ;
        RECT -184.215 5.085 -184.045 5.255 ;
        RECT -185.985 4.895 -185.815 5.065 ;
        RECT -182.445 4.895 -182.275 5.065 ;
        RECT -172.525 5.815 -172.355 5.985 ;
        RECT -166.145 5.815 -165.975 5.985 ;
        RECT -172.525 5.355 -172.355 5.525 ;
        RECT -166.145 5.355 -165.975 5.525 ;
        RECT -174.295 5.085 -174.125 5.255 ;
        RECT -176.065 4.895 -175.895 5.065 ;
        RECT -172.525 4.895 -172.355 5.065 ;
        RECT -162.605 5.815 -162.435 5.985 ;
        RECT -156.225 5.815 -156.055 5.985 ;
        RECT -162.605 5.355 -162.435 5.525 ;
        RECT -156.225 5.355 -156.055 5.525 ;
        RECT -164.375 5.085 -164.205 5.255 ;
        RECT -166.145 4.895 -165.975 5.065 ;
        RECT -162.605 4.895 -162.435 5.065 ;
        RECT -152.685 5.815 -152.515 5.985 ;
        RECT -146.305 5.815 -146.135 5.985 ;
        RECT -152.685 5.355 -152.515 5.525 ;
        RECT -146.305 5.355 -146.135 5.525 ;
        RECT -154.455 5.085 -154.285 5.255 ;
        RECT -156.225 4.895 -156.055 5.065 ;
        RECT -152.685 4.895 -152.515 5.065 ;
        RECT -142.765 5.815 -142.595 5.985 ;
        RECT -136.385 5.815 -136.215 5.985 ;
        RECT -142.765 5.355 -142.595 5.525 ;
        RECT -136.385 5.355 -136.215 5.525 ;
        RECT -144.535 5.085 -144.365 5.255 ;
        RECT -146.305 4.895 -146.135 5.065 ;
        RECT -142.765 4.895 -142.595 5.065 ;
        RECT -132.845 5.815 -132.675 5.985 ;
        RECT -126.465 5.815 -126.295 5.985 ;
        RECT -132.845 5.355 -132.675 5.525 ;
        RECT -126.465 5.355 -126.295 5.525 ;
        RECT -134.615 5.085 -134.445 5.255 ;
        RECT -136.385 4.895 -136.215 5.065 ;
        RECT -132.845 4.895 -132.675 5.065 ;
        RECT -122.925 5.815 -122.755 5.985 ;
        RECT -116.545 5.815 -116.375 5.985 ;
        RECT -122.925 5.355 -122.755 5.525 ;
        RECT -116.545 5.355 -116.375 5.525 ;
        RECT -124.695 5.085 -124.525 5.255 ;
        RECT -126.465 4.895 -126.295 5.065 ;
        RECT -122.925 4.895 -122.755 5.065 ;
        RECT -113.005 5.815 -112.835 5.985 ;
        RECT -106.625 5.815 -106.455 5.985 ;
        RECT -113.005 5.355 -112.835 5.525 ;
        RECT -106.625 5.355 -106.455 5.525 ;
        RECT -114.775 5.085 -114.605 5.255 ;
        RECT -116.545 4.895 -116.375 5.065 ;
        RECT -113.005 4.895 -112.835 5.065 ;
        RECT -103.085 5.815 -102.915 5.985 ;
        RECT -96.705 5.815 -96.535 5.985 ;
        RECT -103.085 5.355 -102.915 5.525 ;
        RECT -96.705 5.355 -96.535 5.525 ;
        RECT -104.855 5.085 -104.685 5.255 ;
        RECT -106.625 4.895 -106.455 5.065 ;
        RECT -103.085 4.895 -102.915 5.065 ;
        RECT -93.165 5.815 -92.995 5.985 ;
        RECT -86.785 5.815 -86.615 5.985 ;
        RECT -93.165 5.355 -92.995 5.525 ;
        RECT -86.785 5.355 -86.615 5.525 ;
        RECT -94.935 5.085 -94.765 5.255 ;
        RECT -96.705 4.895 -96.535 5.065 ;
        RECT -93.165 4.895 -92.995 5.065 ;
        RECT -83.245 5.815 -83.075 5.985 ;
        RECT -76.865 5.815 -76.695 5.985 ;
        RECT -83.245 5.355 -83.075 5.525 ;
        RECT -76.865 5.355 -76.695 5.525 ;
        RECT -85.015 5.085 -84.845 5.255 ;
        RECT -86.785 4.895 -86.615 5.065 ;
        RECT -83.245 4.895 -83.075 5.065 ;
        RECT -73.325 5.815 -73.155 5.985 ;
        RECT -66.945 5.815 -66.775 5.985 ;
        RECT -73.325 5.355 -73.155 5.525 ;
        RECT -66.945 5.355 -66.775 5.525 ;
        RECT -75.095 5.085 -74.925 5.255 ;
        RECT -76.865 4.895 -76.695 5.065 ;
        RECT -73.325 4.895 -73.155 5.065 ;
        RECT -63.405 5.815 -63.235 5.985 ;
        RECT -57.025 5.815 -56.855 5.985 ;
        RECT -63.405 5.355 -63.235 5.525 ;
        RECT -57.025 5.355 -56.855 5.525 ;
        RECT -65.175 5.085 -65.005 5.255 ;
        RECT -66.945 4.895 -66.775 5.065 ;
        RECT -63.405 4.895 -63.235 5.065 ;
        RECT -53.485 5.815 -53.315 5.985 ;
        RECT -47.105 5.815 -46.935 5.985 ;
        RECT -53.485 5.355 -53.315 5.525 ;
        RECT -47.105 5.355 -46.935 5.525 ;
        RECT -55.255 5.085 -55.085 5.255 ;
        RECT -57.025 4.895 -56.855 5.065 ;
        RECT -53.485 4.895 -53.315 5.065 ;
        RECT -43.565 5.815 -43.395 5.985 ;
        RECT -37.185 5.815 -37.015 5.985 ;
        RECT -43.565 5.355 -43.395 5.525 ;
        RECT -37.185 5.355 -37.015 5.525 ;
        RECT -45.335 5.085 -45.165 5.255 ;
        RECT -47.105 4.895 -46.935 5.065 ;
        RECT -43.565 4.895 -43.395 5.065 ;
        RECT -33.645 5.815 -33.475 5.985 ;
        RECT -27.265 5.815 -27.095 5.985 ;
        RECT -33.645 5.355 -33.475 5.525 ;
        RECT -27.265 5.355 -27.095 5.525 ;
        RECT -35.415 5.085 -35.245 5.255 ;
        RECT -37.185 4.895 -37.015 5.065 ;
        RECT -33.645 4.895 -33.475 5.065 ;
        RECT -23.725 5.815 -23.555 5.985 ;
        RECT -17.345 5.815 -17.175 5.985 ;
        RECT -23.725 5.355 -23.555 5.525 ;
        RECT -17.345 5.355 -17.175 5.525 ;
        RECT -25.495 5.085 -25.325 5.255 ;
        RECT -27.265 4.895 -27.095 5.065 ;
        RECT -23.725 4.895 -23.555 5.065 ;
        RECT -13.805 5.815 -13.635 5.985 ;
        RECT -7.425 5.815 -7.255 5.985 ;
        RECT -13.805 5.355 -13.635 5.525 ;
        RECT -7.425 5.355 -7.255 5.525 ;
        RECT -15.575 5.085 -15.405 5.255 ;
        RECT -17.345 4.895 -17.175 5.065 ;
        RECT -13.805 4.895 -13.635 5.065 ;
        RECT -3.885 5.815 -3.715 5.985 ;
        RECT 2.495 5.815 2.665 5.985 ;
        RECT -3.885 5.355 -3.715 5.525 ;
        RECT 2.495 5.355 2.665 5.525 ;
        RECT -5.655 5.085 -5.485 5.255 ;
        RECT -7.425 4.895 -7.255 5.065 ;
        RECT -3.885 4.895 -3.715 5.065 ;
        RECT 6.035 5.815 6.205 5.985 ;
        RECT 12.415 5.815 12.585 5.985 ;
        RECT 6.035 5.355 6.205 5.525 ;
        RECT 12.415 5.355 12.585 5.525 ;
        RECT 4.265 5.085 4.435 5.255 ;
        RECT 2.495 4.895 2.665 5.065 ;
        RECT 6.035 4.895 6.205 5.065 ;
        RECT 15.955 5.815 16.125 5.985 ;
        RECT 15.955 5.355 16.125 5.525 ;
        RECT 14.185 5.085 14.355 5.255 ;
        RECT 12.415 4.895 12.585 5.065 ;
        RECT 15.955 4.895 16.125 5.065 ;
        RECT -289.785 -78.175 -289.615 -78.005 ;
        RECT -288.015 -78.275 -287.845 -78.105 ;
        RECT -286.245 -78.175 -286.075 -78.005 ;
        RECT -289.785 -78.635 -289.615 -78.465 ;
        RECT -289.785 -79.095 -289.615 -78.925 ;
        RECT -279.865 -78.175 -279.695 -78.005 ;
        RECT -278.095 -78.275 -277.925 -78.105 ;
        RECT -276.325 -78.175 -276.155 -78.005 ;
        RECT -286.245 -78.635 -286.075 -78.465 ;
        RECT -279.865 -78.635 -279.695 -78.465 ;
        RECT -286.245 -79.095 -286.075 -78.925 ;
        RECT -279.865 -79.095 -279.695 -78.925 ;
        RECT -269.945 -78.175 -269.775 -78.005 ;
        RECT -268.175 -78.275 -268.005 -78.105 ;
        RECT -266.405 -78.175 -266.235 -78.005 ;
        RECT -276.325 -78.635 -276.155 -78.465 ;
        RECT -269.945 -78.635 -269.775 -78.465 ;
        RECT -276.325 -79.095 -276.155 -78.925 ;
        RECT -269.945 -79.095 -269.775 -78.925 ;
        RECT -260.025 -78.175 -259.855 -78.005 ;
        RECT -258.255 -78.275 -258.085 -78.105 ;
        RECT -256.485 -78.175 -256.315 -78.005 ;
        RECT -266.405 -78.635 -266.235 -78.465 ;
        RECT -260.025 -78.635 -259.855 -78.465 ;
        RECT -266.405 -79.095 -266.235 -78.925 ;
        RECT -260.025 -79.095 -259.855 -78.925 ;
        RECT -250.105 -78.175 -249.935 -78.005 ;
        RECT -248.335 -78.275 -248.165 -78.105 ;
        RECT -246.565 -78.175 -246.395 -78.005 ;
        RECT -256.485 -78.635 -256.315 -78.465 ;
        RECT -250.105 -78.635 -249.935 -78.465 ;
        RECT -256.485 -79.095 -256.315 -78.925 ;
        RECT -250.105 -79.095 -249.935 -78.925 ;
        RECT -240.185 -78.175 -240.015 -78.005 ;
        RECT -238.415 -78.275 -238.245 -78.105 ;
        RECT -236.645 -78.175 -236.475 -78.005 ;
        RECT -246.565 -78.635 -246.395 -78.465 ;
        RECT -240.185 -78.635 -240.015 -78.465 ;
        RECT -246.565 -79.095 -246.395 -78.925 ;
        RECT -240.185 -79.095 -240.015 -78.925 ;
        RECT -230.265 -78.175 -230.095 -78.005 ;
        RECT -228.495 -78.275 -228.325 -78.105 ;
        RECT -226.725 -78.175 -226.555 -78.005 ;
        RECT -236.645 -78.635 -236.475 -78.465 ;
        RECT -230.265 -78.635 -230.095 -78.465 ;
        RECT -236.645 -79.095 -236.475 -78.925 ;
        RECT -230.265 -79.095 -230.095 -78.925 ;
        RECT -220.345 -78.175 -220.175 -78.005 ;
        RECT -218.575 -78.275 -218.405 -78.105 ;
        RECT -216.805 -78.175 -216.635 -78.005 ;
        RECT -226.725 -78.635 -226.555 -78.465 ;
        RECT -220.345 -78.635 -220.175 -78.465 ;
        RECT -226.725 -79.095 -226.555 -78.925 ;
        RECT -220.345 -79.095 -220.175 -78.925 ;
        RECT -210.425 -78.175 -210.255 -78.005 ;
        RECT -208.655 -78.275 -208.485 -78.105 ;
        RECT -206.885 -78.175 -206.715 -78.005 ;
        RECT -216.805 -78.635 -216.635 -78.465 ;
        RECT -210.425 -78.635 -210.255 -78.465 ;
        RECT -216.805 -79.095 -216.635 -78.925 ;
        RECT -210.425 -79.095 -210.255 -78.925 ;
        RECT -200.505 -78.175 -200.335 -78.005 ;
        RECT -198.735 -78.275 -198.565 -78.105 ;
        RECT -196.965 -78.175 -196.795 -78.005 ;
        RECT -206.885 -78.635 -206.715 -78.465 ;
        RECT -200.505 -78.635 -200.335 -78.465 ;
        RECT -206.885 -79.095 -206.715 -78.925 ;
        RECT -200.505 -79.095 -200.335 -78.925 ;
        RECT -190.585 -78.175 -190.415 -78.005 ;
        RECT -188.815 -78.275 -188.645 -78.105 ;
        RECT -187.045 -78.175 -186.875 -78.005 ;
        RECT -196.965 -78.635 -196.795 -78.465 ;
        RECT -190.585 -78.635 -190.415 -78.465 ;
        RECT -196.965 -79.095 -196.795 -78.925 ;
        RECT -190.585 -79.095 -190.415 -78.925 ;
        RECT -180.665 -78.175 -180.495 -78.005 ;
        RECT -178.895 -78.275 -178.725 -78.105 ;
        RECT -177.125 -78.175 -176.955 -78.005 ;
        RECT -187.045 -78.635 -186.875 -78.465 ;
        RECT -180.665 -78.635 -180.495 -78.465 ;
        RECT -187.045 -79.095 -186.875 -78.925 ;
        RECT -180.665 -79.095 -180.495 -78.925 ;
        RECT -170.745 -78.175 -170.575 -78.005 ;
        RECT -168.975 -78.275 -168.805 -78.105 ;
        RECT -167.205 -78.175 -167.035 -78.005 ;
        RECT -177.125 -78.635 -176.955 -78.465 ;
        RECT -170.745 -78.635 -170.575 -78.465 ;
        RECT -177.125 -79.095 -176.955 -78.925 ;
        RECT -170.745 -79.095 -170.575 -78.925 ;
        RECT -160.825 -78.175 -160.655 -78.005 ;
        RECT -159.055 -78.275 -158.885 -78.105 ;
        RECT -157.285 -78.175 -157.115 -78.005 ;
        RECT -167.205 -78.635 -167.035 -78.465 ;
        RECT -160.825 -78.635 -160.655 -78.465 ;
        RECT -167.205 -79.095 -167.035 -78.925 ;
        RECT -160.825 -79.095 -160.655 -78.925 ;
        RECT -150.905 -78.175 -150.735 -78.005 ;
        RECT -149.135 -78.275 -148.965 -78.105 ;
        RECT -147.365 -78.175 -147.195 -78.005 ;
        RECT -157.285 -78.635 -157.115 -78.465 ;
        RECT -150.905 -78.635 -150.735 -78.465 ;
        RECT -157.285 -79.095 -157.115 -78.925 ;
        RECT -150.905 -79.095 -150.735 -78.925 ;
        RECT -140.985 -78.175 -140.815 -78.005 ;
        RECT -139.215 -78.275 -139.045 -78.105 ;
        RECT -137.445 -78.175 -137.275 -78.005 ;
        RECT -147.365 -78.635 -147.195 -78.465 ;
        RECT -140.985 -78.635 -140.815 -78.465 ;
        RECT -147.365 -79.095 -147.195 -78.925 ;
        RECT -140.985 -79.095 -140.815 -78.925 ;
        RECT -131.065 -78.175 -130.895 -78.005 ;
        RECT -129.295 -78.275 -129.125 -78.105 ;
        RECT -127.525 -78.175 -127.355 -78.005 ;
        RECT -137.445 -78.635 -137.275 -78.465 ;
        RECT -131.065 -78.635 -130.895 -78.465 ;
        RECT -137.445 -79.095 -137.275 -78.925 ;
        RECT -131.065 -79.095 -130.895 -78.925 ;
        RECT -121.145 -78.175 -120.975 -78.005 ;
        RECT -119.375 -78.275 -119.205 -78.105 ;
        RECT -117.605 -78.175 -117.435 -78.005 ;
        RECT -127.525 -78.635 -127.355 -78.465 ;
        RECT -121.145 -78.635 -120.975 -78.465 ;
        RECT -127.525 -79.095 -127.355 -78.925 ;
        RECT -121.145 -79.095 -120.975 -78.925 ;
        RECT -111.225 -78.175 -111.055 -78.005 ;
        RECT -109.455 -78.275 -109.285 -78.105 ;
        RECT -107.685 -78.175 -107.515 -78.005 ;
        RECT -117.605 -78.635 -117.435 -78.465 ;
        RECT -111.225 -78.635 -111.055 -78.465 ;
        RECT -117.605 -79.095 -117.435 -78.925 ;
        RECT -111.225 -79.095 -111.055 -78.925 ;
        RECT -101.305 -78.175 -101.135 -78.005 ;
        RECT -99.535 -78.275 -99.365 -78.105 ;
        RECT -97.765 -78.175 -97.595 -78.005 ;
        RECT -107.685 -78.635 -107.515 -78.465 ;
        RECT -101.305 -78.635 -101.135 -78.465 ;
        RECT -107.685 -79.095 -107.515 -78.925 ;
        RECT -101.305 -79.095 -101.135 -78.925 ;
        RECT -91.385 -78.175 -91.215 -78.005 ;
        RECT -89.615 -78.275 -89.445 -78.105 ;
        RECT -87.845 -78.175 -87.675 -78.005 ;
        RECT -97.765 -78.635 -97.595 -78.465 ;
        RECT -91.385 -78.635 -91.215 -78.465 ;
        RECT -97.765 -79.095 -97.595 -78.925 ;
        RECT -91.385 -79.095 -91.215 -78.925 ;
        RECT -81.465 -78.175 -81.295 -78.005 ;
        RECT -79.695 -78.275 -79.525 -78.105 ;
        RECT -77.925 -78.175 -77.755 -78.005 ;
        RECT -87.845 -78.635 -87.675 -78.465 ;
        RECT -81.465 -78.635 -81.295 -78.465 ;
        RECT -87.845 -79.095 -87.675 -78.925 ;
        RECT -81.465 -79.095 -81.295 -78.925 ;
        RECT -71.545 -78.175 -71.375 -78.005 ;
        RECT -69.775 -78.275 -69.605 -78.105 ;
        RECT -68.005 -78.175 -67.835 -78.005 ;
        RECT -77.925 -78.635 -77.755 -78.465 ;
        RECT -71.545 -78.635 -71.375 -78.465 ;
        RECT -77.925 -79.095 -77.755 -78.925 ;
        RECT -71.545 -79.095 -71.375 -78.925 ;
        RECT -61.625 -78.175 -61.455 -78.005 ;
        RECT -59.855 -78.275 -59.685 -78.105 ;
        RECT -58.085 -78.175 -57.915 -78.005 ;
        RECT -68.005 -78.635 -67.835 -78.465 ;
        RECT -61.625 -78.635 -61.455 -78.465 ;
        RECT -68.005 -79.095 -67.835 -78.925 ;
        RECT -61.625 -79.095 -61.455 -78.925 ;
        RECT -51.705 -78.175 -51.535 -78.005 ;
        RECT -49.935 -78.275 -49.765 -78.105 ;
        RECT -48.165 -78.175 -47.995 -78.005 ;
        RECT -58.085 -78.635 -57.915 -78.465 ;
        RECT -51.705 -78.635 -51.535 -78.465 ;
        RECT -58.085 -79.095 -57.915 -78.925 ;
        RECT -51.705 -79.095 -51.535 -78.925 ;
        RECT -41.785 -78.175 -41.615 -78.005 ;
        RECT -40.015 -78.275 -39.845 -78.105 ;
        RECT -38.245 -78.175 -38.075 -78.005 ;
        RECT -48.165 -78.635 -47.995 -78.465 ;
        RECT -41.785 -78.635 -41.615 -78.465 ;
        RECT -48.165 -79.095 -47.995 -78.925 ;
        RECT -41.785 -79.095 -41.615 -78.925 ;
        RECT -31.865 -78.175 -31.695 -78.005 ;
        RECT -30.095 -78.275 -29.925 -78.105 ;
        RECT -28.325 -78.175 -28.155 -78.005 ;
        RECT -38.245 -78.635 -38.075 -78.465 ;
        RECT -31.865 -78.635 -31.695 -78.465 ;
        RECT -38.245 -79.095 -38.075 -78.925 ;
        RECT -31.865 -79.095 -31.695 -78.925 ;
        RECT -21.945 -78.175 -21.775 -78.005 ;
        RECT -20.175 -78.275 -20.005 -78.105 ;
        RECT -18.405 -78.175 -18.235 -78.005 ;
        RECT -28.325 -78.635 -28.155 -78.465 ;
        RECT -21.945 -78.635 -21.775 -78.465 ;
        RECT -28.325 -79.095 -28.155 -78.925 ;
        RECT -21.945 -79.095 -21.775 -78.925 ;
        RECT -12.025 -78.175 -11.855 -78.005 ;
        RECT -10.255 -78.275 -10.085 -78.105 ;
        RECT -8.485 -78.175 -8.315 -78.005 ;
        RECT -18.405 -78.635 -18.235 -78.465 ;
        RECT -12.025 -78.635 -11.855 -78.465 ;
        RECT -18.405 -79.095 -18.235 -78.925 ;
        RECT -12.025 -79.095 -11.855 -78.925 ;
        RECT -2.105 -78.175 -1.935 -78.005 ;
        RECT -0.335 -78.275 -0.165 -78.105 ;
        RECT 1.435 -78.175 1.605 -78.005 ;
        RECT -8.485 -78.635 -8.315 -78.465 ;
        RECT -2.105 -78.635 -1.935 -78.465 ;
        RECT -8.485 -79.095 -8.315 -78.925 ;
        RECT -2.105 -79.095 -1.935 -78.925 ;
        RECT 7.815 -78.175 7.985 -78.005 ;
        RECT 9.585 -78.275 9.755 -78.105 ;
        RECT 11.355 -78.175 11.525 -78.005 ;
        RECT 1.435 -78.635 1.605 -78.465 ;
        RECT 7.815 -78.635 7.985 -78.465 ;
        RECT 1.435 -79.095 1.605 -78.925 ;
        RECT 7.815 -79.095 7.985 -78.925 ;
        RECT 17.735 -78.175 17.905 -78.005 ;
        RECT 19.505 -78.275 19.675 -78.105 ;
        RECT 21.275 -78.175 21.445 -78.005 ;
        RECT 11.355 -78.635 11.525 -78.465 ;
        RECT 17.735 -78.635 17.905 -78.465 ;
        RECT 11.355 -79.095 11.525 -78.925 ;
        RECT 17.735 -79.095 17.905 -78.925 ;
        RECT 21.275 -78.635 21.445 -78.465 ;
        RECT 21.275 -79.095 21.445 -78.925 ;
        RECT -284.435 -79.755 -284.265 -79.585 ;
        RECT -283.975 -79.755 -283.805 -79.585 ;
        RECT -283.515 -79.755 -283.345 -79.585 ;
        RECT -283.055 -79.755 -282.885 -79.585 ;
        RECT -282.595 -79.755 -282.425 -79.585 ;
        RECT -282.135 -79.755 -281.965 -79.585 ;
        RECT -281.675 -79.755 -281.505 -79.585 ;
        RECT -274.515 -79.755 -274.345 -79.585 ;
        RECT -274.055 -79.755 -273.885 -79.585 ;
        RECT -273.595 -79.755 -273.425 -79.585 ;
        RECT -273.135 -79.755 -272.965 -79.585 ;
        RECT -272.675 -79.755 -272.505 -79.585 ;
        RECT -272.215 -79.755 -272.045 -79.585 ;
        RECT -271.755 -79.755 -271.585 -79.585 ;
        RECT -264.595 -79.755 -264.425 -79.585 ;
        RECT -264.135 -79.755 -263.965 -79.585 ;
        RECT -263.675 -79.755 -263.505 -79.585 ;
        RECT -263.215 -79.755 -263.045 -79.585 ;
        RECT -262.755 -79.755 -262.585 -79.585 ;
        RECT -262.295 -79.755 -262.125 -79.585 ;
        RECT -261.835 -79.755 -261.665 -79.585 ;
        RECT -254.675 -79.755 -254.505 -79.585 ;
        RECT -254.215 -79.755 -254.045 -79.585 ;
        RECT -253.755 -79.755 -253.585 -79.585 ;
        RECT -253.295 -79.755 -253.125 -79.585 ;
        RECT -252.835 -79.755 -252.665 -79.585 ;
        RECT -252.375 -79.755 -252.205 -79.585 ;
        RECT -251.915 -79.755 -251.745 -79.585 ;
        RECT -244.755 -79.755 -244.585 -79.585 ;
        RECT -244.295 -79.755 -244.125 -79.585 ;
        RECT -243.835 -79.755 -243.665 -79.585 ;
        RECT -243.375 -79.755 -243.205 -79.585 ;
        RECT -242.915 -79.755 -242.745 -79.585 ;
        RECT -242.455 -79.755 -242.285 -79.585 ;
        RECT -241.995 -79.755 -241.825 -79.585 ;
        RECT -234.835 -79.755 -234.665 -79.585 ;
        RECT -234.375 -79.755 -234.205 -79.585 ;
        RECT -233.915 -79.755 -233.745 -79.585 ;
        RECT -233.455 -79.755 -233.285 -79.585 ;
        RECT -232.995 -79.755 -232.825 -79.585 ;
        RECT -232.535 -79.755 -232.365 -79.585 ;
        RECT -232.075 -79.755 -231.905 -79.585 ;
        RECT -224.915 -79.755 -224.745 -79.585 ;
        RECT -224.455 -79.755 -224.285 -79.585 ;
        RECT -223.995 -79.755 -223.825 -79.585 ;
        RECT -223.535 -79.755 -223.365 -79.585 ;
        RECT -223.075 -79.755 -222.905 -79.585 ;
        RECT -222.615 -79.755 -222.445 -79.585 ;
        RECT -222.155 -79.755 -221.985 -79.585 ;
        RECT -214.995 -79.755 -214.825 -79.585 ;
        RECT -214.535 -79.755 -214.365 -79.585 ;
        RECT -214.075 -79.755 -213.905 -79.585 ;
        RECT -213.615 -79.755 -213.445 -79.585 ;
        RECT -213.155 -79.755 -212.985 -79.585 ;
        RECT -212.695 -79.755 -212.525 -79.585 ;
        RECT -212.235 -79.755 -212.065 -79.585 ;
        RECT -205.075 -79.755 -204.905 -79.585 ;
        RECT -204.615 -79.755 -204.445 -79.585 ;
        RECT -204.155 -79.755 -203.985 -79.585 ;
        RECT -203.695 -79.755 -203.525 -79.585 ;
        RECT -203.235 -79.755 -203.065 -79.585 ;
        RECT -202.775 -79.755 -202.605 -79.585 ;
        RECT -202.315 -79.755 -202.145 -79.585 ;
        RECT -195.155 -79.755 -194.985 -79.585 ;
        RECT -194.695 -79.755 -194.525 -79.585 ;
        RECT -194.235 -79.755 -194.065 -79.585 ;
        RECT -193.775 -79.755 -193.605 -79.585 ;
        RECT -193.315 -79.755 -193.145 -79.585 ;
        RECT -192.855 -79.755 -192.685 -79.585 ;
        RECT -192.395 -79.755 -192.225 -79.585 ;
        RECT -185.235 -79.755 -185.065 -79.585 ;
        RECT -184.775 -79.755 -184.605 -79.585 ;
        RECT -184.315 -79.755 -184.145 -79.585 ;
        RECT -183.855 -79.755 -183.685 -79.585 ;
        RECT -183.395 -79.755 -183.225 -79.585 ;
        RECT -182.935 -79.755 -182.765 -79.585 ;
        RECT -182.475 -79.755 -182.305 -79.585 ;
        RECT -175.315 -79.755 -175.145 -79.585 ;
        RECT -174.855 -79.755 -174.685 -79.585 ;
        RECT -174.395 -79.755 -174.225 -79.585 ;
        RECT -173.935 -79.755 -173.765 -79.585 ;
        RECT -173.475 -79.755 -173.305 -79.585 ;
        RECT -173.015 -79.755 -172.845 -79.585 ;
        RECT -172.555 -79.755 -172.385 -79.585 ;
        RECT -165.395 -79.755 -165.225 -79.585 ;
        RECT -164.935 -79.755 -164.765 -79.585 ;
        RECT -164.475 -79.755 -164.305 -79.585 ;
        RECT -164.015 -79.755 -163.845 -79.585 ;
        RECT -163.555 -79.755 -163.385 -79.585 ;
        RECT -163.095 -79.755 -162.925 -79.585 ;
        RECT -162.635 -79.755 -162.465 -79.585 ;
        RECT -155.475 -79.755 -155.305 -79.585 ;
        RECT -155.015 -79.755 -154.845 -79.585 ;
        RECT -154.555 -79.755 -154.385 -79.585 ;
        RECT -154.095 -79.755 -153.925 -79.585 ;
        RECT -153.635 -79.755 -153.465 -79.585 ;
        RECT -153.175 -79.755 -153.005 -79.585 ;
        RECT -152.715 -79.755 -152.545 -79.585 ;
        RECT -145.555 -79.755 -145.385 -79.585 ;
        RECT -145.095 -79.755 -144.925 -79.585 ;
        RECT -144.635 -79.755 -144.465 -79.585 ;
        RECT -144.175 -79.755 -144.005 -79.585 ;
        RECT -143.715 -79.755 -143.545 -79.585 ;
        RECT -143.255 -79.755 -143.085 -79.585 ;
        RECT -142.795 -79.755 -142.625 -79.585 ;
        RECT -135.635 -79.755 -135.465 -79.585 ;
        RECT -135.175 -79.755 -135.005 -79.585 ;
        RECT -134.715 -79.755 -134.545 -79.585 ;
        RECT -134.255 -79.755 -134.085 -79.585 ;
        RECT -133.795 -79.755 -133.625 -79.585 ;
        RECT -133.335 -79.755 -133.165 -79.585 ;
        RECT -132.875 -79.755 -132.705 -79.585 ;
        RECT -125.715 -79.755 -125.545 -79.585 ;
        RECT -125.255 -79.755 -125.085 -79.585 ;
        RECT -124.795 -79.755 -124.625 -79.585 ;
        RECT -124.335 -79.755 -124.165 -79.585 ;
        RECT -123.875 -79.755 -123.705 -79.585 ;
        RECT -123.415 -79.755 -123.245 -79.585 ;
        RECT -122.955 -79.755 -122.785 -79.585 ;
        RECT -115.795 -79.755 -115.625 -79.585 ;
        RECT -115.335 -79.755 -115.165 -79.585 ;
        RECT -114.875 -79.755 -114.705 -79.585 ;
        RECT -114.415 -79.755 -114.245 -79.585 ;
        RECT -113.955 -79.755 -113.785 -79.585 ;
        RECT -113.495 -79.755 -113.325 -79.585 ;
        RECT -113.035 -79.755 -112.865 -79.585 ;
        RECT -105.875 -79.755 -105.705 -79.585 ;
        RECT -105.415 -79.755 -105.245 -79.585 ;
        RECT -104.955 -79.755 -104.785 -79.585 ;
        RECT -104.495 -79.755 -104.325 -79.585 ;
        RECT -104.035 -79.755 -103.865 -79.585 ;
        RECT -103.575 -79.755 -103.405 -79.585 ;
        RECT -103.115 -79.755 -102.945 -79.585 ;
        RECT -95.955 -79.755 -95.785 -79.585 ;
        RECT -95.495 -79.755 -95.325 -79.585 ;
        RECT -95.035 -79.755 -94.865 -79.585 ;
        RECT -94.575 -79.755 -94.405 -79.585 ;
        RECT -94.115 -79.755 -93.945 -79.585 ;
        RECT -93.655 -79.755 -93.485 -79.585 ;
        RECT -93.195 -79.755 -93.025 -79.585 ;
        RECT -86.035 -79.755 -85.865 -79.585 ;
        RECT -85.575 -79.755 -85.405 -79.585 ;
        RECT -85.115 -79.755 -84.945 -79.585 ;
        RECT -84.655 -79.755 -84.485 -79.585 ;
        RECT -84.195 -79.755 -84.025 -79.585 ;
        RECT -83.735 -79.755 -83.565 -79.585 ;
        RECT -83.275 -79.755 -83.105 -79.585 ;
        RECT -76.115 -79.755 -75.945 -79.585 ;
        RECT -75.655 -79.755 -75.485 -79.585 ;
        RECT -75.195 -79.755 -75.025 -79.585 ;
        RECT -74.735 -79.755 -74.565 -79.585 ;
        RECT -74.275 -79.755 -74.105 -79.585 ;
        RECT -73.815 -79.755 -73.645 -79.585 ;
        RECT -73.355 -79.755 -73.185 -79.585 ;
        RECT -66.195 -79.755 -66.025 -79.585 ;
        RECT -65.735 -79.755 -65.565 -79.585 ;
        RECT -65.275 -79.755 -65.105 -79.585 ;
        RECT -64.815 -79.755 -64.645 -79.585 ;
        RECT -64.355 -79.755 -64.185 -79.585 ;
        RECT -63.895 -79.755 -63.725 -79.585 ;
        RECT -63.435 -79.755 -63.265 -79.585 ;
        RECT -56.275 -79.755 -56.105 -79.585 ;
        RECT -55.815 -79.755 -55.645 -79.585 ;
        RECT -55.355 -79.755 -55.185 -79.585 ;
        RECT -54.895 -79.755 -54.725 -79.585 ;
        RECT -54.435 -79.755 -54.265 -79.585 ;
        RECT -53.975 -79.755 -53.805 -79.585 ;
        RECT -53.515 -79.755 -53.345 -79.585 ;
        RECT -46.355 -79.755 -46.185 -79.585 ;
        RECT -45.895 -79.755 -45.725 -79.585 ;
        RECT -45.435 -79.755 -45.265 -79.585 ;
        RECT -44.975 -79.755 -44.805 -79.585 ;
        RECT -44.515 -79.755 -44.345 -79.585 ;
        RECT -44.055 -79.755 -43.885 -79.585 ;
        RECT -43.595 -79.755 -43.425 -79.585 ;
        RECT -36.435 -79.755 -36.265 -79.585 ;
        RECT -35.975 -79.755 -35.805 -79.585 ;
        RECT -35.515 -79.755 -35.345 -79.585 ;
        RECT -35.055 -79.755 -34.885 -79.585 ;
        RECT -34.595 -79.755 -34.425 -79.585 ;
        RECT -34.135 -79.755 -33.965 -79.585 ;
        RECT -33.675 -79.755 -33.505 -79.585 ;
        RECT -26.515 -79.755 -26.345 -79.585 ;
        RECT -26.055 -79.755 -25.885 -79.585 ;
        RECT -25.595 -79.755 -25.425 -79.585 ;
        RECT -25.135 -79.755 -24.965 -79.585 ;
        RECT -24.675 -79.755 -24.505 -79.585 ;
        RECT -24.215 -79.755 -24.045 -79.585 ;
        RECT -23.755 -79.755 -23.585 -79.585 ;
        RECT -16.595 -79.755 -16.425 -79.585 ;
        RECT -16.135 -79.755 -15.965 -79.585 ;
        RECT -15.675 -79.755 -15.505 -79.585 ;
        RECT -15.215 -79.755 -15.045 -79.585 ;
        RECT -14.755 -79.755 -14.585 -79.585 ;
        RECT -14.295 -79.755 -14.125 -79.585 ;
        RECT -13.835 -79.755 -13.665 -79.585 ;
        RECT -6.675 -79.755 -6.505 -79.585 ;
        RECT -6.215 -79.755 -6.045 -79.585 ;
        RECT -5.755 -79.755 -5.585 -79.585 ;
        RECT -5.295 -79.755 -5.125 -79.585 ;
        RECT -4.835 -79.755 -4.665 -79.585 ;
        RECT -4.375 -79.755 -4.205 -79.585 ;
        RECT -3.915 -79.755 -3.745 -79.585 ;
        RECT 3.245 -79.755 3.415 -79.585 ;
        RECT 3.705 -79.755 3.875 -79.585 ;
        RECT 4.165 -79.755 4.335 -79.585 ;
        RECT 4.625 -79.755 4.795 -79.585 ;
        RECT 5.085 -79.755 5.255 -79.585 ;
        RECT 5.545 -79.755 5.715 -79.585 ;
        RECT 6.005 -79.755 6.175 -79.585 ;
        RECT 13.165 -79.755 13.335 -79.585 ;
        RECT 13.625 -79.755 13.795 -79.585 ;
        RECT 14.085 -79.755 14.255 -79.585 ;
        RECT 14.545 -79.755 14.715 -79.585 ;
        RECT 15.005 -79.755 15.175 -79.585 ;
        RECT 15.465 -79.755 15.635 -79.585 ;
        RECT 15.925 -79.755 16.095 -79.585 ;
        RECT -289.395 -82.475 -289.225 -82.305 ;
        RECT -288.935 -82.475 -288.765 -82.305 ;
        RECT -288.475 -82.475 -288.305 -82.305 ;
        RECT -288.015 -82.475 -287.845 -82.305 ;
        RECT -287.555 -82.475 -287.385 -82.305 ;
        RECT -287.095 -82.475 -286.925 -82.305 ;
        RECT -286.635 -82.475 -286.465 -82.305 ;
        RECT -279.475 -82.475 -279.305 -82.305 ;
        RECT -279.015 -82.475 -278.845 -82.305 ;
        RECT -278.555 -82.475 -278.385 -82.305 ;
        RECT -278.095 -82.475 -277.925 -82.305 ;
        RECT -277.635 -82.475 -277.465 -82.305 ;
        RECT -277.175 -82.475 -277.005 -82.305 ;
        RECT -276.715 -82.475 -276.545 -82.305 ;
        RECT -269.555 -82.475 -269.385 -82.305 ;
        RECT -269.095 -82.475 -268.925 -82.305 ;
        RECT -268.635 -82.475 -268.465 -82.305 ;
        RECT -268.175 -82.475 -268.005 -82.305 ;
        RECT -267.715 -82.475 -267.545 -82.305 ;
        RECT -267.255 -82.475 -267.085 -82.305 ;
        RECT -266.795 -82.475 -266.625 -82.305 ;
        RECT -259.635 -82.475 -259.465 -82.305 ;
        RECT -259.175 -82.475 -259.005 -82.305 ;
        RECT -258.715 -82.475 -258.545 -82.305 ;
        RECT -258.255 -82.475 -258.085 -82.305 ;
        RECT -257.795 -82.475 -257.625 -82.305 ;
        RECT -257.335 -82.475 -257.165 -82.305 ;
        RECT -256.875 -82.475 -256.705 -82.305 ;
        RECT -249.715 -82.475 -249.545 -82.305 ;
        RECT -249.255 -82.475 -249.085 -82.305 ;
        RECT -248.795 -82.475 -248.625 -82.305 ;
        RECT -248.335 -82.475 -248.165 -82.305 ;
        RECT -247.875 -82.475 -247.705 -82.305 ;
        RECT -247.415 -82.475 -247.245 -82.305 ;
        RECT -246.955 -82.475 -246.785 -82.305 ;
        RECT -239.795 -82.475 -239.625 -82.305 ;
        RECT -239.335 -82.475 -239.165 -82.305 ;
        RECT -238.875 -82.475 -238.705 -82.305 ;
        RECT -238.415 -82.475 -238.245 -82.305 ;
        RECT -237.955 -82.475 -237.785 -82.305 ;
        RECT -237.495 -82.475 -237.325 -82.305 ;
        RECT -237.035 -82.475 -236.865 -82.305 ;
        RECT -229.875 -82.475 -229.705 -82.305 ;
        RECT -229.415 -82.475 -229.245 -82.305 ;
        RECT -228.955 -82.475 -228.785 -82.305 ;
        RECT -228.495 -82.475 -228.325 -82.305 ;
        RECT -228.035 -82.475 -227.865 -82.305 ;
        RECT -227.575 -82.475 -227.405 -82.305 ;
        RECT -227.115 -82.475 -226.945 -82.305 ;
        RECT -219.955 -82.475 -219.785 -82.305 ;
        RECT -219.495 -82.475 -219.325 -82.305 ;
        RECT -219.035 -82.475 -218.865 -82.305 ;
        RECT -218.575 -82.475 -218.405 -82.305 ;
        RECT -218.115 -82.475 -217.945 -82.305 ;
        RECT -217.655 -82.475 -217.485 -82.305 ;
        RECT -217.195 -82.475 -217.025 -82.305 ;
        RECT -210.035 -82.475 -209.865 -82.305 ;
        RECT -209.575 -82.475 -209.405 -82.305 ;
        RECT -209.115 -82.475 -208.945 -82.305 ;
        RECT -208.655 -82.475 -208.485 -82.305 ;
        RECT -208.195 -82.475 -208.025 -82.305 ;
        RECT -207.735 -82.475 -207.565 -82.305 ;
        RECT -207.275 -82.475 -207.105 -82.305 ;
        RECT -200.115 -82.475 -199.945 -82.305 ;
        RECT -199.655 -82.475 -199.485 -82.305 ;
        RECT -199.195 -82.475 -199.025 -82.305 ;
        RECT -198.735 -82.475 -198.565 -82.305 ;
        RECT -198.275 -82.475 -198.105 -82.305 ;
        RECT -197.815 -82.475 -197.645 -82.305 ;
        RECT -197.355 -82.475 -197.185 -82.305 ;
        RECT -190.195 -82.475 -190.025 -82.305 ;
        RECT -189.735 -82.475 -189.565 -82.305 ;
        RECT -189.275 -82.475 -189.105 -82.305 ;
        RECT -188.815 -82.475 -188.645 -82.305 ;
        RECT -188.355 -82.475 -188.185 -82.305 ;
        RECT -187.895 -82.475 -187.725 -82.305 ;
        RECT -187.435 -82.475 -187.265 -82.305 ;
        RECT -180.275 -82.475 -180.105 -82.305 ;
        RECT -179.815 -82.475 -179.645 -82.305 ;
        RECT -179.355 -82.475 -179.185 -82.305 ;
        RECT -178.895 -82.475 -178.725 -82.305 ;
        RECT -178.435 -82.475 -178.265 -82.305 ;
        RECT -177.975 -82.475 -177.805 -82.305 ;
        RECT -177.515 -82.475 -177.345 -82.305 ;
        RECT -170.355 -82.475 -170.185 -82.305 ;
        RECT -169.895 -82.475 -169.725 -82.305 ;
        RECT -169.435 -82.475 -169.265 -82.305 ;
        RECT -168.975 -82.475 -168.805 -82.305 ;
        RECT -168.515 -82.475 -168.345 -82.305 ;
        RECT -168.055 -82.475 -167.885 -82.305 ;
        RECT -167.595 -82.475 -167.425 -82.305 ;
        RECT -160.435 -82.475 -160.265 -82.305 ;
        RECT -159.975 -82.475 -159.805 -82.305 ;
        RECT -159.515 -82.475 -159.345 -82.305 ;
        RECT -159.055 -82.475 -158.885 -82.305 ;
        RECT -158.595 -82.475 -158.425 -82.305 ;
        RECT -158.135 -82.475 -157.965 -82.305 ;
        RECT -157.675 -82.475 -157.505 -82.305 ;
        RECT -150.515 -82.475 -150.345 -82.305 ;
        RECT -150.055 -82.475 -149.885 -82.305 ;
        RECT -149.595 -82.475 -149.425 -82.305 ;
        RECT -149.135 -82.475 -148.965 -82.305 ;
        RECT -148.675 -82.475 -148.505 -82.305 ;
        RECT -148.215 -82.475 -148.045 -82.305 ;
        RECT -147.755 -82.475 -147.585 -82.305 ;
        RECT -140.595 -82.475 -140.425 -82.305 ;
        RECT -140.135 -82.475 -139.965 -82.305 ;
        RECT -139.675 -82.475 -139.505 -82.305 ;
        RECT -139.215 -82.475 -139.045 -82.305 ;
        RECT -138.755 -82.475 -138.585 -82.305 ;
        RECT -138.295 -82.475 -138.125 -82.305 ;
        RECT -137.835 -82.475 -137.665 -82.305 ;
        RECT -130.675 -82.475 -130.505 -82.305 ;
        RECT -130.215 -82.475 -130.045 -82.305 ;
        RECT -129.755 -82.475 -129.585 -82.305 ;
        RECT -129.295 -82.475 -129.125 -82.305 ;
        RECT -128.835 -82.475 -128.665 -82.305 ;
        RECT -128.375 -82.475 -128.205 -82.305 ;
        RECT -127.915 -82.475 -127.745 -82.305 ;
        RECT -120.755 -82.475 -120.585 -82.305 ;
        RECT -120.295 -82.475 -120.125 -82.305 ;
        RECT -119.835 -82.475 -119.665 -82.305 ;
        RECT -119.375 -82.475 -119.205 -82.305 ;
        RECT -118.915 -82.475 -118.745 -82.305 ;
        RECT -118.455 -82.475 -118.285 -82.305 ;
        RECT -117.995 -82.475 -117.825 -82.305 ;
        RECT -110.835 -82.475 -110.665 -82.305 ;
        RECT -110.375 -82.475 -110.205 -82.305 ;
        RECT -109.915 -82.475 -109.745 -82.305 ;
        RECT -109.455 -82.475 -109.285 -82.305 ;
        RECT -108.995 -82.475 -108.825 -82.305 ;
        RECT -108.535 -82.475 -108.365 -82.305 ;
        RECT -108.075 -82.475 -107.905 -82.305 ;
        RECT -100.915 -82.475 -100.745 -82.305 ;
        RECT -100.455 -82.475 -100.285 -82.305 ;
        RECT -99.995 -82.475 -99.825 -82.305 ;
        RECT -99.535 -82.475 -99.365 -82.305 ;
        RECT -99.075 -82.475 -98.905 -82.305 ;
        RECT -98.615 -82.475 -98.445 -82.305 ;
        RECT -98.155 -82.475 -97.985 -82.305 ;
        RECT -90.995 -82.475 -90.825 -82.305 ;
        RECT -90.535 -82.475 -90.365 -82.305 ;
        RECT -90.075 -82.475 -89.905 -82.305 ;
        RECT -89.615 -82.475 -89.445 -82.305 ;
        RECT -89.155 -82.475 -88.985 -82.305 ;
        RECT -88.695 -82.475 -88.525 -82.305 ;
        RECT -88.235 -82.475 -88.065 -82.305 ;
        RECT -81.075 -82.475 -80.905 -82.305 ;
        RECT -80.615 -82.475 -80.445 -82.305 ;
        RECT -80.155 -82.475 -79.985 -82.305 ;
        RECT -79.695 -82.475 -79.525 -82.305 ;
        RECT -79.235 -82.475 -79.065 -82.305 ;
        RECT -78.775 -82.475 -78.605 -82.305 ;
        RECT -78.315 -82.475 -78.145 -82.305 ;
        RECT -71.155 -82.475 -70.985 -82.305 ;
        RECT -70.695 -82.475 -70.525 -82.305 ;
        RECT -70.235 -82.475 -70.065 -82.305 ;
        RECT -69.775 -82.475 -69.605 -82.305 ;
        RECT -69.315 -82.475 -69.145 -82.305 ;
        RECT -68.855 -82.475 -68.685 -82.305 ;
        RECT -68.395 -82.475 -68.225 -82.305 ;
        RECT -61.235 -82.475 -61.065 -82.305 ;
        RECT -60.775 -82.475 -60.605 -82.305 ;
        RECT -60.315 -82.475 -60.145 -82.305 ;
        RECT -59.855 -82.475 -59.685 -82.305 ;
        RECT -59.395 -82.475 -59.225 -82.305 ;
        RECT -58.935 -82.475 -58.765 -82.305 ;
        RECT -58.475 -82.475 -58.305 -82.305 ;
        RECT -51.315 -82.475 -51.145 -82.305 ;
        RECT -50.855 -82.475 -50.685 -82.305 ;
        RECT -50.395 -82.475 -50.225 -82.305 ;
        RECT -49.935 -82.475 -49.765 -82.305 ;
        RECT -49.475 -82.475 -49.305 -82.305 ;
        RECT -49.015 -82.475 -48.845 -82.305 ;
        RECT -48.555 -82.475 -48.385 -82.305 ;
        RECT -41.395 -82.475 -41.225 -82.305 ;
        RECT -40.935 -82.475 -40.765 -82.305 ;
        RECT -40.475 -82.475 -40.305 -82.305 ;
        RECT -40.015 -82.475 -39.845 -82.305 ;
        RECT -39.555 -82.475 -39.385 -82.305 ;
        RECT -39.095 -82.475 -38.925 -82.305 ;
        RECT -38.635 -82.475 -38.465 -82.305 ;
        RECT -31.475 -82.475 -31.305 -82.305 ;
        RECT -31.015 -82.475 -30.845 -82.305 ;
        RECT -30.555 -82.475 -30.385 -82.305 ;
        RECT -30.095 -82.475 -29.925 -82.305 ;
        RECT -29.635 -82.475 -29.465 -82.305 ;
        RECT -29.175 -82.475 -29.005 -82.305 ;
        RECT -28.715 -82.475 -28.545 -82.305 ;
        RECT -21.555 -82.475 -21.385 -82.305 ;
        RECT -21.095 -82.475 -20.925 -82.305 ;
        RECT -20.635 -82.475 -20.465 -82.305 ;
        RECT -20.175 -82.475 -20.005 -82.305 ;
        RECT -19.715 -82.475 -19.545 -82.305 ;
        RECT -19.255 -82.475 -19.085 -82.305 ;
        RECT -18.795 -82.475 -18.625 -82.305 ;
        RECT -11.635 -82.475 -11.465 -82.305 ;
        RECT -11.175 -82.475 -11.005 -82.305 ;
        RECT -10.715 -82.475 -10.545 -82.305 ;
        RECT -10.255 -82.475 -10.085 -82.305 ;
        RECT -9.795 -82.475 -9.625 -82.305 ;
        RECT -9.335 -82.475 -9.165 -82.305 ;
        RECT -8.875 -82.475 -8.705 -82.305 ;
        RECT -1.715 -82.475 -1.545 -82.305 ;
        RECT -1.255 -82.475 -1.085 -82.305 ;
        RECT -0.795 -82.475 -0.625 -82.305 ;
        RECT -0.335 -82.475 -0.165 -82.305 ;
        RECT 0.125 -82.475 0.295 -82.305 ;
        RECT 0.585 -82.475 0.755 -82.305 ;
        RECT 1.045 -82.475 1.215 -82.305 ;
        RECT 8.205 -82.475 8.375 -82.305 ;
        RECT 8.665 -82.475 8.835 -82.305 ;
        RECT 9.125 -82.475 9.295 -82.305 ;
        RECT 9.585 -82.475 9.755 -82.305 ;
        RECT 10.045 -82.475 10.215 -82.305 ;
        RECT 10.505 -82.475 10.675 -82.305 ;
        RECT 10.965 -82.475 11.135 -82.305 ;
        RECT 18.125 -82.475 18.295 -82.305 ;
        RECT 18.585 -82.475 18.755 -82.305 ;
        RECT 19.045 -82.475 19.215 -82.305 ;
        RECT 19.505 -82.475 19.675 -82.305 ;
        RECT 19.965 -82.475 20.135 -82.305 ;
        RECT 20.425 -82.475 20.595 -82.305 ;
        RECT 20.885 -82.475 21.055 -82.305 ;
        RECT -284.825 -83.135 -284.655 -82.965 ;
        RECT -284.825 -83.595 -284.655 -83.425 ;
        RECT -281.285 -83.135 -281.115 -82.965 ;
        RECT -274.905 -83.135 -274.735 -82.965 ;
        RECT -281.285 -83.595 -281.115 -83.425 ;
        RECT -274.905 -83.595 -274.735 -83.425 ;
        RECT -283.055 -83.865 -282.885 -83.695 ;
        RECT -284.825 -84.055 -284.655 -83.885 ;
        RECT -281.285 -84.055 -281.115 -83.885 ;
        RECT -271.365 -83.135 -271.195 -82.965 ;
        RECT -264.985 -83.135 -264.815 -82.965 ;
        RECT -271.365 -83.595 -271.195 -83.425 ;
        RECT -264.985 -83.595 -264.815 -83.425 ;
        RECT -273.135 -83.865 -272.965 -83.695 ;
        RECT -274.905 -84.055 -274.735 -83.885 ;
        RECT -271.365 -84.055 -271.195 -83.885 ;
        RECT -261.445 -83.135 -261.275 -82.965 ;
        RECT -255.065 -83.135 -254.895 -82.965 ;
        RECT -261.445 -83.595 -261.275 -83.425 ;
        RECT -255.065 -83.595 -254.895 -83.425 ;
        RECT -263.215 -83.865 -263.045 -83.695 ;
        RECT -264.985 -84.055 -264.815 -83.885 ;
        RECT -261.445 -84.055 -261.275 -83.885 ;
        RECT -251.525 -83.135 -251.355 -82.965 ;
        RECT -245.145 -83.135 -244.975 -82.965 ;
        RECT -251.525 -83.595 -251.355 -83.425 ;
        RECT -245.145 -83.595 -244.975 -83.425 ;
        RECT -253.295 -83.865 -253.125 -83.695 ;
        RECT -255.065 -84.055 -254.895 -83.885 ;
        RECT -251.525 -84.055 -251.355 -83.885 ;
        RECT -241.605 -83.135 -241.435 -82.965 ;
        RECT -235.225 -83.135 -235.055 -82.965 ;
        RECT -241.605 -83.595 -241.435 -83.425 ;
        RECT -235.225 -83.595 -235.055 -83.425 ;
        RECT -243.375 -83.865 -243.205 -83.695 ;
        RECT -245.145 -84.055 -244.975 -83.885 ;
        RECT -241.605 -84.055 -241.435 -83.885 ;
        RECT -231.685 -83.135 -231.515 -82.965 ;
        RECT -225.305 -83.135 -225.135 -82.965 ;
        RECT -231.685 -83.595 -231.515 -83.425 ;
        RECT -225.305 -83.595 -225.135 -83.425 ;
        RECT -233.455 -83.865 -233.285 -83.695 ;
        RECT -235.225 -84.055 -235.055 -83.885 ;
        RECT -231.685 -84.055 -231.515 -83.885 ;
        RECT -221.765 -83.135 -221.595 -82.965 ;
        RECT -215.385 -83.135 -215.215 -82.965 ;
        RECT -221.765 -83.595 -221.595 -83.425 ;
        RECT -215.385 -83.595 -215.215 -83.425 ;
        RECT -223.535 -83.865 -223.365 -83.695 ;
        RECT -225.305 -84.055 -225.135 -83.885 ;
        RECT -221.765 -84.055 -221.595 -83.885 ;
        RECT -211.845 -83.135 -211.675 -82.965 ;
        RECT -205.465 -83.135 -205.295 -82.965 ;
        RECT -211.845 -83.595 -211.675 -83.425 ;
        RECT -205.465 -83.595 -205.295 -83.425 ;
        RECT -213.615 -83.865 -213.445 -83.695 ;
        RECT -215.385 -84.055 -215.215 -83.885 ;
        RECT -211.845 -84.055 -211.675 -83.885 ;
        RECT -201.925 -83.135 -201.755 -82.965 ;
        RECT -195.545 -83.135 -195.375 -82.965 ;
        RECT -201.925 -83.595 -201.755 -83.425 ;
        RECT -195.545 -83.595 -195.375 -83.425 ;
        RECT -203.695 -83.865 -203.525 -83.695 ;
        RECT -205.465 -84.055 -205.295 -83.885 ;
        RECT -201.925 -84.055 -201.755 -83.885 ;
        RECT -192.005 -83.135 -191.835 -82.965 ;
        RECT -185.625 -83.135 -185.455 -82.965 ;
        RECT -192.005 -83.595 -191.835 -83.425 ;
        RECT -185.625 -83.595 -185.455 -83.425 ;
        RECT -193.775 -83.865 -193.605 -83.695 ;
        RECT -195.545 -84.055 -195.375 -83.885 ;
        RECT -192.005 -84.055 -191.835 -83.885 ;
        RECT -182.085 -83.135 -181.915 -82.965 ;
        RECT -175.705 -83.135 -175.535 -82.965 ;
        RECT -182.085 -83.595 -181.915 -83.425 ;
        RECT -175.705 -83.595 -175.535 -83.425 ;
        RECT -183.855 -83.865 -183.685 -83.695 ;
        RECT -185.625 -84.055 -185.455 -83.885 ;
        RECT -182.085 -84.055 -181.915 -83.885 ;
        RECT -172.165 -83.135 -171.995 -82.965 ;
        RECT -165.785 -83.135 -165.615 -82.965 ;
        RECT -172.165 -83.595 -171.995 -83.425 ;
        RECT -165.785 -83.595 -165.615 -83.425 ;
        RECT -173.935 -83.865 -173.765 -83.695 ;
        RECT -175.705 -84.055 -175.535 -83.885 ;
        RECT -172.165 -84.055 -171.995 -83.885 ;
        RECT -162.245 -83.135 -162.075 -82.965 ;
        RECT -155.865 -83.135 -155.695 -82.965 ;
        RECT -162.245 -83.595 -162.075 -83.425 ;
        RECT -155.865 -83.595 -155.695 -83.425 ;
        RECT -164.015 -83.865 -163.845 -83.695 ;
        RECT -165.785 -84.055 -165.615 -83.885 ;
        RECT -162.245 -84.055 -162.075 -83.885 ;
        RECT -152.325 -83.135 -152.155 -82.965 ;
        RECT -145.945 -83.135 -145.775 -82.965 ;
        RECT -152.325 -83.595 -152.155 -83.425 ;
        RECT -145.945 -83.595 -145.775 -83.425 ;
        RECT -154.095 -83.865 -153.925 -83.695 ;
        RECT -155.865 -84.055 -155.695 -83.885 ;
        RECT -152.325 -84.055 -152.155 -83.885 ;
        RECT -142.405 -83.135 -142.235 -82.965 ;
        RECT -136.025 -83.135 -135.855 -82.965 ;
        RECT -142.405 -83.595 -142.235 -83.425 ;
        RECT -136.025 -83.595 -135.855 -83.425 ;
        RECT -144.175 -83.865 -144.005 -83.695 ;
        RECT -145.945 -84.055 -145.775 -83.885 ;
        RECT -142.405 -84.055 -142.235 -83.885 ;
        RECT -132.485 -83.135 -132.315 -82.965 ;
        RECT -126.105 -83.135 -125.935 -82.965 ;
        RECT -132.485 -83.595 -132.315 -83.425 ;
        RECT -126.105 -83.595 -125.935 -83.425 ;
        RECT -134.255 -83.865 -134.085 -83.695 ;
        RECT -136.025 -84.055 -135.855 -83.885 ;
        RECT -132.485 -84.055 -132.315 -83.885 ;
        RECT -122.565 -83.135 -122.395 -82.965 ;
        RECT -116.185 -83.135 -116.015 -82.965 ;
        RECT -122.565 -83.595 -122.395 -83.425 ;
        RECT -116.185 -83.595 -116.015 -83.425 ;
        RECT -124.335 -83.865 -124.165 -83.695 ;
        RECT -126.105 -84.055 -125.935 -83.885 ;
        RECT -122.565 -84.055 -122.395 -83.885 ;
        RECT -112.645 -83.135 -112.475 -82.965 ;
        RECT -106.265 -83.135 -106.095 -82.965 ;
        RECT -112.645 -83.595 -112.475 -83.425 ;
        RECT -106.265 -83.595 -106.095 -83.425 ;
        RECT -114.415 -83.865 -114.245 -83.695 ;
        RECT -116.185 -84.055 -116.015 -83.885 ;
        RECT -112.645 -84.055 -112.475 -83.885 ;
        RECT -102.725 -83.135 -102.555 -82.965 ;
        RECT -96.345 -83.135 -96.175 -82.965 ;
        RECT -102.725 -83.595 -102.555 -83.425 ;
        RECT -96.345 -83.595 -96.175 -83.425 ;
        RECT -104.495 -83.865 -104.325 -83.695 ;
        RECT -106.265 -84.055 -106.095 -83.885 ;
        RECT -102.725 -84.055 -102.555 -83.885 ;
        RECT -92.805 -83.135 -92.635 -82.965 ;
        RECT -86.425 -83.135 -86.255 -82.965 ;
        RECT -92.805 -83.595 -92.635 -83.425 ;
        RECT -86.425 -83.595 -86.255 -83.425 ;
        RECT -94.575 -83.865 -94.405 -83.695 ;
        RECT -96.345 -84.055 -96.175 -83.885 ;
        RECT -92.805 -84.055 -92.635 -83.885 ;
        RECT -82.885 -83.135 -82.715 -82.965 ;
        RECT -76.505 -83.135 -76.335 -82.965 ;
        RECT -82.885 -83.595 -82.715 -83.425 ;
        RECT -76.505 -83.595 -76.335 -83.425 ;
        RECT -84.655 -83.865 -84.485 -83.695 ;
        RECT -86.425 -84.055 -86.255 -83.885 ;
        RECT -82.885 -84.055 -82.715 -83.885 ;
        RECT -72.965 -83.135 -72.795 -82.965 ;
        RECT -66.585 -83.135 -66.415 -82.965 ;
        RECT -72.965 -83.595 -72.795 -83.425 ;
        RECT -66.585 -83.595 -66.415 -83.425 ;
        RECT -74.735 -83.865 -74.565 -83.695 ;
        RECT -76.505 -84.055 -76.335 -83.885 ;
        RECT -72.965 -84.055 -72.795 -83.885 ;
        RECT -63.045 -83.135 -62.875 -82.965 ;
        RECT -56.665 -83.135 -56.495 -82.965 ;
        RECT -63.045 -83.595 -62.875 -83.425 ;
        RECT -56.665 -83.595 -56.495 -83.425 ;
        RECT -64.815 -83.865 -64.645 -83.695 ;
        RECT -66.585 -84.055 -66.415 -83.885 ;
        RECT -63.045 -84.055 -62.875 -83.885 ;
        RECT -53.125 -83.135 -52.955 -82.965 ;
        RECT -46.745 -83.135 -46.575 -82.965 ;
        RECT -53.125 -83.595 -52.955 -83.425 ;
        RECT -46.745 -83.595 -46.575 -83.425 ;
        RECT -54.895 -83.865 -54.725 -83.695 ;
        RECT -56.665 -84.055 -56.495 -83.885 ;
        RECT -53.125 -84.055 -52.955 -83.885 ;
        RECT -43.205 -83.135 -43.035 -82.965 ;
        RECT -36.825 -83.135 -36.655 -82.965 ;
        RECT -43.205 -83.595 -43.035 -83.425 ;
        RECT -36.825 -83.595 -36.655 -83.425 ;
        RECT -44.975 -83.865 -44.805 -83.695 ;
        RECT -46.745 -84.055 -46.575 -83.885 ;
        RECT -43.205 -84.055 -43.035 -83.885 ;
        RECT -33.285 -83.135 -33.115 -82.965 ;
        RECT -26.905 -83.135 -26.735 -82.965 ;
        RECT -33.285 -83.595 -33.115 -83.425 ;
        RECT -26.905 -83.595 -26.735 -83.425 ;
        RECT -35.055 -83.865 -34.885 -83.695 ;
        RECT -36.825 -84.055 -36.655 -83.885 ;
        RECT -33.285 -84.055 -33.115 -83.885 ;
        RECT -23.365 -83.135 -23.195 -82.965 ;
        RECT -16.985 -83.135 -16.815 -82.965 ;
        RECT -23.365 -83.595 -23.195 -83.425 ;
        RECT -16.985 -83.595 -16.815 -83.425 ;
        RECT -25.135 -83.865 -24.965 -83.695 ;
        RECT -26.905 -84.055 -26.735 -83.885 ;
        RECT -23.365 -84.055 -23.195 -83.885 ;
        RECT -13.445 -83.135 -13.275 -82.965 ;
        RECT -7.065 -83.135 -6.895 -82.965 ;
        RECT -13.445 -83.595 -13.275 -83.425 ;
        RECT -7.065 -83.595 -6.895 -83.425 ;
        RECT -15.215 -83.865 -15.045 -83.695 ;
        RECT -16.985 -84.055 -16.815 -83.885 ;
        RECT -13.445 -84.055 -13.275 -83.885 ;
        RECT -3.525 -83.135 -3.355 -82.965 ;
        RECT 2.855 -83.135 3.025 -82.965 ;
        RECT -3.525 -83.595 -3.355 -83.425 ;
        RECT 2.855 -83.595 3.025 -83.425 ;
        RECT -5.295 -83.865 -5.125 -83.695 ;
        RECT -7.065 -84.055 -6.895 -83.885 ;
        RECT -3.525 -84.055 -3.355 -83.885 ;
        RECT 6.395 -83.135 6.565 -82.965 ;
        RECT 12.775 -83.135 12.945 -82.965 ;
        RECT 6.395 -83.595 6.565 -83.425 ;
        RECT 12.775 -83.595 12.945 -83.425 ;
        RECT 4.625 -83.865 4.795 -83.695 ;
        RECT 2.855 -84.055 3.025 -83.885 ;
        RECT 6.395 -84.055 6.565 -83.885 ;
        RECT 16.315 -83.135 16.485 -82.965 ;
        RECT 16.315 -83.595 16.485 -83.425 ;
        RECT 14.545 -83.865 14.715 -83.695 ;
        RECT 12.775 -84.055 12.945 -83.885 ;
        RECT 16.315 -84.055 16.485 -83.885 ;
        RECT -291.545 -172.755 -291.375 -172.585 ;
        RECT -289.775 -172.855 -289.605 -172.685 ;
        RECT -288.005 -172.755 -287.835 -172.585 ;
        RECT -291.545 -173.215 -291.375 -173.045 ;
        RECT -291.545 -173.675 -291.375 -173.505 ;
        RECT -281.625 -172.755 -281.455 -172.585 ;
        RECT -279.855 -172.855 -279.685 -172.685 ;
        RECT -278.085 -172.755 -277.915 -172.585 ;
        RECT -288.005 -173.215 -287.835 -173.045 ;
        RECT -281.625 -173.215 -281.455 -173.045 ;
        RECT -288.005 -173.675 -287.835 -173.505 ;
        RECT -281.625 -173.675 -281.455 -173.505 ;
        RECT -271.705 -172.755 -271.535 -172.585 ;
        RECT -269.935 -172.855 -269.765 -172.685 ;
        RECT -268.165 -172.755 -267.995 -172.585 ;
        RECT -278.085 -173.215 -277.915 -173.045 ;
        RECT -271.705 -173.215 -271.535 -173.045 ;
        RECT -278.085 -173.675 -277.915 -173.505 ;
        RECT -271.705 -173.675 -271.535 -173.505 ;
        RECT -261.785 -172.755 -261.615 -172.585 ;
        RECT -260.015 -172.855 -259.845 -172.685 ;
        RECT -258.245 -172.755 -258.075 -172.585 ;
        RECT -268.165 -173.215 -267.995 -173.045 ;
        RECT -261.785 -173.215 -261.615 -173.045 ;
        RECT -268.165 -173.675 -267.995 -173.505 ;
        RECT -261.785 -173.675 -261.615 -173.505 ;
        RECT -251.865 -172.755 -251.695 -172.585 ;
        RECT -250.095 -172.855 -249.925 -172.685 ;
        RECT -248.325 -172.755 -248.155 -172.585 ;
        RECT -258.245 -173.215 -258.075 -173.045 ;
        RECT -251.865 -173.215 -251.695 -173.045 ;
        RECT -258.245 -173.675 -258.075 -173.505 ;
        RECT -251.865 -173.675 -251.695 -173.505 ;
        RECT -241.945 -172.755 -241.775 -172.585 ;
        RECT -240.175 -172.855 -240.005 -172.685 ;
        RECT -238.405 -172.755 -238.235 -172.585 ;
        RECT -248.325 -173.215 -248.155 -173.045 ;
        RECT -241.945 -173.215 -241.775 -173.045 ;
        RECT -248.325 -173.675 -248.155 -173.505 ;
        RECT -241.945 -173.675 -241.775 -173.505 ;
        RECT -232.025 -172.755 -231.855 -172.585 ;
        RECT -230.255 -172.855 -230.085 -172.685 ;
        RECT -228.485 -172.755 -228.315 -172.585 ;
        RECT -238.405 -173.215 -238.235 -173.045 ;
        RECT -232.025 -173.215 -231.855 -173.045 ;
        RECT -238.405 -173.675 -238.235 -173.505 ;
        RECT -232.025 -173.675 -231.855 -173.505 ;
        RECT -222.105 -172.755 -221.935 -172.585 ;
        RECT -220.335 -172.855 -220.165 -172.685 ;
        RECT -218.565 -172.755 -218.395 -172.585 ;
        RECT -228.485 -173.215 -228.315 -173.045 ;
        RECT -222.105 -173.215 -221.935 -173.045 ;
        RECT -228.485 -173.675 -228.315 -173.505 ;
        RECT -222.105 -173.675 -221.935 -173.505 ;
        RECT -212.185 -172.755 -212.015 -172.585 ;
        RECT -210.415 -172.855 -210.245 -172.685 ;
        RECT -208.645 -172.755 -208.475 -172.585 ;
        RECT -218.565 -173.215 -218.395 -173.045 ;
        RECT -212.185 -173.215 -212.015 -173.045 ;
        RECT -218.565 -173.675 -218.395 -173.505 ;
        RECT -212.185 -173.675 -212.015 -173.505 ;
        RECT -202.265 -172.755 -202.095 -172.585 ;
        RECT -200.495 -172.855 -200.325 -172.685 ;
        RECT -198.725 -172.755 -198.555 -172.585 ;
        RECT -208.645 -173.215 -208.475 -173.045 ;
        RECT -202.265 -173.215 -202.095 -173.045 ;
        RECT -208.645 -173.675 -208.475 -173.505 ;
        RECT -202.265 -173.675 -202.095 -173.505 ;
        RECT -192.345 -172.755 -192.175 -172.585 ;
        RECT -190.575 -172.855 -190.405 -172.685 ;
        RECT -188.805 -172.755 -188.635 -172.585 ;
        RECT -198.725 -173.215 -198.555 -173.045 ;
        RECT -192.345 -173.215 -192.175 -173.045 ;
        RECT -198.725 -173.675 -198.555 -173.505 ;
        RECT -192.345 -173.675 -192.175 -173.505 ;
        RECT -182.425 -172.755 -182.255 -172.585 ;
        RECT -180.655 -172.855 -180.485 -172.685 ;
        RECT -178.885 -172.755 -178.715 -172.585 ;
        RECT -188.805 -173.215 -188.635 -173.045 ;
        RECT -182.425 -173.215 -182.255 -173.045 ;
        RECT -188.805 -173.675 -188.635 -173.505 ;
        RECT -182.425 -173.675 -182.255 -173.505 ;
        RECT -172.505 -172.755 -172.335 -172.585 ;
        RECT -170.735 -172.855 -170.565 -172.685 ;
        RECT -168.965 -172.755 -168.795 -172.585 ;
        RECT -178.885 -173.215 -178.715 -173.045 ;
        RECT -172.505 -173.215 -172.335 -173.045 ;
        RECT -178.885 -173.675 -178.715 -173.505 ;
        RECT -172.505 -173.675 -172.335 -173.505 ;
        RECT -162.585 -172.755 -162.415 -172.585 ;
        RECT -160.815 -172.855 -160.645 -172.685 ;
        RECT -159.045 -172.755 -158.875 -172.585 ;
        RECT -168.965 -173.215 -168.795 -173.045 ;
        RECT -162.585 -173.215 -162.415 -173.045 ;
        RECT -168.965 -173.675 -168.795 -173.505 ;
        RECT -162.585 -173.675 -162.415 -173.505 ;
        RECT -152.665 -172.755 -152.495 -172.585 ;
        RECT -150.895 -172.855 -150.725 -172.685 ;
        RECT -149.125 -172.755 -148.955 -172.585 ;
        RECT -159.045 -173.215 -158.875 -173.045 ;
        RECT -152.665 -173.215 -152.495 -173.045 ;
        RECT -159.045 -173.675 -158.875 -173.505 ;
        RECT -152.665 -173.675 -152.495 -173.505 ;
        RECT -142.745 -172.755 -142.575 -172.585 ;
        RECT -140.975 -172.855 -140.805 -172.685 ;
        RECT -139.205 -172.755 -139.035 -172.585 ;
        RECT -149.125 -173.215 -148.955 -173.045 ;
        RECT -142.745 -173.215 -142.575 -173.045 ;
        RECT -149.125 -173.675 -148.955 -173.505 ;
        RECT -142.745 -173.675 -142.575 -173.505 ;
        RECT -132.825 -172.755 -132.655 -172.585 ;
        RECT -131.055 -172.855 -130.885 -172.685 ;
        RECT -129.285 -172.755 -129.115 -172.585 ;
        RECT -139.205 -173.215 -139.035 -173.045 ;
        RECT -132.825 -173.215 -132.655 -173.045 ;
        RECT -139.205 -173.675 -139.035 -173.505 ;
        RECT -132.825 -173.675 -132.655 -173.505 ;
        RECT -122.905 -172.755 -122.735 -172.585 ;
        RECT -121.135 -172.855 -120.965 -172.685 ;
        RECT -119.365 -172.755 -119.195 -172.585 ;
        RECT -129.285 -173.215 -129.115 -173.045 ;
        RECT -122.905 -173.215 -122.735 -173.045 ;
        RECT -129.285 -173.675 -129.115 -173.505 ;
        RECT -122.905 -173.675 -122.735 -173.505 ;
        RECT -112.985 -172.755 -112.815 -172.585 ;
        RECT -111.215 -172.855 -111.045 -172.685 ;
        RECT -109.445 -172.755 -109.275 -172.585 ;
        RECT -119.365 -173.215 -119.195 -173.045 ;
        RECT -112.985 -173.215 -112.815 -173.045 ;
        RECT -119.365 -173.675 -119.195 -173.505 ;
        RECT -112.985 -173.675 -112.815 -173.505 ;
        RECT -103.065 -172.755 -102.895 -172.585 ;
        RECT -101.295 -172.855 -101.125 -172.685 ;
        RECT -99.525 -172.755 -99.355 -172.585 ;
        RECT -109.445 -173.215 -109.275 -173.045 ;
        RECT -103.065 -173.215 -102.895 -173.045 ;
        RECT -109.445 -173.675 -109.275 -173.505 ;
        RECT -103.065 -173.675 -102.895 -173.505 ;
        RECT -93.145 -172.755 -92.975 -172.585 ;
        RECT -91.375 -172.855 -91.205 -172.685 ;
        RECT -89.605 -172.755 -89.435 -172.585 ;
        RECT -99.525 -173.215 -99.355 -173.045 ;
        RECT -93.145 -173.215 -92.975 -173.045 ;
        RECT -99.525 -173.675 -99.355 -173.505 ;
        RECT -93.145 -173.675 -92.975 -173.505 ;
        RECT -83.225 -172.755 -83.055 -172.585 ;
        RECT -81.455 -172.855 -81.285 -172.685 ;
        RECT -79.685 -172.755 -79.515 -172.585 ;
        RECT -89.605 -173.215 -89.435 -173.045 ;
        RECT -83.225 -173.215 -83.055 -173.045 ;
        RECT -89.605 -173.675 -89.435 -173.505 ;
        RECT -83.225 -173.675 -83.055 -173.505 ;
        RECT -73.305 -172.755 -73.135 -172.585 ;
        RECT -71.535 -172.855 -71.365 -172.685 ;
        RECT -69.765 -172.755 -69.595 -172.585 ;
        RECT -79.685 -173.215 -79.515 -173.045 ;
        RECT -73.305 -173.215 -73.135 -173.045 ;
        RECT -79.685 -173.675 -79.515 -173.505 ;
        RECT -73.305 -173.675 -73.135 -173.505 ;
        RECT -63.385 -172.755 -63.215 -172.585 ;
        RECT -61.615 -172.855 -61.445 -172.685 ;
        RECT -59.845 -172.755 -59.675 -172.585 ;
        RECT -69.765 -173.215 -69.595 -173.045 ;
        RECT -63.385 -173.215 -63.215 -173.045 ;
        RECT -69.765 -173.675 -69.595 -173.505 ;
        RECT -63.385 -173.675 -63.215 -173.505 ;
        RECT -53.465 -172.755 -53.295 -172.585 ;
        RECT -51.695 -172.855 -51.525 -172.685 ;
        RECT -49.925 -172.755 -49.755 -172.585 ;
        RECT -59.845 -173.215 -59.675 -173.045 ;
        RECT -53.465 -173.215 -53.295 -173.045 ;
        RECT -59.845 -173.675 -59.675 -173.505 ;
        RECT -53.465 -173.675 -53.295 -173.505 ;
        RECT -43.545 -172.755 -43.375 -172.585 ;
        RECT -41.775 -172.855 -41.605 -172.685 ;
        RECT -40.005 -172.755 -39.835 -172.585 ;
        RECT -49.925 -173.215 -49.755 -173.045 ;
        RECT -43.545 -173.215 -43.375 -173.045 ;
        RECT -49.925 -173.675 -49.755 -173.505 ;
        RECT -43.545 -173.675 -43.375 -173.505 ;
        RECT -33.625 -172.755 -33.455 -172.585 ;
        RECT -31.855 -172.855 -31.685 -172.685 ;
        RECT -30.085 -172.755 -29.915 -172.585 ;
        RECT -40.005 -173.215 -39.835 -173.045 ;
        RECT -33.625 -173.215 -33.455 -173.045 ;
        RECT -40.005 -173.675 -39.835 -173.505 ;
        RECT -33.625 -173.675 -33.455 -173.505 ;
        RECT -23.705 -172.755 -23.535 -172.585 ;
        RECT -21.935 -172.855 -21.765 -172.685 ;
        RECT -20.165 -172.755 -19.995 -172.585 ;
        RECT -30.085 -173.215 -29.915 -173.045 ;
        RECT -23.705 -173.215 -23.535 -173.045 ;
        RECT -30.085 -173.675 -29.915 -173.505 ;
        RECT -23.705 -173.675 -23.535 -173.505 ;
        RECT -13.785 -172.755 -13.615 -172.585 ;
        RECT -12.015 -172.855 -11.845 -172.685 ;
        RECT -10.245 -172.755 -10.075 -172.585 ;
        RECT -20.165 -173.215 -19.995 -173.045 ;
        RECT -13.785 -173.215 -13.615 -173.045 ;
        RECT -20.165 -173.675 -19.995 -173.505 ;
        RECT -13.785 -173.675 -13.615 -173.505 ;
        RECT -3.865 -172.755 -3.695 -172.585 ;
        RECT -2.095 -172.855 -1.925 -172.685 ;
        RECT -0.325 -172.755 -0.155 -172.585 ;
        RECT -10.245 -173.215 -10.075 -173.045 ;
        RECT -3.865 -173.215 -3.695 -173.045 ;
        RECT -10.245 -173.675 -10.075 -173.505 ;
        RECT -3.865 -173.675 -3.695 -173.505 ;
        RECT 6.055 -172.755 6.225 -172.585 ;
        RECT 7.825 -172.855 7.995 -172.685 ;
        RECT 9.595 -172.755 9.765 -172.585 ;
        RECT -0.325 -173.215 -0.155 -173.045 ;
        RECT 6.055 -173.215 6.225 -173.045 ;
        RECT -0.325 -173.675 -0.155 -173.505 ;
        RECT 6.055 -173.675 6.225 -173.505 ;
        RECT 15.975 -172.755 16.145 -172.585 ;
        RECT 17.745 -172.855 17.915 -172.685 ;
        RECT 19.515 -172.755 19.685 -172.585 ;
        RECT 9.595 -173.215 9.765 -173.045 ;
        RECT 15.975 -173.215 16.145 -173.045 ;
        RECT 9.595 -173.675 9.765 -173.505 ;
        RECT 15.975 -173.675 16.145 -173.505 ;
        RECT 19.515 -173.215 19.685 -173.045 ;
        RECT 19.515 -173.675 19.685 -173.505 ;
        RECT -286.195 -174.335 -286.025 -174.165 ;
        RECT -285.735 -174.335 -285.565 -174.165 ;
        RECT -285.275 -174.335 -285.105 -174.165 ;
        RECT -284.815 -174.335 -284.645 -174.165 ;
        RECT -284.355 -174.335 -284.185 -174.165 ;
        RECT -283.895 -174.335 -283.725 -174.165 ;
        RECT -283.435 -174.335 -283.265 -174.165 ;
        RECT -276.275 -174.335 -276.105 -174.165 ;
        RECT -275.815 -174.335 -275.645 -174.165 ;
        RECT -275.355 -174.335 -275.185 -174.165 ;
        RECT -274.895 -174.335 -274.725 -174.165 ;
        RECT -274.435 -174.335 -274.265 -174.165 ;
        RECT -273.975 -174.335 -273.805 -174.165 ;
        RECT -273.515 -174.335 -273.345 -174.165 ;
        RECT -266.355 -174.335 -266.185 -174.165 ;
        RECT -265.895 -174.335 -265.725 -174.165 ;
        RECT -265.435 -174.335 -265.265 -174.165 ;
        RECT -264.975 -174.335 -264.805 -174.165 ;
        RECT -264.515 -174.335 -264.345 -174.165 ;
        RECT -264.055 -174.335 -263.885 -174.165 ;
        RECT -263.595 -174.335 -263.425 -174.165 ;
        RECT -256.435 -174.335 -256.265 -174.165 ;
        RECT -255.975 -174.335 -255.805 -174.165 ;
        RECT -255.515 -174.335 -255.345 -174.165 ;
        RECT -255.055 -174.335 -254.885 -174.165 ;
        RECT -254.595 -174.335 -254.425 -174.165 ;
        RECT -254.135 -174.335 -253.965 -174.165 ;
        RECT -253.675 -174.335 -253.505 -174.165 ;
        RECT -246.515 -174.335 -246.345 -174.165 ;
        RECT -246.055 -174.335 -245.885 -174.165 ;
        RECT -245.595 -174.335 -245.425 -174.165 ;
        RECT -245.135 -174.335 -244.965 -174.165 ;
        RECT -244.675 -174.335 -244.505 -174.165 ;
        RECT -244.215 -174.335 -244.045 -174.165 ;
        RECT -243.755 -174.335 -243.585 -174.165 ;
        RECT -236.595 -174.335 -236.425 -174.165 ;
        RECT -236.135 -174.335 -235.965 -174.165 ;
        RECT -235.675 -174.335 -235.505 -174.165 ;
        RECT -235.215 -174.335 -235.045 -174.165 ;
        RECT -234.755 -174.335 -234.585 -174.165 ;
        RECT -234.295 -174.335 -234.125 -174.165 ;
        RECT -233.835 -174.335 -233.665 -174.165 ;
        RECT -226.675 -174.335 -226.505 -174.165 ;
        RECT -226.215 -174.335 -226.045 -174.165 ;
        RECT -225.755 -174.335 -225.585 -174.165 ;
        RECT -225.295 -174.335 -225.125 -174.165 ;
        RECT -224.835 -174.335 -224.665 -174.165 ;
        RECT -224.375 -174.335 -224.205 -174.165 ;
        RECT -223.915 -174.335 -223.745 -174.165 ;
        RECT -216.755 -174.335 -216.585 -174.165 ;
        RECT -216.295 -174.335 -216.125 -174.165 ;
        RECT -215.835 -174.335 -215.665 -174.165 ;
        RECT -215.375 -174.335 -215.205 -174.165 ;
        RECT -214.915 -174.335 -214.745 -174.165 ;
        RECT -214.455 -174.335 -214.285 -174.165 ;
        RECT -213.995 -174.335 -213.825 -174.165 ;
        RECT -206.835 -174.335 -206.665 -174.165 ;
        RECT -206.375 -174.335 -206.205 -174.165 ;
        RECT -205.915 -174.335 -205.745 -174.165 ;
        RECT -205.455 -174.335 -205.285 -174.165 ;
        RECT -204.995 -174.335 -204.825 -174.165 ;
        RECT -204.535 -174.335 -204.365 -174.165 ;
        RECT -204.075 -174.335 -203.905 -174.165 ;
        RECT -196.915 -174.335 -196.745 -174.165 ;
        RECT -196.455 -174.335 -196.285 -174.165 ;
        RECT -195.995 -174.335 -195.825 -174.165 ;
        RECT -195.535 -174.335 -195.365 -174.165 ;
        RECT -195.075 -174.335 -194.905 -174.165 ;
        RECT -194.615 -174.335 -194.445 -174.165 ;
        RECT -194.155 -174.335 -193.985 -174.165 ;
        RECT -186.995 -174.335 -186.825 -174.165 ;
        RECT -186.535 -174.335 -186.365 -174.165 ;
        RECT -186.075 -174.335 -185.905 -174.165 ;
        RECT -185.615 -174.335 -185.445 -174.165 ;
        RECT -185.155 -174.335 -184.985 -174.165 ;
        RECT -184.695 -174.335 -184.525 -174.165 ;
        RECT -184.235 -174.335 -184.065 -174.165 ;
        RECT -177.075 -174.335 -176.905 -174.165 ;
        RECT -176.615 -174.335 -176.445 -174.165 ;
        RECT -176.155 -174.335 -175.985 -174.165 ;
        RECT -175.695 -174.335 -175.525 -174.165 ;
        RECT -175.235 -174.335 -175.065 -174.165 ;
        RECT -174.775 -174.335 -174.605 -174.165 ;
        RECT -174.315 -174.335 -174.145 -174.165 ;
        RECT -167.155 -174.335 -166.985 -174.165 ;
        RECT -166.695 -174.335 -166.525 -174.165 ;
        RECT -166.235 -174.335 -166.065 -174.165 ;
        RECT -165.775 -174.335 -165.605 -174.165 ;
        RECT -165.315 -174.335 -165.145 -174.165 ;
        RECT -164.855 -174.335 -164.685 -174.165 ;
        RECT -164.395 -174.335 -164.225 -174.165 ;
        RECT -157.235 -174.335 -157.065 -174.165 ;
        RECT -156.775 -174.335 -156.605 -174.165 ;
        RECT -156.315 -174.335 -156.145 -174.165 ;
        RECT -155.855 -174.335 -155.685 -174.165 ;
        RECT -155.395 -174.335 -155.225 -174.165 ;
        RECT -154.935 -174.335 -154.765 -174.165 ;
        RECT -154.475 -174.335 -154.305 -174.165 ;
        RECT -147.315 -174.335 -147.145 -174.165 ;
        RECT -146.855 -174.335 -146.685 -174.165 ;
        RECT -146.395 -174.335 -146.225 -174.165 ;
        RECT -145.935 -174.335 -145.765 -174.165 ;
        RECT -145.475 -174.335 -145.305 -174.165 ;
        RECT -145.015 -174.335 -144.845 -174.165 ;
        RECT -144.555 -174.335 -144.385 -174.165 ;
        RECT -137.395 -174.335 -137.225 -174.165 ;
        RECT -136.935 -174.335 -136.765 -174.165 ;
        RECT -136.475 -174.335 -136.305 -174.165 ;
        RECT -136.015 -174.335 -135.845 -174.165 ;
        RECT -135.555 -174.335 -135.385 -174.165 ;
        RECT -135.095 -174.335 -134.925 -174.165 ;
        RECT -134.635 -174.335 -134.465 -174.165 ;
        RECT -127.475 -174.335 -127.305 -174.165 ;
        RECT -127.015 -174.335 -126.845 -174.165 ;
        RECT -126.555 -174.335 -126.385 -174.165 ;
        RECT -126.095 -174.335 -125.925 -174.165 ;
        RECT -125.635 -174.335 -125.465 -174.165 ;
        RECT -125.175 -174.335 -125.005 -174.165 ;
        RECT -124.715 -174.335 -124.545 -174.165 ;
        RECT -117.555 -174.335 -117.385 -174.165 ;
        RECT -117.095 -174.335 -116.925 -174.165 ;
        RECT -116.635 -174.335 -116.465 -174.165 ;
        RECT -116.175 -174.335 -116.005 -174.165 ;
        RECT -115.715 -174.335 -115.545 -174.165 ;
        RECT -115.255 -174.335 -115.085 -174.165 ;
        RECT -114.795 -174.335 -114.625 -174.165 ;
        RECT -107.635 -174.335 -107.465 -174.165 ;
        RECT -107.175 -174.335 -107.005 -174.165 ;
        RECT -106.715 -174.335 -106.545 -174.165 ;
        RECT -106.255 -174.335 -106.085 -174.165 ;
        RECT -105.795 -174.335 -105.625 -174.165 ;
        RECT -105.335 -174.335 -105.165 -174.165 ;
        RECT -104.875 -174.335 -104.705 -174.165 ;
        RECT -97.715 -174.335 -97.545 -174.165 ;
        RECT -97.255 -174.335 -97.085 -174.165 ;
        RECT -96.795 -174.335 -96.625 -174.165 ;
        RECT -96.335 -174.335 -96.165 -174.165 ;
        RECT -95.875 -174.335 -95.705 -174.165 ;
        RECT -95.415 -174.335 -95.245 -174.165 ;
        RECT -94.955 -174.335 -94.785 -174.165 ;
        RECT -87.795 -174.335 -87.625 -174.165 ;
        RECT -87.335 -174.335 -87.165 -174.165 ;
        RECT -86.875 -174.335 -86.705 -174.165 ;
        RECT -86.415 -174.335 -86.245 -174.165 ;
        RECT -85.955 -174.335 -85.785 -174.165 ;
        RECT -85.495 -174.335 -85.325 -174.165 ;
        RECT -85.035 -174.335 -84.865 -174.165 ;
        RECT -77.875 -174.335 -77.705 -174.165 ;
        RECT -77.415 -174.335 -77.245 -174.165 ;
        RECT -76.955 -174.335 -76.785 -174.165 ;
        RECT -76.495 -174.335 -76.325 -174.165 ;
        RECT -76.035 -174.335 -75.865 -174.165 ;
        RECT -75.575 -174.335 -75.405 -174.165 ;
        RECT -75.115 -174.335 -74.945 -174.165 ;
        RECT -67.955 -174.335 -67.785 -174.165 ;
        RECT -67.495 -174.335 -67.325 -174.165 ;
        RECT -67.035 -174.335 -66.865 -174.165 ;
        RECT -66.575 -174.335 -66.405 -174.165 ;
        RECT -66.115 -174.335 -65.945 -174.165 ;
        RECT -65.655 -174.335 -65.485 -174.165 ;
        RECT -65.195 -174.335 -65.025 -174.165 ;
        RECT -58.035 -174.335 -57.865 -174.165 ;
        RECT -57.575 -174.335 -57.405 -174.165 ;
        RECT -57.115 -174.335 -56.945 -174.165 ;
        RECT -56.655 -174.335 -56.485 -174.165 ;
        RECT -56.195 -174.335 -56.025 -174.165 ;
        RECT -55.735 -174.335 -55.565 -174.165 ;
        RECT -55.275 -174.335 -55.105 -174.165 ;
        RECT -48.115 -174.335 -47.945 -174.165 ;
        RECT -47.655 -174.335 -47.485 -174.165 ;
        RECT -47.195 -174.335 -47.025 -174.165 ;
        RECT -46.735 -174.335 -46.565 -174.165 ;
        RECT -46.275 -174.335 -46.105 -174.165 ;
        RECT -45.815 -174.335 -45.645 -174.165 ;
        RECT -45.355 -174.335 -45.185 -174.165 ;
        RECT -38.195 -174.335 -38.025 -174.165 ;
        RECT -37.735 -174.335 -37.565 -174.165 ;
        RECT -37.275 -174.335 -37.105 -174.165 ;
        RECT -36.815 -174.335 -36.645 -174.165 ;
        RECT -36.355 -174.335 -36.185 -174.165 ;
        RECT -35.895 -174.335 -35.725 -174.165 ;
        RECT -35.435 -174.335 -35.265 -174.165 ;
        RECT -28.275 -174.335 -28.105 -174.165 ;
        RECT -27.815 -174.335 -27.645 -174.165 ;
        RECT -27.355 -174.335 -27.185 -174.165 ;
        RECT -26.895 -174.335 -26.725 -174.165 ;
        RECT -26.435 -174.335 -26.265 -174.165 ;
        RECT -25.975 -174.335 -25.805 -174.165 ;
        RECT -25.515 -174.335 -25.345 -174.165 ;
        RECT -18.355 -174.335 -18.185 -174.165 ;
        RECT -17.895 -174.335 -17.725 -174.165 ;
        RECT -17.435 -174.335 -17.265 -174.165 ;
        RECT -16.975 -174.335 -16.805 -174.165 ;
        RECT -16.515 -174.335 -16.345 -174.165 ;
        RECT -16.055 -174.335 -15.885 -174.165 ;
        RECT -15.595 -174.335 -15.425 -174.165 ;
        RECT -8.435 -174.335 -8.265 -174.165 ;
        RECT -7.975 -174.335 -7.805 -174.165 ;
        RECT -7.515 -174.335 -7.345 -174.165 ;
        RECT -7.055 -174.335 -6.885 -174.165 ;
        RECT -6.595 -174.335 -6.425 -174.165 ;
        RECT -6.135 -174.335 -5.965 -174.165 ;
        RECT -5.675 -174.335 -5.505 -174.165 ;
        RECT 1.485 -174.335 1.655 -174.165 ;
        RECT 1.945 -174.335 2.115 -174.165 ;
        RECT 2.405 -174.335 2.575 -174.165 ;
        RECT 2.865 -174.335 3.035 -174.165 ;
        RECT 3.325 -174.335 3.495 -174.165 ;
        RECT 3.785 -174.335 3.955 -174.165 ;
        RECT 4.245 -174.335 4.415 -174.165 ;
        RECT 11.405 -174.335 11.575 -174.165 ;
        RECT 11.865 -174.335 12.035 -174.165 ;
        RECT 12.325 -174.335 12.495 -174.165 ;
        RECT 12.785 -174.335 12.955 -174.165 ;
        RECT 13.245 -174.335 13.415 -174.165 ;
        RECT 13.705 -174.335 13.875 -174.165 ;
        RECT 14.165 -174.335 14.335 -174.165 ;
        RECT -291.155 -177.055 -290.985 -176.885 ;
        RECT -290.695 -177.055 -290.525 -176.885 ;
        RECT -290.235 -177.055 -290.065 -176.885 ;
        RECT -289.775 -177.055 -289.605 -176.885 ;
        RECT -289.315 -177.055 -289.145 -176.885 ;
        RECT -288.855 -177.055 -288.685 -176.885 ;
        RECT -288.395 -177.055 -288.225 -176.885 ;
        RECT -281.235 -177.055 -281.065 -176.885 ;
        RECT -280.775 -177.055 -280.605 -176.885 ;
        RECT -280.315 -177.055 -280.145 -176.885 ;
        RECT -279.855 -177.055 -279.685 -176.885 ;
        RECT -279.395 -177.055 -279.225 -176.885 ;
        RECT -278.935 -177.055 -278.765 -176.885 ;
        RECT -278.475 -177.055 -278.305 -176.885 ;
        RECT -271.315 -177.055 -271.145 -176.885 ;
        RECT -270.855 -177.055 -270.685 -176.885 ;
        RECT -270.395 -177.055 -270.225 -176.885 ;
        RECT -269.935 -177.055 -269.765 -176.885 ;
        RECT -269.475 -177.055 -269.305 -176.885 ;
        RECT -269.015 -177.055 -268.845 -176.885 ;
        RECT -268.555 -177.055 -268.385 -176.885 ;
        RECT -261.395 -177.055 -261.225 -176.885 ;
        RECT -260.935 -177.055 -260.765 -176.885 ;
        RECT -260.475 -177.055 -260.305 -176.885 ;
        RECT -260.015 -177.055 -259.845 -176.885 ;
        RECT -259.555 -177.055 -259.385 -176.885 ;
        RECT -259.095 -177.055 -258.925 -176.885 ;
        RECT -258.635 -177.055 -258.465 -176.885 ;
        RECT -251.475 -177.055 -251.305 -176.885 ;
        RECT -251.015 -177.055 -250.845 -176.885 ;
        RECT -250.555 -177.055 -250.385 -176.885 ;
        RECT -250.095 -177.055 -249.925 -176.885 ;
        RECT -249.635 -177.055 -249.465 -176.885 ;
        RECT -249.175 -177.055 -249.005 -176.885 ;
        RECT -248.715 -177.055 -248.545 -176.885 ;
        RECT -241.555 -177.055 -241.385 -176.885 ;
        RECT -241.095 -177.055 -240.925 -176.885 ;
        RECT -240.635 -177.055 -240.465 -176.885 ;
        RECT -240.175 -177.055 -240.005 -176.885 ;
        RECT -239.715 -177.055 -239.545 -176.885 ;
        RECT -239.255 -177.055 -239.085 -176.885 ;
        RECT -238.795 -177.055 -238.625 -176.885 ;
        RECT -231.635 -177.055 -231.465 -176.885 ;
        RECT -231.175 -177.055 -231.005 -176.885 ;
        RECT -230.715 -177.055 -230.545 -176.885 ;
        RECT -230.255 -177.055 -230.085 -176.885 ;
        RECT -229.795 -177.055 -229.625 -176.885 ;
        RECT -229.335 -177.055 -229.165 -176.885 ;
        RECT -228.875 -177.055 -228.705 -176.885 ;
        RECT -221.715 -177.055 -221.545 -176.885 ;
        RECT -221.255 -177.055 -221.085 -176.885 ;
        RECT -220.795 -177.055 -220.625 -176.885 ;
        RECT -220.335 -177.055 -220.165 -176.885 ;
        RECT -219.875 -177.055 -219.705 -176.885 ;
        RECT -219.415 -177.055 -219.245 -176.885 ;
        RECT -218.955 -177.055 -218.785 -176.885 ;
        RECT -211.795 -177.055 -211.625 -176.885 ;
        RECT -211.335 -177.055 -211.165 -176.885 ;
        RECT -210.875 -177.055 -210.705 -176.885 ;
        RECT -210.415 -177.055 -210.245 -176.885 ;
        RECT -209.955 -177.055 -209.785 -176.885 ;
        RECT -209.495 -177.055 -209.325 -176.885 ;
        RECT -209.035 -177.055 -208.865 -176.885 ;
        RECT -201.875 -177.055 -201.705 -176.885 ;
        RECT -201.415 -177.055 -201.245 -176.885 ;
        RECT -200.955 -177.055 -200.785 -176.885 ;
        RECT -200.495 -177.055 -200.325 -176.885 ;
        RECT -200.035 -177.055 -199.865 -176.885 ;
        RECT -199.575 -177.055 -199.405 -176.885 ;
        RECT -199.115 -177.055 -198.945 -176.885 ;
        RECT -191.955 -177.055 -191.785 -176.885 ;
        RECT -191.495 -177.055 -191.325 -176.885 ;
        RECT -191.035 -177.055 -190.865 -176.885 ;
        RECT -190.575 -177.055 -190.405 -176.885 ;
        RECT -190.115 -177.055 -189.945 -176.885 ;
        RECT -189.655 -177.055 -189.485 -176.885 ;
        RECT -189.195 -177.055 -189.025 -176.885 ;
        RECT -182.035 -177.055 -181.865 -176.885 ;
        RECT -181.575 -177.055 -181.405 -176.885 ;
        RECT -181.115 -177.055 -180.945 -176.885 ;
        RECT -180.655 -177.055 -180.485 -176.885 ;
        RECT -180.195 -177.055 -180.025 -176.885 ;
        RECT -179.735 -177.055 -179.565 -176.885 ;
        RECT -179.275 -177.055 -179.105 -176.885 ;
        RECT -172.115 -177.055 -171.945 -176.885 ;
        RECT -171.655 -177.055 -171.485 -176.885 ;
        RECT -171.195 -177.055 -171.025 -176.885 ;
        RECT -170.735 -177.055 -170.565 -176.885 ;
        RECT -170.275 -177.055 -170.105 -176.885 ;
        RECT -169.815 -177.055 -169.645 -176.885 ;
        RECT -169.355 -177.055 -169.185 -176.885 ;
        RECT -162.195 -177.055 -162.025 -176.885 ;
        RECT -161.735 -177.055 -161.565 -176.885 ;
        RECT -161.275 -177.055 -161.105 -176.885 ;
        RECT -160.815 -177.055 -160.645 -176.885 ;
        RECT -160.355 -177.055 -160.185 -176.885 ;
        RECT -159.895 -177.055 -159.725 -176.885 ;
        RECT -159.435 -177.055 -159.265 -176.885 ;
        RECT -152.275 -177.055 -152.105 -176.885 ;
        RECT -151.815 -177.055 -151.645 -176.885 ;
        RECT -151.355 -177.055 -151.185 -176.885 ;
        RECT -150.895 -177.055 -150.725 -176.885 ;
        RECT -150.435 -177.055 -150.265 -176.885 ;
        RECT -149.975 -177.055 -149.805 -176.885 ;
        RECT -149.515 -177.055 -149.345 -176.885 ;
        RECT -142.355 -177.055 -142.185 -176.885 ;
        RECT -141.895 -177.055 -141.725 -176.885 ;
        RECT -141.435 -177.055 -141.265 -176.885 ;
        RECT -140.975 -177.055 -140.805 -176.885 ;
        RECT -140.515 -177.055 -140.345 -176.885 ;
        RECT -140.055 -177.055 -139.885 -176.885 ;
        RECT -139.595 -177.055 -139.425 -176.885 ;
        RECT -132.435 -177.055 -132.265 -176.885 ;
        RECT -131.975 -177.055 -131.805 -176.885 ;
        RECT -131.515 -177.055 -131.345 -176.885 ;
        RECT -131.055 -177.055 -130.885 -176.885 ;
        RECT -130.595 -177.055 -130.425 -176.885 ;
        RECT -130.135 -177.055 -129.965 -176.885 ;
        RECT -129.675 -177.055 -129.505 -176.885 ;
        RECT -122.515 -177.055 -122.345 -176.885 ;
        RECT -122.055 -177.055 -121.885 -176.885 ;
        RECT -121.595 -177.055 -121.425 -176.885 ;
        RECT -121.135 -177.055 -120.965 -176.885 ;
        RECT -120.675 -177.055 -120.505 -176.885 ;
        RECT -120.215 -177.055 -120.045 -176.885 ;
        RECT -119.755 -177.055 -119.585 -176.885 ;
        RECT -112.595 -177.055 -112.425 -176.885 ;
        RECT -112.135 -177.055 -111.965 -176.885 ;
        RECT -111.675 -177.055 -111.505 -176.885 ;
        RECT -111.215 -177.055 -111.045 -176.885 ;
        RECT -110.755 -177.055 -110.585 -176.885 ;
        RECT -110.295 -177.055 -110.125 -176.885 ;
        RECT -109.835 -177.055 -109.665 -176.885 ;
        RECT -102.675 -177.055 -102.505 -176.885 ;
        RECT -102.215 -177.055 -102.045 -176.885 ;
        RECT -101.755 -177.055 -101.585 -176.885 ;
        RECT -101.295 -177.055 -101.125 -176.885 ;
        RECT -100.835 -177.055 -100.665 -176.885 ;
        RECT -100.375 -177.055 -100.205 -176.885 ;
        RECT -99.915 -177.055 -99.745 -176.885 ;
        RECT -92.755 -177.055 -92.585 -176.885 ;
        RECT -92.295 -177.055 -92.125 -176.885 ;
        RECT -91.835 -177.055 -91.665 -176.885 ;
        RECT -91.375 -177.055 -91.205 -176.885 ;
        RECT -90.915 -177.055 -90.745 -176.885 ;
        RECT -90.455 -177.055 -90.285 -176.885 ;
        RECT -89.995 -177.055 -89.825 -176.885 ;
        RECT -82.835 -177.055 -82.665 -176.885 ;
        RECT -82.375 -177.055 -82.205 -176.885 ;
        RECT -81.915 -177.055 -81.745 -176.885 ;
        RECT -81.455 -177.055 -81.285 -176.885 ;
        RECT -80.995 -177.055 -80.825 -176.885 ;
        RECT -80.535 -177.055 -80.365 -176.885 ;
        RECT -80.075 -177.055 -79.905 -176.885 ;
        RECT -72.915 -177.055 -72.745 -176.885 ;
        RECT -72.455 -177.055 -72.285 -176.885 ;
        RECT -71.995 -177.055 -71.825 -176.885 ;
        RECT -71.535 -177.055 -71.365 -176.885 ;
        RECT -71.075 -177.055 -70.905 -176.885 ;
        RECT -70.615 -177.055 -70.445 -176.885 ;
        RECT -70.155 -177.055 -69.985 -176.885 ;
        RECT -62.995 -177.055 -62.825 -176.885 ;
        RECT -62.535 -177.055 -62.365 -176.885 ;
        RECT -62.075 -177.055 -61.905 -176.885 ;
        RECT -61.615 -177.055 -61.445 -176.885 ;
        RECT -61.155 -177.055 -60.985 -176.885 ;
        RECT -60.695 -177.055 -60.525 -176.885 ;
        RECT -60.235 -177.055 -60.065 -176.885 ;
        RECT -53.075 -177.055 -52.905 -176.885 ;
        RECT -52.615 -177.055 -52.445 -176.885 ;
        RECT -52.155 -177.055 -51.985 -176.885 ;
        RECT -51.695 -177.055 -51.525 -176.885 ;
        RECT -51.235 -177.055 -51.065 -176.885 ;
        RECT -50.775 -177.055 -50.605 -176.885 ;
        RECT -50.315 -177.055 -50.145 -176.885 ;
        RECT -43.155 -177.055 -42.985 -176.885 ;
        RECT -42.695 -177.055 -42.525 -176.885 ;
        RECT -42.235 -177.055 -42.065 -176.885 ;
        RECT -41.775 -177.055 -41.605 -176.885 ;
        RECT -41.315 -177.055 -41.145 -176.885 ;
        RECT -40.855 -177.055 -40.685 -176.885 ;
        RECT -40.395 -177.055 -40.225 -176.885 ;
        RECT -33.235 -177.055 -33.065 -176.885 ;
        RECT -32.775 -177.055 -32.605 -176.885 ;
        RECT -32.315 -177.055 -32.145 -176.885 ;
        RECT -31.855 -177.055 -31.685 -176.885 ;
        RECT -31.395 -177.055 -31.225 -176.885 ;
        RECT -30.935 -177.055 -30.765 -176.885 ;
        RECT -30.475 -177.055 -30.305 -176.885 ;
        RECT -23.315 -177.055 -23.145 -176.885 ;
        RECT -22.855 -177.055 -22.685 -176.885 ;
        RECT -22.395 -177.055 -22.225 -176.885 ;
        RECT -21.935 -177.055 -21.765 -176.885 ;
        RECT -21.475 -177.055 -21.305 -176.885 ;
        RECT -21.015 -177.055 -20.845 -176.885 ;
        RECT -20.555 -177.055 -20.385 -176.885 ;
        RECT -13.395 -177.055 -13.225 -176.885 ;
        RECT -12.935 -177.055 -12.765 -176.885 ;
        RECT -12.475 -177.055 -12.305 -176.885 ;
        RECT -12.015 -177.055 -11.845 -176.885 ;
        RECT -11.555 -177.055 -11.385 -176.885 ;
        RECT -11.095 -177.055 -10.925 -176.885 ;
        RECT -10.635 -177.055 -10.465 -176.885 ;
        RECT -3.475 -177.055 -3.305 -176.885 ;
        RECT -3.015 -177.055 -2.845 -176.885 ;
        RECT -2.555 -177.055 -2.385 -176.885 ;
        RECT -2.095 -177.055 -1.925 -176.885 ;
        RECT -1.635 -177.055 -1.465 -176.885 ;
        RECT -1.175 -177.055 -1.005 -176.885 ;
        RECT -0.715 -177.055 -0.545 -176.885 ;
        RECT 6.445 -177.055 6.615 -176.885 ;
        RECT 6.905 -177.055 7.075 -176.885 ;
        RECT 7.365 -177.055 7.535 -176.885 ;
        RECT 7.825 -177.055 7.995 -176.885 ;
        RECT 8.285 -177.055 8.455 -176.885 ;
        RECT 8.745 -177.055 8.915 -176.885 ;
        RECT 9.205 -177.055 9.375 -176.885 ;
        RECT 16.365 -177.055 16.535 -176.885 ;
        RECT 16.825 -177.055 16.995 -176.885 ;
        RECT 17.285 -177.055 17.455 -176.885 ;
        RECT 17.745 -177.055 17.915 -176.885 ;
        RECT 18.205 -177.055 18.375 -176.885 ;
        RECT 18.665 -177.055 18.835 -176.885 ;
        RECT 19.125 -177.055 19.295 -176.885 ;
        RECT -286.585 -177.715 -286.415 -177.545 ;
        RECT -286.585 -178.175 -286.415 -178.005 ;
        RECT -283.045 -177.715 -282.875 -177.545 ;
        RECT -276.665 -177.715 -276.495 -177.545 ;
        RECT -283.045 -178.175 -282.875 -178.005 ;
        RECT -276.665 -178.175 -276.495 -178.005 ;
        RECT -284.815 -178.445 -284.645 -178.275 ;
        RECT -286.585 -178.635 -286.415 -178.465 ;
        RECT -283.045 -178.635 -282.875 -178.465 ;
        RECT -273.125 -177.715 -272.955 -177.545 ;
        RECT -266.745 -177.715 -266.575 -177.545 ;
        RECT -273.125 -178.175 -272.955 -178.005 ;
        RECT -266.745 -178.175 -266.575 -178.005 ;
        RECT -274.895 -178.445 -274.725 -178.275 ;
        RECT -276.665 -178.635 -276.495 -178.465 ;
        RECT -273.125 -178.635 -272.955 -178.465 ;
        RECT -263.205 -177.715 -263.035 -177.545 ;
        RECT -256.825 -177.715 -256.655 -177.545 ;
        RECT -263.205 -178.175 -263.035 -178.005 ;
        RECT -256.825 -178.175 -256.655 -178.005 ;
        RECT -264.975 -178.445 -264.805 -178.275 ;
        RECT -266.745 -178.635 -266.575 -178.465 ;
        RECT -263.205 -178.635 -263.035 -178.465 ;
        RECT -253.285 -177.715 -253.115 -177.545 ;
        RECT -246.905 -177.715 -246.735 -177.545 ;
        RECT -253.285 -178.175 -253.115 -178.005 ;
        RECT -246.905 -178.175 -246.735 -178.005 ;
        RECT -255.055 -178.445 -254.885 -178.275 ;
        RECT -256.825 -178.635 -256.655 -178.465 ;
        RECT -253.285 -178.635 -253.115 -178.465 ;
        RECT -243.365 -177.715 -243.195 -177.545 ;
        RECT -236.985 -177.715 -236.815 -177.545 ;
        RECT -243.365 -178.175 -243.195 -178.005 ;
        RECT -236.985 -178.175 -236.815 -178.005 ;
        RECT -245.135 -178.445 -244.965 -178.275 ;
        RECT -246.905 -178.635 -246.735 -178.465 ;
        RECT -243.365 -178.635 -243.195 -178.465 ;
        RECT -233.445 -177.715 -233.275 -177.545 ;
        RECT -227.065 -177.715 -226.895 -177.545 ;
        RECT -233.445 -178.175 -233.275 -178.005 ;
        RECT -227.065 -178.175 -226.895 -178.005 ;
        RECT -235.215 -178.445 -235.045 -178.275 ;
        RECT -236.985 -178.635 -236.815 -178.465 ;
        RECT -233.445 -178.635 -233.275 -178.465 ;
        RECT -223.525 -177.715 -223.355 -177.545 ;
        RECT -217.145 -177.715 -216.975 -177.545 ;
        RECT -223.525 -178.175 -223.355 -178.005 ;
        RECT -217.145 -178.175 -216.975 -178.005 ;
        RECT -225.295 -178.445 -225.125 -178.275 ;
        RECT -227.065 -178.635 -226.895 -178.465 ;
        RECT -223.525 -178.635 -223.355 -178.465 ;
        RECT -213.605 -177.715 -213.435 -177.545 ;
        RECT -207.225 -177.715 -207.055 -177.545 ;
        RECT -213.605 -178.175 -213.435 -178.005 ;
        RECT -207.225 -178.175 -207.055 -178.005 ;
        RECT -215.375 -178.445 -215.205 -178.275 ;
        RECT -217.145 -178.635 -216.975 -178.465 ;
        RECT -213.605 -178.635 -213.435 -178.465 ;
        RECT -203.685 -177.715 -203.515 -177.545 ;
        RECT -197.305 -177.715 -197.135 -177.545 ;
        RECT -203.685 -178.175 -203.515 -178.005 ;
        RECT -197.305 -178.175 -197.135 -178.005 ;
        RECT -205.455 -178.445 -205.285 -178.275 ;
        RECT -207.225 -178.635 -207.055 -178.465 ;
        RECT -203.685 -178.635 -203.515 -178.465 ;
        RECT -193.765 -177.715 -193.595 -177.545 ;
        RECT -187.385 -177.715 -187.215 -177.545 ;
        RECT -193.765 -178.175 -193.595 -178.005 ;
        RECT -187.385 -178.175 -187.215 -178.005 ;
        RECT -195.535 -178.445 -195.365 -178.275 ;
        RECT -197.305 -178.635 -197.135 -178.465 ;
        RECT -193.765 -178.635 -193.595 -178.465 ;
        RECT -183.845 -177.715 -183.675 -177.545 ;
        RECT -177.465 -177.715 -177.295 -177.545 ;
        RECT -183.845 -178.175 -183.675 -178.005 ;
        RECT -177.465 -178.175 -177.295 -178.005 ;
        RECT -185.615 -178.445 -185.445 -178.275 ;
        RECT -187.385 -178.635 -187.215 -178.465 ;
        RECT -183.845 -178.635 -183.675 -178.465 ;
        RECT -173.925 -177.715 -173.755 -177.545 ;
        RECT -167.545 -177.715 -167.375 -177.545 ;
        RECT -173.925 -178.175 -173.755 -178.005 ;
        RECT -167.545 -178.175 -167.375 -178.005 ;
        RECT -175.695 -178.445 -175.525 -178.275 ;
        RECT -177.465 -178.635 -177.295 -178.465 ;
        RECT -173.925 -178.635 -173.755 -178.465 ;
        RECT -164.005 -177.715 -163.835 -177.545 ;
        RECT -157.625 -177.715 -157.455 -177.545 ;
        RECT -164.005 -178.175 -163.835 -178.005 ;
        RECT -157.625 -178.175 -157.455 -178.005 ;
        RECT -165.775 -178.445 -165.605 -178.275 ;
        RECT -167.545 -178.635 -167.375 -178.465 ;
        RECT -164.005 -178.635 -163.835 -178.465 ;
        RECT -154.085 -177.715 -153.915 -177.545 ;
        RECT -147.705 -177.715 -147.535 -177.545 ;
        RECT -154.085 -178.175 -153.915 -178.005 ;
        RECT -147.705 -178.175 -147.535 -178.005 ;
        RECT -155.855 -178.445 -155.685 -178.275 ;
        RECT -157.625 -178.635 -157.455 -178.465 ;
        RECT -154.085 -178.635 -153.915 -178.465 ;
        RECT -144.165 -177.715 -143.995 -177.545 ;
        RECT -137.785 -177.715 -137.615 -177.545 ;
        RECT -144.165 -178.175 -143.995 -178.005 ;
        RECT -137.785 -178.175 -137.615 -178.005 ;
        RECT -145.935 -178.445 -145.765 -178.275 ;
        RECT -147.705 -178.635 -147.535 -178.465 ;
        RECT -144.165 -178.635 -143.995 -178.465 ;
        RECT -134.245 -177.715 -134.075 -177.545 ;
        RECT -127.865 -177.715 -127.695 -177.545 ;
        RECT -134.245 -178.175 -134.075 -178.005 ;
        RECT -127.865 -178.175 -127.695 -178.005 ;
        RECT -136.015 -178.445 -135.845 -178.275 ;
        RECT -137.785 -178.635 -137.615 -178.465 ;
        RECT -134.245 -178.635 -134.075 -178.465 ;
        RECT -124.325 -177.715 -124.155 -177.545 ;
        RECT -117.945 -177.715 -117.775 -177.545 ;
        RECT -124.325 -178.175 -124.155 -178.005 ;
        RECT -117.945 -178.175 -117.775 -178.005 ;
        RECT -126.095 -178.445 -125.925 -178.275 ;
        RECT -127.865 -178.635 -127.695 -178.465 ;
        RECT -124.325 -178.635 -124.155 -178.465 ;
        RECT -114.405 -177.715 -114.235 -177.545 ;
        RECT -108.025 -177.715 -107.855 -177.545 ;
        RECT -114.405 -178.175 -114.235 -178.005 ;
        RECT -108.025 -178.175 -107.855 -178.005 ;
        RECT -116.175 -178.445 -116.005 -178.275 ;
        RECT -117.945 -178.635 -117.775 -178.465 ;
        RECT -114.405 -178.635 -114.235 -178.465 ;
        RECT -104.485 -177.715 -104.315 -177.545 ;
        RECT -98.105 -177.715 -97.935 -177.545 ;
        RECT -104.485 -178.175 -104.315 -178.005 ;
        RECT -98.105 -178.175 -97.935 -178.005 ;
        RECT -106.255 -178.445 -106.085 -178.275 ;
        RECT -108.025 -178.635 -107.855 -178.465 ;
        RECT -104.485 -178.635 -104.315 -178.465 ;
        RECT -94.565 -177.715 -94.395 -177.545 ;
        RECT -88.185 -177.715 -88.015 -177.545 ;
        RECT -94.565 -178.175 -94.395 -178.005 ;
        RECT -88.185 -178.175 -88.015 -178.005 ;
        RECT -96.335 -178.445 -96.165 -178.275 ;
        RECT -98.105 -178.635 -97.935 -178.465 ;
        RECT -94.565 -178.635 -94.395 -178.465 ;
        RECT -84.645 -177.715 -84.475 -177.545 ;
        RECT -78.265 -177.715 -78.095 -177.545 ;
        RECT -84.645 -178.175 -84.475 -178.005 ;
        RECT -78.265 -178.175 -78.095 -178.005 ;
        RECT -86.415 -178.445 -86.245 -178.275 ;
        RECT -88.185 -178.635 -88.015 -178.465 ;
        RECT -84.645 -178.635 -84.475 -178.465 ;
        RECT -74.725 -177.715 -74.555 -177.545 ;
        RECT -68.345 -177.715 -68.175 -177.545 ;
        RECT -74.725 -178.175 -74.555 -178.005 ;
        RECT -68.345 -178.175 -68.175 -178.005 ;
        RECT -76.495 -178.445 -76.325 -178.275 ;
        RECT -78.265 -178.635 -78.095 -178.465 ;
        RECT -74.725 -178.635 -74.555 -178.465 ;
        RECT -64.805 -177.715 -64.635 -177.545 ;
        RECT -58.425 -177.715 -58.255 -177.545 ;
        RECT -64.805 -178.175 -64.635 -178.005 ;
        RECT -58.425 -178.175 -58.255 -178.005 ;
        RECT -66.575 -178.445 -66.405 -178.275 ;
        RECT -68.345 -178.635 -68.175 -178.465 ;
        RECT -64.805 -178.635 -64.635 -178.465 ;
        RECT -54.885 -177.715 -54.715 -177.545 ;
        RECT -48.505 -177.715 -48.335 -177.545 ;
        RECT -54.885 -178.175 -54.715 -178.005 ;
        RECT -48.505 -178.175 -48.335 -178.005 ;
        RECT -56.655 -178.445 -56.485 -178.275 ;
        RECT -58.425 -178.635 -58.255 -178.465 ;
        RECT -54.885 -178.635 -54.715 -178.465 ;
        RECT -44.965 -177.715 -44.795 -177.545 ;
        RECT -38.585 -177.715 -38.415 -177.545 ;
        RECT -44.965 -178.175 -44.795 -178.005 ;
        RECT -38.585 -178.175 -38.415 -178.005 ;
        RECT -46.735 -178.445 -46.565 -178.275 ;
        RECT -48.505 -178.635 -48.335 -178.465 ;
        RECT -44.965 -178.635 -44.795 -178.465 ;
        RECT -35.045 -177.715 -34.875 -177.545 ;
        RECT -28.665 -177.715 -28.495 -177.545 ;
        RECT -35.045 -178.175 -34.875 -178.005 ;
        RECT -28.665 -178.175 -28.495 -178.005 ;
        RECT -36.815 -178.445 -36.645 -178.275 ;
        RECT -38.585 -178.635 -38.415 -178.465 ;
        RECT -35.045 -178.635 -34.875 -178.465 ;
        RECT -25.125 -177.715 -24.955 -177.545 ;
        RECT -18.745 -177.715 -18.575 -177.545 ;
        RECT -25.125 -178.175 -24.955 -178.005 ;
        RECT -18.745 -178.175 -18.575 -178.005 ;
        RECT -26.895 -178.445 -26.725 -178.275 ;
        RECT -28.665 -178.635 -28.495 -178.465 ;
        RECT -25.125 -178.635 -24.955 -178.465 ;
        RECT -15.205 -177.715 -15.035 -177.545 ;
        RECT -8.825 -177.715 -8.655 -177.545 ;
        RECT -15.205 -178.175 -15.035 -178.005 ;
        RECT -8.825 -178.175 -8.655 -178.005 ;
        RECT -16.975 -178.445 -16.805 -178.275 ;
        RECT -18.745 -178.635 -18.575 -178.465 ;
        RECT -15.205 -178.635 -15.035 -178.465 ;
        RECT -5.285 -177.715 -5.115 -177.545 ;
        RECT 1.095 -177.715 1.265 -177.545 ;
        RECT -5.285 -178.175 -5.115 -178.005 ;
        RECT 1.095 -178.175 1.265 -178.005 ;
        RECT -7.055 -178.445 -6.885 -178.275 ;
        RECT -8.825 -178.635 -8.655 -178.465 ;
        RECT -5.285 -178.635 -5.115 -178.465 ;
        RECT 4.635 -177.715 4.805 -177.545 ;
        RECT 11.015 -177.715 11.185 -177.545 ;
        RECT 4.635 -178.175 4.805 -178.005 ;
        RECT 11.015 -178.175 11.185 -178.005 ;
        RECT 2.865 -178.445 3.035 -178.275 ;
        RECT 1.095 -178.635 1.265 -178.465 ;
        RECT 4.635 -178.635 4.805 -178.465 ;
        RECT 14.555 -177.715 14.725 -177.545 ;
        RECT 14.555 -178.175 14.725 -178.005 ;
        RECT 12.785 -178.445 12.955 -178.275 ;
        RECT 11.015 -178.635 11.185 -178.465 ;
        RECT 14.555 -178.635 14.725 -178.465 ;
      LAYER met1 ;
        RECT -288.280 93.760 -284.260 95.140 ;
        RECT -278.360 93.760 -274.340 95.140 ;
        RECT -268.440 93.760 -264.420 95.140 ;
        RECT -258.520 93.760 -254.500 95.140 ;
        RECT -248.600 93.760 -244.580 95.140 ;
        RECT -238.680 93.760 -234.660 95.140 ;
        RECT -228.760 93.760 -224.740 95.140 ;
        RECT -218.840 93.760 -214.820 95.140 ;
        RECT -208.920 93.760 -204.900 95.140 ;
        RECT -199.000 93.760 -194.980 95.140 ;
        RECT -189.080 93.760 -185.060 95.140 ;
        RECT -179.160 93.760 -175.140 95.140 ;
        RECT -169.240 93.760 -165.220 95.140 ;
        RECT -159.320 93.760 -155.300 95.140 ;
        RECT -149.400 93.760 -145.380 95.140 ;
        RECT -139.480 93.760 -135.460 95.140 ;
        RECT -129.560 93.760 -125.540 95.140 ;
        RECT -119.640 93.760 -115.620 95.140 ;
        RECT -109.720 93.760 -105.700 95.140 ;
        RECT -99.800 93.760 -95.780 95.140 ;
        RECT -89.880 93.760 -85.860 95.140 ;
        RECT -79.960 93.760 -75.940 95.140 ;
        RECT -70.040 93.760 -66.020 95.140 ;
        RECT -60.120 93.760 -56.100 95.140 ;
        RECT -50.200 93.760 -46.180 95.140 ;
        RECT -40.280 93.760 -36.260 95.140 ;
        RECT -30.360 93.760 -26.340 95.140 ;
        RECT -20.440 93.760 -16.420 95.140 ;
        RECT -10.520 93.760 -6.500 95.140 ;
        RECT -0.600 93.760 3.420 95.140 ;
        RECT 9.320 93.760 13.340 95.140 ;
        RECT 19.240 93.760 23.260 95.140 ;
        RECT -282.920 93.090 -279.700 93.570 ;
        RECT -273.000 93.090 -269.780 93.570 ;
        RECT -263.080 93.090 -259.860 93.570 ;
        RECT -253.160 93.090 -249.940 93.570 ;
        RECT -243.240 93.090 -240.020 93.570 ;
        RECT -233.320 93.090 -230.100 93.570 ;
        RECT -223.400 93.090 -220.180 93.570 ;
        RECT -213.480 93.090 -210.260 93.570 ;
        RECT -203.560 93.090 -200.340 93.570 ;
        RECT -193.640 93.090 -190.420 93.570 ;
        RECT -183.720 93.090 -180.500 93.570 ;
        RECT -173.800 93.090 -170.580 93.570 ;
        RECT -163.880 93.090 -160.660 93.570 ;
        RECT -153.960 93.090 -150.740 93.570 ;
        RECT -144.040 93.090 -140.820 93.570 ;
        RECT -134.120 93.090 -130.900 93.570 ;
        RECT -124.200 93.090 -120.980 93.570 ;
        RECT -114.280 93.090 -111.060 93.570 ;
        RECT -104.360 93.090 -101.140 93.570 ;
        RECT -94.440 93.090 -91.220 93.570 ;
        RECT -84.520 93.090 -81.300 93.570 ;
        RECT -74.600 93.090 -71.380 93.570 ;
        RECT -64.680 93.090 -61.460 93.570 ;
        RECT -54.760 93.090 -51.540 93.570 ;
        RECT -44.840 93.090 -41.620 93.570 ;
        RECT -34.920 93.090 -31.700 93.570 ;
        RECT -25.000 93.090 -21.780 93.570 ;
        RECT -15.080 93.090 -11.860 93.570 ;
        RECT -5.160 93.090 -1.940 93.570 ;
        RECT 4.760 93.090 7.980 93.570 ;
        RECT 14.680 93.090 17.900 93.570 ;
        RECT -287.880 90.370 -284.660 90.850 ;
        RECT -277.960 90.370 -274.740 90.850 ;
        RECT -268.040 90.370 -264.820 90.850 ;
        RECT -258.120 90.370 -254.900 90.850 ;
        RECT -248.200 90.370 -244.980 90.850 ;
        RECT -238.280 90.370 -235.060 90.850 ;
        RECT -228.360 90.370 -225.140 90.850 ;
        RECT -218.440 90.370 -215.220 90.850 ;
        RECT -208.520 90.370 -205.300 90.850 ;
        RECT -198.600 90.370 -195.380 90.850 ;
        RECT -188.680 90.370 -185.460 90.850 ;
        RECT -178.760 90.370 -175.540 90.850 ;
        RECT -168.840 90.370 -165.620 90.850 ;
        RECT -158.920 90.370 -155.700 90.850 ;
        RECT -149.000 90.370 -145.780 90.850 ;
        RECT -139.080 90.370 -135.860 90.850 ;
        RECT -129.160 90.370 -125.940 90.850 ;
        RECT -119.240 90.370 -116.020 90.850 ;
        RECT -109.320 90.370 -106.100 90.850 ;
        RECT -99.400 90.370 -96.180 90.850 ;
        RECT -89.480 90.370 -86.260 90.850 ;
        RECT -79.560 90.370 -76.340 90.850 ;
        RECT -69.640 90.370 -66.420 90.850 ;
        RECT -59.720 90.370 -56.500 90.850 ;
        RECT -49.800 90.370 -46.580 90.850 ;
        RECT -39.880 90.370 -36.660 90.850 ;
        RECT -29.960 90.370 -26.740 90.850 ;
        RECT -20.040 90.370 -16.820 90.850 ;
        RECT -10.120 90.370 -6.900 90.850 ;
        RECT -0.200 90.370 3.020 90.850 ;
        RECT 9.720 90.370 12.940 90.850 ;
        RECT 19.640 90.370 22.860 90.850 ;
        RECT -283.320 88.800 -279.300 90.180 ;
        RECT -273.400 88.800 -269.380 90.180 ;
        RECT -263.480 88.800 -259.460 90.180 ;
        RECT -253.560 88.800 -249.540 90.180 ;
        RECT -243.640 88.800 -239.620 90.180 ;
        RECT -233.720 88.800 -229.700 90.180 ;
        RECT -223.800 88.800 -219.780 90.180 ;
        RECT -213.880 88.800 -209.860 90.180 ;
        RECT -203.960 88.800 -199.940 90.180 ;
        RECT -194.040 88.800 -190.020 90.180 ;
        RECT -184.120 88.800 -180.100 90.180 ;
        RECT -174.200 88.800 -170.180 90.180 ;
        RECT -164.280 88.800 -160.260 90.180 ;
        RECT -154.360 88.800 -150.340 90.180 ;
        RECT -144.440 88.800 -140.420 90.180 ;
        RECT -134.520 88.800 -130.500 90.180 ;
        RECT -124.600 88.800 -120.580 90.180 ;
        RECT -114.680 88.800 -110.660 90.180 ;
        RECT -104.760 88.800 -100.740 90.180 ;
        RECT -94.840 88.800 -90.820 90.180 ;
        RECT -84.920 88.800 -80.900 90.180 ;
        RECT -75.000 88.800 -70.980 90.180 ;
        RECT -65.080 88.800 -61.060 90.180 ;
        RECT -55.160 88.800 -51.140 90.180 ;
        RECT -45.240 88.800 -41.220 90.180 ;
        RECT -35.320 88.800 -31.300 90.180 ;
        RECT -25.400 88.800 -21.380 90.180 ;
        RECT -15.480 88.800 -11.460 90.180 ;
        RECT -5.560 88.800 -1.540 90.180 ;
        RECT 4.360 88.800 8.380 90.180 ;
        RECT 14.280 88.800 18.300 90.180 ;
        RECT -290.300 9.710 -286.280 11.090 ;
        RECT -280.380 9.710 -276.360 11.090 ;
        RECT -270.460 9.710 -266.440 11.090 ;
        RECT -260.540 9.710 -256.520 11.090 ;
        RECT -250.620 9.710 -246.600 11.090 ;
        RECT -240.700 9.710 -236.680 11.090 ;
        RECT -230.780 9.710 -226.760 11.090 ;
        RECT -220.860 9.710 -216.840 11.090 ;
        RECT -210.940 9.710 -206.920 11.090 ;
        RECT -201.020 9.710 -197.000 11.090 ;
        RECT -191.100 9.710 -187.080 11.090 ;
        RECT -181.180 9.710 -177.160 11.090 ;
        RECT -171.260 9.710 -167.240 11.090 ;
        RECT -161.340 9.710 -157.320 11.090 ;
        RECT -151.420 9.710 -147.400 11.090 ;
        RECT -141.500 9.710 -137.480 11.090 ;
        RECT -131.580 9.710 -127.560 11.090 ;
        RECT -121.660 9.710 -117.640 11.090 ;
        RECT -111.740 9.710 -107.720 11.090 ;
        RECT -101.820 9.710 -97.800 11.090 ;
        RECT -91.900 9.710 -87.880 11.090 ;
        RECT -81.980 9.710 -77.960 11.090 ;
        RECT -72.060 9.710 -68.040 11.090 ;
        RECT -62.140 9.710 -58.120 11.090 ;
        RECT -52.220 9.710 -48.200 11.090 ;
        RECT -42.300 9.710 -38.280 11.090 ;
        RECT -32.380 9.710 -28.360 11.090 ;
        RECT -22.460 9.710 -18.440 11.090 ;
        RECT -12.540 9.710 -8.520 11.090 ;
        RECT -2.620 9.710 1.400 11.090 ;
        RECT 7.300 9.710 11.320 11.090 ;
        RECT 17.220 9.710 21.240 11.090 ;
        RECT -284.940 9.040 -281.720 9.520 ;
        RECT -275.020 9.040 -271.800 9.520 ;
        RECT -265.100 9.040 -261.880 9.520 ;
        RECT -255.180 9.040 -251.960 9.520 ;
        RECT -245.260 9.040 -242.040 9.520 ;
        RECT -235.340 9.040 -232.120 9.520 ;
        RECT -225.420 9.040 -222.200 9.520 ;
        RECT -215.500 9.040 -212.280 9.520 ;
        RECT -205.580 9.040 -202.360 9.520 ;
        RECT -195.660 9.040 -192.440 9.520 ;
        RECT -185.740 9.040 -182.520 9.520 ;
        RECT -175.820 9.040 -172.600 9.520 ;
        RECT -165.900 9.040 -162.680 9.520 ;
        RECT -155.980 9.040 -152.760 9.520 ;
        RECT -146.060 9.040 -142.840 9.520 ;
        RECT -136.140 9.040 -132.920 9.520 ;
        RECT -126.220 9.040 -123.000 9.520 ;
        RECT -116.300 9.040 -113.080 9.520 ;
        RECT -106.380 9.040 -103.160 9.520 ;
        RECT -96.460 9.040 -93.240 9.520 ;
        RECT -86.540 9.040 -83.320 9.520 ;
        RECT -76.620 9.040 -73.400 9.520 ;
        RECT -66.700 9.040 -63.480 9.520 ;
        RECT -56.780 9.040 -53.560 9.520 ;
        RECT -46.860 9.040 -43.640 9.520 ;
        RECT -36.940 9.040 -33.720 9.520 ;
        RECT -27.020 9.040 -23.800 9.520 ;
        RECT -17.100 9.040 -13.880 9.520 ;
        RECT -7.180 9.040 -3.960 9.520 ;
        RECT 2.740 9.040 5.960 9.520 ;
        RECT 12.660 9.040 15.880 9.520 ;
        RECT -289.900 6.320 -286.680 6.800 ;
        RECT -279.980 6.320 -276.760 6.800 ;
        RECT -270.060 6.320 -266.840 6.800 ;
        RECT -260.140 6.320 -256.920 6.800 ;
        RECT -250.220 6.320 -247.000 6.800 ;
        RECT -240.300 6.320 -237.080 6.800 ;
        RECT -230.380 6.320 -227.160 6.800 ;
        RECT -220.460 6.320 -217.240 6.800 ;
        RECT -210.540 6.320 -207.320 6.800 ;
        RECT -200.620 6.320 -197.400 6.800 ;
        RECT -190.700 6.320 -187.480 6.800 ;
        RECT -180.780 6.320 -177.560 6.800 ;
        RECT -170.860 6.320 -167.640 6.800 ;
        RECT -160.940 6.320 -157.720 6.800 ;
        RECT -151.020 6.320 -147.800 6.800 ;
        RECT -141.100 6.320 -137.880 6.800 ;
        RECT -131.180 6.320 -127.960 6.800 ;
        RECT -121.260 6.320 -118.040 6.800 ;
        RECT -111.340 6.320 -108.120 6.800 ;
        RECT -101.420 6.320 -98.200 6.800 ;
        RECT -91.500 6.320 -88.280 6.800 ;
        RECT -81.580 6.320 -78.360 6.800 ;
        RECT -71.660 6.320 -68.440 6.800 ;
        RECT -61.740 6.320 -58.520 6.800 ;
        RECT -51.820 6.320 -48.600 6.800 ;
        RECT -41.900 6.320 -38.680 6.800 ;
        RECT -31.980 6.320 -28.760 6.800 ;
        RECT -22.060 6.320 -18.840 6.800 ;
        RECT -12.140 6.320 -8.920 6.800 ;
        RECT -2.220 6.320 1.000 6.800 ;
        RECT 7.700 6.320 10.920 6.800 ;
        RECT 17.620 6.320 20.840 6.800 ;
        RECT -285.340 4.750 -281.320 6.130 ;
        RECT -275.420 4.750 -271.400 6.130 ;
        RECT -265.500 4.750 -261.480 6.130 ;
        RECT -255.580 4.750 -251.560 6.130 ;
        RECT -245.660 4.750 -241.640 6.130 ;
        RECT -235.740 4.750 -231.720 6.130 ;
        RECT -225.820 4.750 -221.800 6.130 ;
        RECT -215.900 4.750 -211.880 6.130 ;
        RECT -205.980 4.750 -201.960 6.130 ;
        RECT -196.060 4.750 -192.040 6.130 ;
        RECT -186.140 4.750 -182.120 6.130 ;
        RECT -176.220 4.750 -172.200 6.130 ;
        RECT -166.300 4.750 -162.280 6.130 ;
        RECT -156.380 4.750 -152.360 6.130 ;
        RECT -146.460 4.750 -142.440 6.130 ;
        RECT -136.540 4.750 -132.520 6.130 ;
        RECT -126.620 4.750 -122.600 6.130 ;
        RECT -116.700 4.750 -112.680 6.130 ;
        RECT -106.780 4.750 -102.760 6.130 ;
        RECT -96.860 4.750 -92.840 6.130 ;
        RECT -86.940 4.750 -82.920 6.130 ;
        RECT -77.020 4.750 -73.000 6.130 ;
        RECT -67.100 4.750 -63.080 6.130 ;
        RECT -57.180 4.750 -53.160 6.130 ;
        RECT -47.260 4.750 -43.240 6.130 ;
        RECT -37.340 4.750 -33.320 6.130 ;
        RECT -27.420 4.750 -23.400 6.130 ;
        RECT -17.500 4.750 -13.480 6.130 ;
        RECT -7.580 4.750 -3.560 6.130 ;
        RECT 2.340 4.750 6.360 6.130 ;
        RECT 12.260 4.750 16.280 6.130 ;
        RECT -289.940 -79.240 -285.920 -77.860 ;
        RECT -280.020 -79.240 -276.000 -77.860 ;
        RECT -270.100 -79.240 -266.080 -77.860 ;
        RECT -260.180 -79.240 -256.160 -77.860 ;
        RECT -250.260 -79.240 -246.240 -77.860 ;
        RECT -240.340 -79.240 -236.320 -77.860 ;
        RECT -230.420 -79.240 -226.400 -77.860 ;
        RECT -220.500 -79.240 -216.480 -77.860 ;
        RECT -210.580 -79.240 -206.560 -77.860 ;
        RECT -200.660 -79.240 -196.640 -77.860 ;
        RECT -190.740 -79.240 -186.720 -77.860 ;
        RECT -180.820 -79.240 -176.800 -77.860 ;
        RECT -170.900 -79.240 -166.880 -77.860 ;
        RECT -160.980 -79.240 -156.960 -77.860 ;
        RECT -151.060 -79.240 -147.040 -77.860 ;
        RECT -141.140 -79.240 -137.120 -77.860 ;
        RECT -131.220 -79.240 -127.200 -77.860 ;
        RECT -121.300 -79.240 -117.280 -77.860 ;
        RECT -111.380 -79.240 -107.360 -77.860 ;
        RECT -101.460 -79.240 -97.440 -77.860 ;
        RECT -91.540 -79.240 -87.520 -77.860 ;
        RECT -81.620 -79.240 -77.600 -77.860 ;
        RECT -71.700 -79.240 -67.680 -77.860 ;
        RECT -61.780 -79.240 -57.760 -77.860 ;
        RECT -51.860 -79.240 -47.840 -77.860 ;
        RECT -41.940 -79.240 -37.920 -77.860 ;
        RECT -32.020 -79.240 -28.000 -77.860 ;
        RECT -22.100 -79.240 -18.080 -77.860 ;
        RECT -12.180 -79.240 -8.160 -77.860 ;
        RECT -2.260 -79.240 1.760 -77.860 ;
        RECT 7.660 -79.240 11.680 -77.860 ;
        RECT 17.580 -79.240 21.600 -77.860 ;
        RECT -284.580 -79.910 -281.360 -79.430 ;
        RECT -274.660 -79.910 -271.440 -79.430 ;
        RECT -264.740 -79.910 -261.520 -79.430 ;
        RECT -254.820 -79.910 -251.600 -79.430 ;
        RECT -244.900 -79.910 -241.680 -79.430 ;
        RECT -234.980 -79.910 -231.760 -79.430 ;
        RECT -225.060 -79.910 -221.840 -79.430 ;
        RECT -215.140 -79.910 -211.920 -79.430 ;
        RECT -205.220 -79.910 -202.000 -79.430 ;
        RECT -195.300 -79.910 -192.080 -79.430 ;
        RECT -185.380 -79.910 -182.160 -79.430 ;
        RECT -175.460 -79.910 -172.240 -79.430 ;
        RECT -165.540 -79.910 -162.320 -79.430 ;
        RECT -155.620 -79.910 -152.400 -79.430 ;
        RECT -145.700 -79.910 -142.480 -79.430 ;
        RECT -135.780 -79.910 -132.560 -79.430 ;
        RECT -125.860 -79.910 -122.640 -79.430 ;
        RECT -115.940 -79.910 -112.720 -79.430 ;
        RECT -106.020 -79.910 -102.800 -79.430 ;
        RECT -96.100 -79.910 -92.880 -79.430 ;
        RECT -86.180 -79.910 -82.960 -79.430 ;
        RECT -76.260 -79.910 -73.040 -79.430 ;
        RECT -66.340 -79.910 -63.120 -79.430 ;
        RECT -56.420 -79.910 -53.200 -79.430 ;
        RECT -46.500 -79.910 -43.280 -79.430 ;
        RECT -36.580 -79.910 -33.360 -79.430 ;
        RECT -26.660 -79.910 -23.440 -79.430 ;
        RECT -16.740 -79.910 -13.520 -79.430 ;
        RECT -6.820 -79.910 -3.600 -79.430 ;
        RECT 3.100 -79.910 6.320 -79.430 ;
        RECT 13.020 -79.910 16.240 -79.430 ;
        RECT -289.540 -82.630 -286.320 -82.150 ;
        RECT -279.620 -82.630 -276.400 -82.150 ;
        RECT -269.700 -82.630 -266.480 -82.150 ;
        RECT -259.780 -82.630 -256.560 -82.150 ;
        RECT -249.860 -82.630 -246.640 -82.150 ;
        RECT -239.940 -82.630 -236.720 -82.150 ;
        RECT -230.020 -82.630 -226.800 -82.150 ;
        RECT -220.100 -82.630 -216.880 -82.150 ;
        RECT -210.180 -82.630 -206.960 -82.150 ;
        RECT -200.260 -82.630 -197.040 -82.150 ;
        RECT -190.340 -82.630 -187.120 -82.150 ;
        RECT -180.420 -82.630 -177.200 -82.150 ;
        RECT -170.500 -82.630 -167.280 -82.150 ;
        RECT -160.580 -82.630 -157.360 -82.150 ;
        RECT -150.660 -82.630 -147.440 -82.150 ;
        RECT -140.740 -82.630 -137.520 -82.150 ;
        RECT -130.820 -82.630 -127.600 -82.150 ;
        RECT -120.900 -82.630 -117.680 -82.150 ;
        RECT -110.980 -82.630 -107.760 -82.150 ;
        RECT -101.060 -82.630 -97.840 -82.150 ;
        RECT -91.140 -82.630 -87.920 -82.150 ;
        RECT -81.220 -82.630 -78.000 -82.150 ;
        RECT -71.300 -82.630 -68.080 -82.150 ;
        RECT -61.380 -82.630 -58.160 -82.150 ;
        RECT -51.460 -82.630 -48.240 -82.150 ;
        RECT -41.540 -82.630 -38.320 -82.150 ;
        RECT -31.620 -82.630 -28.400 -82.150 ;
        RECT -21.700 -82.630 -18.480 -82.150 ;
        RECT -11.780 -82.630 -8.560 -82.150 ;
        RECT -1.860 -82.630 1.360 -82.150 ;
        RECT 8.060 -82.630 11.280 -82.150 ;
        RECT 17.980 -82.630 21.200 -82.150 ;
        RECT -284.980 -84.200 -280.960 -82.820 ;
        RECT -275.060 -84.200 -271.040 -82.820 ;
        RECT -265.140 -84.200 -261.120 -82.820 ;
        RECT -255.220 -84.200 -251.200 -82.820 ;
        RECT -245.300 -84.200 -241.280 -82.820 ;
        RECT -235.380 -84.200 -231.360 -82.820 ;
        RECT -225.460 -84.200 -221.440 -82.820 ;
        RECT -215.540 -84.200 -211.520 -82.820 ;
        RECT -205.620 -84.200 -201.600 -82.820 ;
        RECT -195.700 -84.200 -191.680 -82.820 ;
        RECT -185.780 -84.200 -181.760 -82.820 ;
        RECT -175.860 -84.200 -171.840 -82.820 ;
        RECT -165.940 -84.200 -161.920 -82.820 ;
        RECT -156.020 -84.200 -152.000 -82.820 ;
        RECT -146.100 -84.200 -142.080 -82.820 ;
        RECT -136.180 -84.200 -132.160 -82.820 ;
        RECT -126.260 -84.200 -122.240 -82.820 ;
        RECT -116.340 -84.200 -112.320 -82.820 ;
        RECT -106.420 -84.200 -102.400 -82.820 ;
        RECT -96.500 -84.200 -92.480 -82.820 ;
        RECT -86.580 -84.200 -82.560 -82.820 ;
        RECT -76.660 -84.200 -72.640 -82.820 ;
        RECT -66.740 -84.200 -62.720 -82.820 ;
        RECT -56.820 -84.200 -52.800 -82.820 ;
        RECT -46.900 -84.200 -42.880 -82.820 ;
        RECT -36.980 -84.200 -32.960 -82.820 ;
        RECT -27.060 -84.200 -23.040 -82.820 ;
        RECT -17.140 -84.200 -13.120 -82.820 ;
        RECT -7.220 -84.200 -3.200 -82.820 ;
        RECT 2.700 -84.200 6.720 -82.820 ;
        RECT 12.620 -84.200 16.640 -82.820 ;
        RECT -291.700 -173.820 -287.680 -172.440 ;
        RECT -281.780 -173.820 -277.760 -172.440 ;
        RECT -271.860 -173.820 -267.840 -172.440 ;
        RECT -261.940 -173.820 -257.920 -172.440 ;
        RECT -252.020 -173.820 -248.000 -172.440 ;
        RECT -242.100 -173.820 -238.080 -172.440 ;
        RECT -232.180 -173.820 -228.160 -172.440 ;
        RECT -222.260 -173.820 -218.240 -172.440 ;
        RECT -212.340 -173.820 -208.320 -172.440 ;
        RECT -202.420 -173.820 -198.400 -172.440 ;
        RECT -192.500 -173.820 -188.480 -172.440 ;
        RECT -182.580 -173.820 -178.560 -172.440 ;
        RECT -172.660 -173.820 -168.640 -172.440 ;
        RECT -162.740 -173.820 -158.720 -172.440 ;
        RECT -152.820 -173.820 -148.800 -172.440 ;
        RECT -142.900 -173.820 -138.880 -172.440 ;
        RECT -132.980 -173.820 -128.960 -172.440 ;
        RECT -123.060 -173.820 -119.040 -172.440 ;
        RECT -113.140 -173.820 -109.120 -172.440 ;
        RECT -103.220 -173.820 -99.200 -172.440 ;
        RECT -93.300 -173.820 -89.280 -172.440 ;
        RECT -83.380 -173.820 -79.360 -172.440 ;
        RECT -73.460 -173.820 -69.440 -172.440 ;
        RECT -63.540 -173.820 -59.520 -172.440 ;
        RECT -53.620 -173.820 -49.600 -172.440 ;
        RECT -43.700 -173.820 -39.680 -172.440 ;
        RECT -33.780 -173.820 -29.760 -172.440 ;
        RECT -23.860 -173.820 -19.840 -172.440 ;
        RECT -13.940 -173.820 -9.920 -172.440 ;
        RECT -4.020 -173.820 0.000 -172.440 ;
        RECT 5.900 -173.820 9.920 -172.440 ;
        RECT 15.820 -173.820 19.840 -172.440 ;
        RECT -286.340 -174.490 -283.120 -174.010 ;
        RECT -276.420 -174.490 -273.200 -174.010 ;
        RECT -266.500 -174.490 -263.280 -174.010 ;
        RECT -256.580 -174.490 -253.360 -174.010 ;
        RECT -246.660 -174.490 -243.440 -174.010 ;
        RECT -236.740 -174.490 -233.520 -174.010 ;
        RECT -226.820 -174.490 -223.600 -174.010 ;
        RECT -216.900 -174.490 -213.680 -174.010 ;
        RECT -206.980 -174.490 -203.760 -174.010 ;
        RECT -197.060 -174.490 -193.840 -174.010 ;
        RECT -187.140 -174.490 -183.920 -174.010 ;
        RECT -177.220 -174.490 -174.000 -174.010 ;
        RECT -167.300 -174.490 -164.080 -174.010 ;
        RECT -157.380 -174.490 -154.160 -174.010 ;
        RECT -147.460 -174.490 -144.240 -174.010 ;
        RECT -137.540 -174.490 -134.320 -174.010 ;
        RECT -127.620 -174.490 -124.400 -174.010 ;
        RECT -117.700 -174.490 -114.480 -174.010 ;
        RECT -107.780 -174.490 -104.560 -174.010 ;
        RECT -97.860 -174.490 -94.640 -174.010 ;
        RECT -87.940 -174.490 -84.720 -174.010 ;
        RECT -78.020 -174.490 -74.800 -174.010 ;
        RECT -68.100 -174.490 -64.880 -174.010 ;
        RECT -58.180 -174.490 -54.960 -174.010 ;
        RECT -48.260 -174.490 -45.040 -174.010 ;
        RECT -38.340 -174.490 -35.120 -174.010 ;
        RECT -28.420 -174.490 -25.200 -174.010 ;
        RECT -18.500 -174.490 -15.280 -174.010 ;
        RECT -8.580 -174.490 -5.360 -174.010 ;
        RECT 1.340 -174.490 4.560 -174.010 ;
        RECT 11.260 -174.490 14.480 -174.010 ;
        RECT -291.300 -177.210 -288.080 -176.730 ;
        RECT -281.380 -177.210 -278.160 -176.730 ;
        RECT -271.460 -177.210 -268.240 -176.730 ;
        RECT -261.540 -177.210 -258.320 -176.730 ;
        RECT -251.620 -177.210 -248.400 -176.730 ;
        RECT -241.700 -177.210 -238.480 -176.730 ;
        RECT -231.780 -177.210 -228.560 -176.730 ;
        RECT -221.860 -177.210 -218.640 -176.730 ;
        RECT -211.940 -177.210 -208.720 -176.730 ;
        RECT -202.020 -177.210 -198.800 -176.730 ;
        RECT -192.100 -177.210 -188.880 -176.730 ;
        RECT -182.180 -177.210 -178.960 -176.730 ;
        RECT -172.260 -177.210 -169.040 -176.730 ;
        RECT -162.340 -177.210 -159.120 -176.730 ;
        RECT -152.420 -177.210 -149.200 -176.730 ;
        RECT -142.500 -177.210 -139.280 -176.730 ;
        RECT -132.580 -177.210 -129.360 -176.730 ;
        RECT -122.660 -177.210 -119.440 -176.730 ;
        RECT -112.740 -177.210 -109.520 -176.730 ;
        RECT -102.820 -177.210 -99.600 -176.730 ;
        RECT -92.900 -177.210 -89.680 -176.730 ;
        RECT -82.980 -177.210 -79.760 -176.730 ;
        RECT -73.060 -177.210 -69.840 -176.730 ;
        RECT -63.140 -177.210 -59.920 -176.730 ;
        RECT -53.220 -177.210 -50.000 -176.730 ;
        RECT -43.300 -177.210 -40.080 -176.730 ;
        RECT -33.380 -177.210 -30.160 -176.730 ;
        RECT -23.460 -177.210 -20.240 -176.730 ;
        RECT -13.540 -177.210 -10.320 -176.730 ;
        RECT -3.620 -177.210 -0.400 -176.730 ;
        RECT 6.300 -177.210 9.520 -176.730 ;
        RECT 16.220 -177.210 19.440 -176.730 ;
        RECT -286.740 -178.780 -282.720 -177.400 ;
        RECT -276.820 -178.780 -272.800 -177.400 ;
        RECT -266.900 -178.780 -262.880 -177.400 ;
        RECT -256.980 -178.780 -252.960 -177.400 ;
        RECT -247.060 -178.780 -243.040 -177.400 ;
        RECT -237.140 -178.780 -233.120 -177.400 ;
        RECT -227.220 -178.780 -223.200 -177.400 ;
        RECT -217.300 -178.780 -213.280 -177.400 ;
        RECT -207.380 -178.780 -203.360 -177.400 ;
        RECT -197.460 -178.780 -193.440 -177.400 ;
        RECT -187.540 -178.780 -183.520 -177.400 ;
        RECT -177.620 -178.780 -173.600 -177.400 ;
        RECT -167.700 -178.780 -163.680 -177.400 ;
        RECT -157.780 -178.780 -153.760 -177.400 ;
        RECT -147.860 -178.780 -143.840 -177.400 ;
        RECT -137.940 -178.780 -133.920 -177.400 ;
        RECT -128.020 -178.780 -124.000 -177.400 ;
        RECT -118.100 -178.780 -114.080 -177.400 ;
        RECT -108.180 -178.780 -104.160 -177.400 ;
        RECT -98.260 -178.780 -94.240 -177.400 ;
        RECT -88.340 -178.780 -84.320 -177.400 ;
        RECT -78.420 -178.780 -74.400 -177.400 ;
        RECT -68.500 -178.780 -64.480 -177.400 ;
        RECT -58.580 -178.780 -54.560 -177.400 ;
        RECT -48.660 -178.780 -44.640 -177.400 ;
        RECT -38.740 -178.780 -34.720 -177.400 ;
        RECT -28.820 -178.780 -24.800 -177.400 ;
        RECT -18.900 -178.780 -14.880 -177.400 ;
        RECT -8.980 -178.780 -4.960 -177.400 ;
        RECT 0.940 -178.780 4.960 -177.400 ;
        RECT 10.860 -178.780 14.880 -177.400 ;
      LAYER via ;
        RECT -287.700 94.070 -287.425 94.335 ;
        RECT -277.780 94.070 -277.505 94.335 ;
        RECT -267.860 94.070 -267.585 94.335 ;
        RECT -257.940 94.070 -257.665 94.335 ;
        RECT -248.020 94.070 -247.745 94.335 ;
        RECT -238.100 94.070 -237.825 94.335 ;
        RECT -228.180 94.070 -227.905 94.335 ;
        RECT -218.260 94.070 -217.985 94.335 ;
        RECT -208.340 94.070 -208.065 94.335 ;
        RECT -198.420 94.070 -198.145 94.335 ;
        RECT -188.500 94.070 -188.225 94.335 ;
        RECT -178.580 94.070 -178.305 94.335 ;
        RECT -168.660 94.070 -168.385 94.335 ;
        RECT -158.740 94.070 -158.465 94.335 ;
        RECT -148.820 94.070 -148.545 94.335 ;
        RECT -138.900 94.070 -138.625 94.335 ;
        RECT -128.980 94.070 -128.705 94.335 ;
        RECT -119.060 94.070 -118.785 94.335 ;
        RECT -109.140 94.070 -108.865 94.335 ;
        RECT -99.220 94.070 -98.945 94.335 ;
        RECT -89.300 94.070 -89.025 94.335 ;
        RECT -79.380 94.070 -79.105 94.335 ;
        RECT -69.460 94.070 -69.185 94.335 ;
        RECT -59.540 94.070 -59.265 94.335 ;
        RECT -49.620 94.070 -49.345 94.335 ;
        RECT -39.700 94.070 -39.425 94.335 ;
        RECT -29.780 94.070 -29.505 94.335 ;
        RECT -19.860 94.070 -19.585 94.335 ;
        RECT -9.940 94.070 -9.665 94.335 ;
        RECT -0.020 94.070 0.255 94.335 ;
        RECT 9.900 94.070 10.175 94.335 ;
        RECT 19.820 94.070 20.095 94.335 ;
        RECT -280.530 93.200 -280.255 93.465 ;
        RECT -280.060 93.200 -279.785 93.465 ;
        RECT -270.610 93.200 -270.335 93.465 ;
        RECT -270.140 93.200 -269.865 93.465 ;
        RECT -260.690 93.200 -260.415 93.465 ;
        RECT -260.220 93.200 -259.945 93.465 ;
        RECT -250.770 93.200 -250.495 93.465 ;
        RECT -250.300 93.200 -250.025 93.465 ;
        RECT -240.850 93.200 -240.575 93.465 ;
        RECT -240.380 93.200 -240.105 93.465 ;
        RECT -230.930 93.200 -230.655 93.465 ;
        RECT -230.460 93.200 -230.185 93.465 ;
        RECT -221.010 93.200 -220.735 93.465 ;
        RECT -220.540 93.200 -220.265 93.465 ;
        RECT -211.090 93.200 -210.815 93.465 ;
        RECT -210.620 93.200 -210.345 93.465 ;
        RECT -201.170 93.200 -200.895 93.465 ;
        RECT -200.700 93.200 -200.425 93.465 ;
        RECT -191.250 93.200 -190.975 93.465 ;
        RECT -190.780 93.200 -190.505 93.465 ;
        RECT -181.330 93.200 -181.055 93.465 ;
        RECT -180.860 93.200 -180.585 93.465 ;
        RECT -171.410 93.200 -171.135 93.465 ;
        RECT -170.940 93.200 -170.665 93.465 ;
        RECT -161.490 93.200 -161.215 93.465 ;
        RECT -161.020 93.200 -160.745 93.465 ;
        RECT -151.570 93.200 -151.295 93.465 ;
        RECT -151.100 93.200 -150.825 93.465 ;
        RECT -141.650 93.200 -141.375 93.465 ;
        RECT -141.180 93.200 -140.905 93.465 ;
        RECT -131.730 93.200 -131.455 93.465 ;
        RECT -131.260 93.200 -130.985 93.465 ;
        RECT -121.810 93.200 -121.535 93.465 ;
        RECT -121.340 93.200 -121.065 93.465 ;
        RECT -111.890 93.200 -111.615 93.465 ;
        RECT -111.420 93.200 -111.145 93.465 ;
        RECT -101.970 93.200 -101.695 93.465 ;
        RECT -101.500 93.200 -101.225 93.465 ;
        RECT -92.050 93.200 -91.775 93.465 ;
        RECT -91.580 93.200 -91.305 93.465 ;
        RECT -82.130 93.200 -81.855 93.465 ;
        RECT -81.660 93.200 -81.385 93.465 ;
        RECT -72.210 93.200 -71.935 93.465 ;
        RECT -71.740 93.200 -71.465 93.465 ;
        RECT -62.290 93.200 -62.015 93.465 ;
        RECT -61.820 93.200 -61.545 93.465 ;
        RECT -52.370 93.200 -52.095 93.465 ;
        RECT -51.900 93.200 -51.625 93.465 ;
        RECT -42.450 93.200 -42.175 93.465 ;
        RECT -41.980 93.200 -41.705 93.465 ;
        RECT -32.530 93.200 -32.255 93.465 ;
        RECT -32.060 93.200 -31.785 93.465 ;
        RECT -22.610 93.200 -22.335 93.465 ;
        RECT -22.140 93.200 -21.865 93.465 ;
        RECT -12.690 93.200 -12.415 93.465 ;
        RECT -12.220 93.200 -11.945 93.465 ;
        RECT -2.770 93.200 -2.495 93.465 ;
        RECT -2.300 93.200 -2.025 93.465 ;
        RECT 7.150 93.200 7.425 93.465 ;
        RECT 7.620 93.200 7.895 93.465 ;
        RECT 17.070 93.200 17.345 93.465 ;
        RECT 17.540 93.200 17.815 93.465 ;
        RECT -287.790 90.470 -287.515 90.735 ;
        RECT -287.330 90.480 -287.055 90.745 ;
        RECT -277.870 90.470 -277.595 90.735 ;
        RECT -277.410 90.480 -277.135 90.745 ;
        RECT -267.950 90.470 -267.675 90.735 ;
        RECT -267.490 90.480 -267.215 90.745 ;
        RECT -258.030 90.470 -257.755 90.735 ;
        RECT -257.570 90.480 -257.295 90.745 ;
        RECT -248.110 90.470 -247.835 90.735 ;
        RECT -247.650 90.480 -247.375 90.745 ;
        RECT -238.190 90.470 -237.915 90.735 ;
        RECT -237.730 90.480 -237.455 90.745 ;
        RECT -228.270 90.470 -227.995 90.735 ;
        RECT -227.810 90.480 -227.535 90.745 ;
        RECT -218.350 90.470 -218.075 90.735 ;
        RECT -217.890 90.480 -217.615 90.745 ;
        RECT -208.430 90.470 -208.155 90.735 ;
        RECT -207.970 90.480 -207.695 90.745 ;
        RECT -198.510 90.470 -198.235 90.735 ;
        RECT -198.050 90.480 -197.775 90.745 ;
        RECT -188.590 90.470 -188.315 90.735 ;
        RECT -188.130 90.480 -187.855 90.745 ;
        RECT -178.670 90.470 -178.395 90.735 ;
        RECT -178.210 90.480 -177.935 90.745 ;
        RECT -168.750 90.470 -168.475 90.735 ;
        RECT -168.290 90.480 -168.015 90.745 ;
        RECT -158.830 90.470 -158.555 90.735 ;
        RECT -158.370 90.480 -158.095 90.745 ;
        RECT -148.910 90.470 -148.635 90.735 ;
        RECT -148.450 90.480 -148.175 90.745 ;
        RECT -138.990 90.470 -138.715 90.735 ;
        RECT -138.530 90.480 -138.255 90.745 ;
        RECT -129.070 90.470 -128.795 90.735 ;
        RECT -128.610 90.480 -128.335 90.745 ;
        RECT -119.150 90.470 -118.875 90.735 ;
        RECT -118.690 90.480 -118.415 90.745 ;
        RECT -109.230 90.470 -108.955 90.735 ;
        RECT -108.770 90.480 -108.495 90.745 ;
        RECT -99.310 90.470 -99.035 90.735 ;
        RECT -98.850 90.480 -98.575 90.745 ;
        RECT -89.390 90.470 -89.115 90.735 ;
        RECT -88.930 90.480 -88.655 90.745 ;
        RECT -79.470 90.470 -79.195 90.735 ;
        RECT -79.010 90.480 -78.735 90.745 ;
        RECT -69.550 90.470 -69.275 90.735 ;
        RECT -69.090 90.480 -68.815 90.745 ;
        RECT -59.630 90.470 -59.355 90.735 ;
        RECT -59.170 90.480 -58.895 90.745 ;
        RECT -49.710 90.470 -49.435 90.735 ;
        RECT -49.250 90.480 -48.975 90.745 ;
        RECT -39.790 90.470 -39.515 90.735 ;
        RECT -39.330 90.480 -39.055 90.745 ;
        RECT -29.870 90.470 -29.595 90.735 ;
        RECT -29.410 90.480 -29.135 90.745 ;
        RECT -19.950 90.470 -19.675 90.735 ;
        RECT -19.490 90.480 -19.215 90.745 ;
        RECT -10.030 90.470 -9.755 90.735 ;
        RECT -9.570 90.480 -9.295 90.745 ;
        RECT -0.110 90.470 0.165 90.735 ;
        RECT 0.350 90.480 0.625 90.745 ;
        RECT 9.810 90.470 10.085 90.735 ;
        RECT 10.270 90.480 10.545 90.745 ;
        RECT 19.730 90.470 20.005 90.735 ;
        RECT 20.190 90.480 20.465 90.745 ;
        RECT -280.140 89.710 -279.865 89.975 ;
        RECT -270.220 89.710 -269.945 89.975 ;
        RECT -260.300 89.710 -260.025 89.975 ;
        RECT -250.380 89.710 -250.105 89.975 ;
        RECT -240.460 89.710 -240.185 89.975 ;
        RECT -230.540 89.710 -230.265 89.975 ;
        RECT -220.620 89.710 -220.345 89.975 ;
        RECT -210.700 89.710 -210.425 89.975 ;
        RECT -200.780 89.710 -200.505 89.975 ;
        RECT -190.860 89.710 -190.585 89.975 ;
        RECT -180.940 89.710 -180.665 89.975 ;
        RECT -171.020 89.710 -170.745 89.975 ;
        RECT -161.100 89.710 -160.825 89.975 ;
        RECT -151.180 89.710 -150.905 89.975 ;
        RECT -141.260 89.710 -140.985 89.975 ;
        RECT -131.340 89.710 -131.065 89.975 ;
        RECT -121.420 89.710 -121.145 89.975 ;
        RECT -111.500 89.710 -111.225 89.975 ;
        RECT -101.580 89.710 -101.305 89.975 ;
        RECT -91.660 89.710 -91.385 89.975 ;
        RECT -81.740 89.710 -81.465 89.975 ;
        RECT -71.820 89.710 -71.545 89.975 ;
        RECT -61.900 89.710 -61.625 89.975 ;
        RECT -51.980 89.710 -51.705 89.975 ;
        RECT -42.060 89.710 -41.785 89.975 ;
        RECT -32.140 89.710 -31.865 89.975 ;
        RECT -22.220 89.710 -21.945 89.975 ;
        RECT -12.300 89.710 -12.025 89.975 ;
        RECT -2.380 89.710 -2.105 89.975 ;
        RECT 7.540 89.710 7.815 89.975 ;
        RECT 17.460 89.710 17.735 89.975 ;
        RECT -289.720 10.020 -289.445 10.285 ;
        RECT -279.800 10.020 -279.525 10.285 ;
        RECT -269.880 10.020 -269.605 10.285 ;
        RECT -259.960 10.020 -259.685 10.285 ;
        RECT -250.040 10.020 -249.765 10.285 ;
        RECT -240.120 10.020 -239.845 10.285 ;
        RECT -230.200 10.020 -229.925 10.285 ;
        RECT -220.280 10.020 -220.005 10.285 ;
        RECT -210.360 10.020 -210.085 10.285 ;
        RECT -200.440 10.020 -200.165 10.285 ;
        RECT -190.520 10.020 -190.245 10.285 ;
        RECT -180.600 10.020 -180.325 10.285 ;
        RECT -170.680 10.020 -170.405 10.285 ;
        RECT -160.760 10.020 -160.485 10.285 ;
        RECT -150.840 10.020 -150.565 10.285 ;
        RECT -140.920 10.020 -140.645 10.285 ;
        RECT -131.000 10.020 -130.725 10.285 ;
        RECT -121.080 10.020 -120.805 10.285 ;
        RECT -111.160 10.020 -110.885 10.285 ;
        RECT -101.240 10.020 -100.965 10.285 ;
        RECT -91.320 10.020 -91.045 10.285 ;
        RECT -81.400 10.020 -81.125 10.285 ;
        RECT -71.480 10.020 -71.205 10.285 ;
        RECT -61.560 10.020 -61.285 10.285 ;
        RECT -51.640 10.020 -51.365 10.285 ;
        RECT -41.720 10.020 -41.445 10.285 ;
        RECT -31.800 10.020 -31.525 10.285 ;
        RECT -21.880 10.020 -21.605 10.285 ;
        RECT -11.960 10.020 -11.685 10.285 ;
        RECT -2.040 10.020 -1.765 10.285 ;
        RECT 7.880 10.020 8.155 10.285 ;
        RECT 17.800 10.020 18.075 10.285 ;
        RECT -282.550 9.150 -282.275 9.415 ;
        RECT -282.080 9.150 -281.805 9.415 ;
        RECT -272.630 9.150 -272.355 9.415 ;
        RECT -272.160 9.150 -271.885 9.415 ;
        RECT -262.710 9.150 -262.435 9.415 ;
        RECT -262.240 9.150 -261.965 9.415 ;
        RECT -252.790 9.150 -252.515 9.415 ;
        RECT -252.320 9.150 -252.045 9.415 ;
        RECT -242.870 9.150 -242.595 9.415 ;
        RECT -242.400 9.150 -242.125 9.415 ;
        RECT -232.950 9.150 -232.675 9.415 ;
        RECT -232.480 9.150 -232.205 9.415 ;
        RECT -223.030 9.150 -222.755 9.415 ;
        RECT -222.560 9.150 -222.285 9.415 ;
        RECT -213.110 9.150 -212.835 9.415 ;
        RECT -212.640 9.150 -212.365 9.415 ;
        RECT -203.190 9.150 -202.915 9.415 ;
        RECT -202.720 9.150 -202.445 9.415 ;
        RECT -193.270 9.150 -192.995 9.415 ;
        RECT -192.800 9.150 -192.525 9.415 ;
        RECT -183.350 9.150 -183.075 9.415 ;
        RECT -182.880 9.150 -182.605 9.415 ;
        RECT -173.430 9.150 -173.155 9.415 ;
        RECT -172.960 9.150 -172.685 9.415 ;
        RECT -163.510 9.150 -163.235 9.415 ;
        RECT -163.040 9.150 -162.765 9.415 ;
        RECT -153.590 9.150 -153.315 9.415 ;
        RECT -153.120 9.150 -152.845 9.415 ;
        RECT -143.670 9.150 -143.395 9.415 ;
        RECT -143.200 9.150 -142.925 9.415 ;
        RECT -133.750 9.150 -133.475 9.415 ;
        RECT -133.280 9.150 -133.005 9.415 ;
        RECT -123.830 9.150 -123.555 9.415 ;
        RECT -123.360 9.150 -123.085 9.415 ;
        RECT -113.910 9.150 -113.635 9.415 ;
        RECT -113.440 9.150 -113.165 9.415 ;
        RECT -103.990 9.150 -103.715 9.415 ;
        RECT -103.520 9.150 -103.245 9.415 ;
        RECT -94.070 9.150 -93.795 9.415 ;
        RECT -93.600 9.150 -93.325 9.415 ;
        RECT -84.150 9.150 -83.875 9.415 ;
        RECT -83.680 9.150 -83.405 9.415 ;
        RECT -74.230 9.150 -73.955 9.415 ;
        RECT -73.760 9.150 -73.485 9.415 ;
        RECT -64.310 9.150 -64.035 9.415 ;
        RECT -63.840 9.150 -63.565 9.415 ;
        RECT -54.390 9.150 -54.115 9.415 ;
        RECT -53.920 9.150 -53.645 9.415 ;
        RECT -44.470 9.150 -44.195 9.415 ;
        RECT -44.000 9.150 -43.725 9.415 ;
        RECT -34.550 9.150 -34.275 9.415 ;
        RECT -34.080 9.150 -33.805 9.415 ;
        RECT -24.630 9.150 -24.355 9.415 ;
        RECT -24.160 9.150 -23.885 9.415 ;
        RECT -14.710 9.150 -14.435 9.415 ;
        RECT -14.240 9.150 -13.965 9.415 ;
        RECT -4.790 9.150 -4.515 9.415 ;
        RECT -4.320 9.150 -4.045 9.415 ;
        RECT 5.130 9.150 5.405 9.415 ;
        RECT 5.600 9.150 5.875 9.415 ;
        RECT 15.050 9.150 15.325 9.415 ;
        RECT 15.520 9.150 15.795 9.415 ;
        RECT -289.810 6.420 -289.535 6.685 ;
        RECT -289.350 6.430 -289.075 6.695 ;
        RECT -279.890 6.420 -279.615 6.685 ;
        RECT -279.430 6.430 -279.155 6.695 ;
        RECT -269.970 6.420 -269.695 6.685 ;
        RECT -269.510 6.430 -269.235 6.695 ;
        RECT -260.050 6.420 -259.775 6.685 ;
        RECT -259.590 6.430 -259.315 6.695 ;
        RECT -250.130 6.420 -249.855 6.685 ;
        RECT -249.670 6.430 -249.395 6.695 ;
        RECT -240.210 6.420 -239.935 6.685 ;
        RECT -239.750 6.430 -239.475 6.695 ;
        RECT -230.290 6.420 -230.015 6.685 ;
        RECT -229.830 6.430 -229.555 6.695 ;
        RECT -220.370 6.420 -220.095 6.685 ;
        RECT -219.910 6.430 -219.635 6.695 ;
        RECT -210.450 6.420 -210.175 6.685 ;
        RECT -209.990 6.430 -209.715 6.695 ;
        RECT -200.530 6.420 -200.255 6.685 ;
        RECT -200.070 6.430 -199.795 6.695 ;
        RECT -190.610 6.420 -190.335 6.685 ;
        RECT -190.150 6.430 -189.875 6.695 ;
        RECT -180.690 6.420 -180.415 6.685 ;
        RECT -180.230 6.430 -179.955 6.695 ;
        RECT -170.770 6.420 -170.495 6.685 ;
        RECT -170.310 6.430 -170.035 6.695 ;
        RECT -160.850 6.420 -160.575 6.685 ;
        RECT -160.390 6.430 -160.115 6.695 ;
        RECT -150.930 6.420 -150.655 6.685 ;
        RECT -150.470 6.430 -150.195 6.695 ;
        RECT -141.010 6.420 -140.735 6.685 ;
        RECT -140.550 6.430 -140.275 6.695 ;
        RECT -131.090 6.420 -130.815 6.685 ;
        RECT -130.630 6.430 -130.355 6.695 ;
        RECT -121.170 6.420 -120.895 6.685 ;
        RECT -120.710 6.430 -120.435 6.695 ;
        RECT -111.250 6.420 -110.975 6.685 ;
        RECT -110.790 6.430 -110.515 6.695 ;
        RECT -101.330 6.420 -101.055 6.685 ;
        RECT -100.870 6.430 -100.595 6.695 ;
        RECT -91.410 6.420 -91.135 6.685 ;
        RECT -90.950 6.430 -90.675 6.695 ;
        RECT -81.490 6.420 -81.215 6.685 ;
        RECT -81.030 6.430 -80.755 6.695 ;
        RECT -71.570 6.420 -71.295 6.685 ;
        RECT -71.110 6.430 -70.835 6.695 ;
        RECT -61.650 6.420 -61.375 6.685 ;
        RECT -61.190 6.430 -60.915 6.695 ;
        RECT -51.730 6.420 -51.455 6.685 ;
        RECT -51.270 6.430 -50.995 6.695 ;
        RECT -41.810 6.420 -41.535 6.685 ;
        RECT -41.350 6.430 -41.075 6.695 ;
        RECT -31.890 6.420 -31.615 6.685 ;
        RECT -31.430 6.430 -31.155 6.695 ;
        RECT -21.970 6.420 -21.695 6.685 ;
        RECT -21.510 6.430 -21.235 6.695 ;
        RECT -12.050 6.420 -11.775 6.685 ;
        RECT -11.590 6.430 -11.315 6.695 ;
        RECT -2.130 6.420 -1.855 6.685 ;
        RECT -1.670 6.430 -1.395 6.695 ;
        RECT 7.790 6.420 8.065 6.685 ;
        RECT 8.250 6.430 8.525 6.695 ;
        RECT 17.710 6.420 17.985 6.685 ;
        RECT 18.170 6.430 18.445 6.695 ;
        RECT -282.160 5.660 -281.885 5.925 ;
        RECT -272.240 5.660 -271.965 5.925 ;
        RECT -262.320 5.660 -262.045 5.925 ;
        RECT -252.400 5.660 -252.125 5.925 ;
        RECT -242.480 5.660 -242.205 5.925 ;
        RECT -232.560 5.660 -232.285 5.925 ;
        RECT -222.640 5.660 -222.365 5.925 ;
        RECT -212.720 5.660 -212.445 5.925 ;
        RECT -202.800 5.660 -202.525 5.925 ;
        RECT -192.880 5.660 -192.605 5.925 ;
        RECT -182.960 5.660 -182.685 5.925 ;
        RECT -173.040 5.660 -172.765 5.925 ;
        RECT -163.120 5.660 -162.845 5.925 ;
        RECT -153.200 5.660 -152.925 5.925 ;
        RECT -143.280 5.660 -143.005 5.925 ;
        RECT -133.360 5.660 -133.085 5.925 ;
        RECT -123.440 5.660 -123.165 5.925 ;
        RECT -113.520 5.660 -113.245 5.925 ;
        RECT -103.600 5.660 -103.325 5.925 ;
        RECT -93.680 5.660 -93.405 5.925 ;
        RECT -83.760 5.660 -83.485 5.925 ;
        RECT -73.840 5.660 -73.565 5.925 ;
        RECT -63.920 5.660 -63.645 5.925 ;
        RECT -54.000 5.660 -53.725 5.925 ;
        RECT -44.080 5.660 -43.805 5.925 ;
        RECT -34.160 5.660 -33.885 5.925 ;
        RECT -24.240 5.660 -23.965 5.925 ;
        RECT -14.320 5.660 -14.045 5.925 ;
        RECT -4.400 5.660 -4.125 5.925 ;
        RECT 5.520 5.660 5.795 5.925 ;
        RECT 15.440 5.660 15.715 5.925 ;
        RECT -289.360 -78.930 -289.085 -78.665 ;
        RECT -279.440 -78.930 -279.165 -78.665 ;
        RECT -269.520 -78.930 -269.245 -78.665 ;
        RECT -259.600 -78.930 -259.325 -78.665 ;
        RECT -249.680 -78.930 -249.405 -78.665 ;
        RECT -239.760 -78.930 -239.485 -78.665 ;
        RECT -229.840 -78.930 -229.565 -78.665 ;
        RECT -219.920 -78.930 -219.645 -78.665 ;
        RECT -210.000 -78.930 -209.725 -78.665 ;
        RECT -200.080 -78.930 -199.805 -78.665 ;
        RECT -190.160 -78.930 -189.885 -78.665 ;
        RECT -180.240 -78.930 -179.965 -78.665 ;
        RECT -170.320 -78.930 -170.045 -78.665 ;
        RECT -160.400 -78.930 -160.125 -78.665 ;
        RECT -150.480 -78.930 -150.205 -78.665 ;
        RECT -140.560 -78.930 -140.285 -78.665 ;
        RECT -130.640 -78.930 -130.365 -78.665 ;
        RECT -120.720 -78.930 -120.445 -78.665 ;
        RECT -110.800 -78.930 -110.525 -78.665 ;
        RECT -100.880 -78.930 -100.605 -78.665 ;
        RECT -90.960 -78.930 -90.685 -78.665 ;
        RECT -81.040 -78.930 -80.765 -78.665 ;
        RECT -71.120 -78.930 -70.845 -78.665 ;
        RECT -61.200 -78.930 -60.925 -78.665 ;
        RECT -51.280 -78.930 -51.005 -78.665 ;
        RECT -41.360 -78.930 -41.085 -78.665 ;
        RECT -31.440 -78.930 -31.165 -78.665 ;
        RECT -21.520 -78.930 -21.245 -78.665 ;
        RECT -11.600 -78.930 -11.325 -78.665 ;
        RECT -1.680 -78.930 -1.405 -78.665 ;
        RECT 8.240 -78.930 8.515 -78.665 ;
        RECT 18.160 -78.930 18.435 -78.665 ;
        RECT -282.190 -79.800 -281.915 -79.535 ;
        RECT -281.720 -79.800 -281.445 -79.535 ;
        RECT -272.270 -79.800 -271.995 -79.535 ;
        RECT -271.800 -79.800 -271.525 -79.535 ;
        RECT -262.350 -79.800 -262.075 -79.535 ;
        RECT -261.880 -79.800 -261.605 -79.535 ;
        RECT -252.430 -79.800 -252.155 -79.535 ;
        RECT -251.960 -79.800 -251.685 -79.535 ;
        RECT -242.510 -79.800 -242.235 -79.535 ;
        RECT -242.040 -79.800 -241.765 -79.535 ;
        RECT -232.590 -79.800 -232.315 -79.535 ;
        RECT -232.120 -79.800 -231.845 -79.535 ;
        RECT -222.670 -79.800 -222.395 -79.535 ;
        RECT -222.200 -79.800 -221.925 -79.535 ;
        RECT -212.750 -79.800 -212.475 -79.535 ;
        RECT -212.280 -79.800 -212.005 -79.535 ;
        RECT -202.830 -79.800 -202.555 -79.535 ;
        RECT -202.360 -79.800 -202.085 -79.535 ;
        RECT -192.910 -79.800 -192.635 -79.535 ;
        RECT -192.440 -79.800 -192.165 -79.535 ;
        RECT -182.990 -79.800 -182.715 -79.535 ;
        RECT -182.520 -79.800 -182.245 -79.535 ;
        RECT -173.070 -79.800 -172.795 -79.535 ;
        RECT -172.600 -79.800 -172.325 -79.535 ;
        RECT -163.150 -79.800 -162.875 -79.535 ;
        RECT -162.680 -79.800 -162.405 -79.535 ;
        RECT -153.230 -79.800 -152.955 -79.535 ;
        RECT -152.760 -79.800 -152.485 -79.535 ;
        RECT -143.310 -79.800 -143.035 -79.535 ;
        RECT -142.840 -79.800 -142.565 -79.535 ;
        RECT -133.390 -79.800 -133.115 -79.535 ;
        RECT -132.920 -79.800 -132.645 -79.535 ;
        RECT -123.470 -79.800 -123.195 -79.535 ;
        RECT -123.000 -79.800 -122.725 -79.535 ;
        RECT -113.550 -79.800 -113.275 -79.535 ;
        RECT -113.080 -79.800 -112.805 -79.535 ;
        RECT -103.630 -79.800 -103.355 -79.535 ;
        RECT -103.160 -79.800 -102.885 -79.535 ;
        RECT -93.710 -79.800 -93.435 -79.535 ;
        RECT -93.240 -79.800 -92.965 -79.535 ;
        RECT -83.790 -79.800 -83.515 -79.535 ;
        RECT -83.320 -79.800 -83.045 -79.535 ;
        RECT -73.870 -79.800 -73.595 -79.535 ;
        RECT -73.400 -79.800 -73.125 -79.535 ;
        RECT -63.950 -79.800 -63.675 -79.535 ;
        RECT -63.480 -79.800 -63.205 -79.535 ;
        RECT -54.030 -79.800 -53.755 -79.535 ;
        RECT -53.560 -79.800 -53.285 -79.535 ;
        RECT -44.110 -79.800 -43.835 -79.535 ;
        RECT -43.640 -79.800 -43.365 -79.535 ;
        RECT -34.190 -79.800 -33.915 -79.535 ;
        RECT -33.720 -79.800 -33.445 -79.535 ;
        RECT -24.270 -79.800 -23.995 -79.535 ;
        RECT -23.800 -79.800 -23.525 -79.535 ;
        RECT -14.350 -79.800 -14.075 -79.535 ;
        RECT -13.880 -79.800 -13.605 -79.535 ;
        RECT -4.430 -79.800 -4.155 -79.535 ;
        RECT -3.960 -79.800 -3.685 -79.535 ;
        RECT 5.490 -79.800 5.765 -79.535 ;
        RECT 5.960 -79.800 6.235 -79.535 ;
        RECT 15.410 -79.800 15.685 -79.535 ;
        RECT 15.880 -79.800 16.155 -79.535 ;
        RECT -289.450 -82.530 -289.175 -82.265 ;
        RECT -288.990 -82.520 -288.715 -82.255 ;
        RECT -279.530 -82.530 -279.255 -82.265 ;
        RECT -279.070 -82.520 -278.795 -82.255 ;
        RECT -269.610 -82.530 -269.335 -82.265 ;
        RECT -269.150 -82.520 -268.875 -82.255 ;
        RECT -259.690 -82.530 -259.415 -82.265 ;
        RECT -259.230 -82.520 -258.955 -82.255 ;
        RECT -249.770 -82.530 -249.495 -82.265 ;
        RECT -249.310 -82.520 -249.035 -82.255 ;
        RECT -239.850 -82.530 -239.575 -82.265 ;
        RECT -239.390 -82.520 -239.115 -82.255 ;
        RECT -229.930 -82.530 -229.655 -82.265 ;
        RECT -229.470 -82.520 -229.195 -82.255 ;
        RECT -220.010 -82.530 -219.735 -82.265 ;
        RECT -219.550 -82.520 -219.275 -82.255 ;
        RECT -210.090 -82.530 -209.815 -82.265 ;
        RECT -209.630 -82.520 -209.355 -82.255 ;
        RECT -200.170 -82.530 -199.895 -82.265 ;
        RECT -199.710 -82.520 -199.435 -82.255 ;
        RECT -190.250 -82.530 -189.975 -82.265 ;
        RECT -189.790 -82.520 -189.515 -82.255 ;
        RECT -180.330 -82.530 -180.055 -82.265 ;
        RECT -179.870 -82.520 -179.595 -82.255 ;
        RECT -170.410 -82.530 -170.135 -82.265 ;
        RECT -169.950 -82.520 -169.675 -82.255 ;
        RECT -160.490 -82.530 -160.215 -82.265 ;
        RECT -160.030 -82.520 -159.755 -82.255 ;
        RECT -150.570 -82.530 -150.295 -82.265 ;
        RECT -150.110 -82.520 -149.835 -82.255 ;
        RECT -140.650 -82.530 -140.375 -82.265 ;
        RECT -140.190 -82.520 -139.915 -82.255 ;
        RECT -130.730 -82.530 -130.455 -82.265 ;
        RECT -130.270 -82.520 -129.995 -82.255 ;
        RECT -120.810 -82.530 -120.535 -82.265 ;
        RECT -120.350 -82.520 -120.075 -82.255 ;
        RECT -110.890 -82.530 -110.615 -82.265 ;
        RECT -110.430 -82.520 -110.155 -82.255 ;
        RECT -100.970 -82.530 -100.695 -82.265 ;
        RECT -100.510 -82.520 -100.235 -82.255 ;
        RECT -91.050 -82.530 -90.775 -82.265 ;
        RECT -90.590 -82.520 -90.315 -82.255 ;
        RECT -81.130 -82.530 -80.855 -82.265 ;
        RECT -80.670 -82.520 -80.395 -82.255 ;
        RECT -71.210 -82.530 -70.935 -82.265 ;
        RECT -70.750 -82.520 -70.475 -82.255 ;
        RECT -61.290 -82.530 -61.015 -82.265 ;
        RECT -60.830 -82.520 -60.555 -82.255 ;
        RECT -51.370 -82.530 -51.095 -82.265 ;
        RECT -50.910 -82.520 -50.635 -82.255 ;
        RECT -41.450 -82.530 -41.175 -82.265 ;
        RECT -40.990 -82.520 -40.715 -82.255 ;
        RECT -31.530 -82.530 -31.255 -82.265 ;
        RECT -31.070 -82.520 -30.795 -82.255 ;
        RECT -21.610 -82.530 -21.335 -82.265 ;
        RECT -21.150 -82.520 -20.875 -82.255 ;
        RECT -11.690 -82.530 -11.415 -82.265 ;
        RECT -11.230 -82.520 -10.955 -82.255 ;
        RECT -1.770 -82.530 -1.495 -82.265 ;
        RECT -1.310 -82.520 -1.035 -82.255 ;
        RECT 8.150 -82.530 8.425 -82.265 ;
        RECT 8.610 -82.520 8.885 -82.255 ;
        RECT 18.070 -82.530 18.345 -82.265 ;
        RECT 18.530 -82.520 18.805 -82.255 ;
        RECT -281.800 -83.290 -281.525 -83.025 ;
        RECT -271.880 -83.290 -271.605 -83.025 ;
        RECT -261.960 -83.290 -261.685 -83.025 ;
        RECT -252.040 -83.290 -251.765 -83.025 ;
        RECT -242.120 -83.290 -241.845 -83.025 ;
        RECT -232.200 -83.290 -231.925 -83.025 ;
        RECT -222.280 -83.290 -222.005 -83.025 ;
        RECT -212.360 -83.290 -212.085 -83.025 ;
        RECT -202.440 -83.290 -202.165 -83.025 ;
        RECT -192.520 -83.290 -192.245 -83.025 ;
        RECT -182.600 -83.290 -182.325 -83.025 ;
        RECT -172.680 -83.290 -172.405 -83.025 ;
        RECT -162.760 -83.290 -162.485 -83.025 ;
        RECT -152.840 -83.290 -152.565 -83.025 ;
        RECT -142.920 -83.290 -142.645 -83.025 ;
        RECT -133.000 -83.290 -132.725 -83.025 ;
        RECT -123.080 -83.290 -122.805 -83.025 ;
        RECT -113.160 -83.290 -112.885 -83.025 ;
        RECT -103.240 -83.290 -102.965 -83.025 ;
        RECT -93.320 -83.290 -93.045 -83.025 ;
        RECT -83.400 -83.290 -83.125 -83.025 ;
        RECT -73.480 -83.290 -73.205 -83.025 ;
        RECT -63.560 -83.290 -63.285 -83.025 ;
        RECT -53.640 -83.290 -53.365 -83.025 ;
        RECT -43.720 -83.290 -43.445 -83.025 ;
        RECT -33.800 -83.290 -33.525 -83.025 ;
        RECT -23.880 -83.290 -23.605 -83.025 ;
        RECT -13.960 -83.290 -13.685 -83.025 ;
        RECT -4.040 -83.290 -3.765 -83.025 ;
        RECT 5.880 -83.290 6.155 -83.025 ;
        RECT 15.800 -83.290 16.075 -83.025 ;
        RECT -291.120 -173.510 -290.845 -173.245 ;
        RECT -281.200 -173.510 -280.925 -173.245 ;
        RECT -271.280 -173.510 -271.005 -173.245 ;
        RECT -261.360 -173.510 -261.085 -173.245 ;
        RECT -251.440 -173.510 -251.165 -173.245 ;
        RECT -241.520 -173.510 -241.245 -173.245 ;
        RECT -231.600 -173.510 -231.325 -173.245 ;
        RECT -221.680 -173.510 -221.405 -173.245 ;
        RECT -211.760 -173.510 -211.485 -173.245 ;
        RECT -201.840 -173.510 -201.565 -173.245 ;
        RECT -191.920 -173.510 -191.645 -173.245 ;
        RECT -182.000 -173.510 -181.725 -173.245 ;
        RECT -172.080 -173.510 -171.805 -173.245 ;
        RECT -162.160 -173.510 -161.885 -173.245 ;
        RECT -152.240 -173.510 -151.965 -173.245 ;
        RECT -142.320 -173.510 -142.045 -173.245 ;
        RECT -132.400 -173.510 -132.125 -173.245 ;
        RECT -122.480 -173.510 -122.205 -173.245 ;
        RECT -112.560 -173.510 -112.285 -173.245 ;
        RECT -102.640 -173.510 -102.365 -173.245 ;
        RECT -92.720 -173.510 -92.445 -173.245 ;
        RECT -82.800 -173.510 -82.525 -173.245 ;
        RECT -72.880 -173.510 -72.605 -173.245 ;
        RECT -62.960 -173.510 -62.685 -173.245 ;
        RECT -53.040 -173.510 -52.765 -173.245 ;
        RECT -43.120 -173.510 -42.845 -173.245 ;
        RECT -33.200 -173.510 -32.925 -173.245 ;
        RECT -23.280 -173.510 -23.005 -173.245 ;
        RECT -13.360 -173.510 -13.085 -173.245 ;
        RECT -3.440 -173.510 -3.165 -173.245 ;
        RECT 6.480 -173.510 6.755 -173.245 ;
        RECT 16.400 -173.510 16.675 -173.245 ;
        RECT -283.950 -174.380 -283.675 -174.115 ;
        RECT -283.480 -174.380 -283.205 -174.115 ;
        RECT -274.030 -174.380 -273.755 -174.115 ;
        RECT -273.560 -174.380 -273.285 -174.115 ;
        RECT -264.110 -174.380 -263.835 -174.115 ;
        RECT -263.640 -174.380 -263.365 -174.115 ;
        RECT -254.190 -174.380 -253.915 -174.115 ;
        RECT -253.720 -174.380 -253.445 -174.115 ;
        RECT -244.270 -174.380 -243.995 -174.115 ;
        RECT -243.800 -174.380 -243.525 -174.115 ;
        RECT -234.350 -174.380 -234.075 -174.115 ;
        RECT -233.880 -174.380 -233.605 -174.115 ;
        RECT -224.430 -174.380 -224.155 -174.115 ;
        RECT -223.960 -174.380 -223.685 -174.115 ;
        RECT -214.510 -174.380 -214.235 -174.115 ;
        RECT -214.040 -174.380 -213.765 -174.115 ;
        RECT -204.590 -174.380 -204.315 -174.115 ;
        RECT -204.120 -174.380 -203.845 -174.115 ;
        RECT -194.670 -174.380 -194.395 -174.115 ;
        RECT -194.200 -174.380 -193.925 -174.115 ;
        RECT -184.750 -174.380 -184.475 -174.115 ;
        RECT -184.280 -174.380 -184.005 -174.115 ;
        RECT -174.830 -174.380 -174.555 -174.115 ;
        RECT -174.360 -174.380 -174.085 -174.115 ;
        RECT -164.910 -174.380 -164.635 -174.115 ;
        RECT -164.440 -174.380 -164.165 -174.115 ;
        RECT -154.990 -174.380 -154.715 -174.115 ;
        RECT -154.520 -174.380 -154.245 -174.115 ;
        RECT -145.070 -174.380 -144.795 -174.115 ;
        RECT -144.600 -174.380 -144.325 -174.115 ;
        RECT -135.150 -174.380 -134.875 -174.115 ;
        RECT -134.680 -174.380 -134.405 -174.115 ;
        RECT -125.230 -174.380 -124.955 -174.115 ;
        RECT -124.760 -174.380 -124.485 -174.115 ;
        RECT -115.310 -174.380 -115.035 -174.115 ;
        RECT -114.840 -174.380 -114.565 -174.115 ;
        RECT -105.390 -174.380 -105.115 -174.115 ;
        RECT -104.920 -174.380 -104.645 -174.115 ;
        RECT -95.470 -174.380 -95.195 -174.115 ;
        RECT -95.000 -174.380 -94.725 -174.115 ;
        RECT -85.550 -174.380 -85.275 -174.115 ;
        RECT -85.080 -174.380 -84.805 -174.115 ;
        RECT -75.630 -174.380 -75.355 -174.115 ;
        RECT -75.160 -174.380 -74.885 -174.115 ;
        RECT -65.710 -174.380 -65.435 -174.115 ;
        RECT -65.240 -174.380 -64.965 -174.115 ;
        RECT -55.790 -174.380 -55.515 -174.115 ;
        RECT -55.320 -174.380 -55.045 -174.115 ;
        RECT -45.870 -174.380 -45.595 -174.115 ;
        RECT -45.400 -174.380 -45.125 -174.115 ;
        RECT -35.950 -174.380 -35.675 -174.115 ;
        RECT -35.480 -174.380 -35.205 -174.115 ;
        RECT -26.030 -174.380 -25.755 -174.115 ;
        RECT -25.560 -174.380 -25.285 -174.115 ;
        RECT -16.110 -174.380 -15.835 -174.115 ;
        RECT -15.640 -174.380 -15.365 -174.115 ;
        RECT -6.190 -174.380 -5.915 -174.115 ;
        RECT -5.720 -174.380 -5.445 -174.115 ;
        RECT 3.730 -174.380 4.005 -174.115 ;
        RECT 4.200 -174.380 4.475 -174.115 ;
        RECT 13.650 -174.380 13.925 -174.115 ;
        RECT 14.120 -174.380 14.395 -174.115 ;
        RECT -291.210 -177.110 -290.935 -176.845 ;
        RECT -290.750 -177.100 -290.475 -176.835 ;
        RECT -281.290 -177.110 -281.015 -176.845 ;
        RECT -280.830 -177.100 -280.555 -176.835 ;
        RECT -271.370 -177.110 -271.095 -176.845 ;
        RECT -270.910 -177.100 -270.635 -176.835 ;
        RECT -261.450 -177.110 -261.175 -176.845 ;
        RECT -260.990 -177.100 -260.715 -176.835 ;
        RECT -251.530 -177.110 -251.255 -176.845 ;
        RECT -251.070 -177.100 -250.795 -176.835 ;
        RECT -241.610 -177.110 -241.335 -176.845 ;
        RECT -241.150 -177.100 -240.875 -176.835 ;
        RECT -231.690 -177.110 -231.415 -176.845 ;
        RECT -231.230 -177.100 -230.955 -176.835 ;
        RECT -221.770 -177.110 -221.495 -176.845 ;
        RECT -221.310 -177.100 -221.035 -176.835 ;
        RECT -211.850 -177.110 -211.575 -176.845 ;
        RECT -211.390 -177.100 -211.115 -176.835 ;
        RECT -201.930 -177.110 -201.655 -176.845 ;
        RECT -201.470 -177.100 -201.195 -176.835 ;
        RECT -192.010 -177.110 -191.735 -176.845 ;
        RECT -191.550 -177.100 -191.275 -176.835 ;
        RECT -182.090 -177.110 -181.815 -176.845 ;
        RECT -181.630 -177.100 -181.355 -176.835 ;
        RECT -172.170 -177.110 -171.895 -176.845 ;
        RECT -171.710 -177.100 -171.435 -176.835 ;
        RECT -162.250 -177.110 -161.975 -176.845 ;
        RECT -161.790 -177.100 -161.515 -176.835 ;
        RECT -152.330 -177.110 -152.055 -176.845 ;
        RECT -151.870 -177.100 -151.595 -176.835 ;
        RECT -142.410 -177.110 -142.135 -176.845 ;
        RECT -141.950 -177.100 -141.675 -176.835 ;
        RECT -132.490 -177.110 -132.215 -176.845 ;
        RECT -132.030 -177.100 -131.755 -176.835 ;
        RECT -122.570 -177.110 -122.295 -176.845 ;
        RECT -122.110 -177.100 -121.835 -176.835 ;
        RECT -112.650 -177.110 -112.375 -176.845 ;
        RECT -112.190 -177.100 -111.915 -176.835 ;
        RECT -102.730 -177.110 -102.455 -176.845 ;
        RECT -102.270 -177.100 -101.995 -176.835 ;
        RECT -92.810 -177.110 -92.535 -176.845 ;
        RECT -92.350 -177.100 -92.075 -176.835 ;
        RECT -82.890 -177.110 -82.615 -176.845 ;
        RECT -82.430 -177.100 -82.155 -176.835 ;
        RECT -72.970 -177.110 -72.695 -176.845 ;
        RECT -72.510 -177.100 -72.235 -176.835 ;
        RECT -63.050 -177.110 -62.775 -176.845 ;
        RECT -62.590 -177.100 -62.315 -176.835 ;
        RECT -53.130 -177.110 -52.855 -176.845 ;
        RECT -52.670 -177.100 -52.395 -176.835 ;
        RECT -43.210 -177.110 -42.935 -176.845 ;
        RECT -42.750 -177.100 -42.475 -176.835 ;
        RECT -33.290 -177.110 -33.015 -176.845 ;
        RECT -32.830 -177.100 -32.555 -176.835 ;
        RECT -23.370 -177.110 -23.095 -176.845 ;
        RECT -22.910 -177.100 -22.635 -176.835 ;
        RECT -13.450 -177.110 -13.175 -176.845 ;
        RECT -12.990 -177.100 -12.715 -176.835 ;
        RECT -3.530 -177.110 -3.255 -176.845 ;
        RECT -3.070 -177.100 -2.795 -176.835 ;
        RECT 6.390 -177.110 6.665 -176.845 ;
        RECT 6.850 -177.100 7.125 -176.835 ;
        RECT 16.310 -177.110 16.585 -176.845 ;
        RECT 16.770 -177.100 17.045 -176.835 ;
        RECT -283.560 -177.870 -283.285 -177.605 ;
        RECT -273.640 -177.870 -273.365 -177.605 ;
        RECT -263.720 -177.870 -263.445 -177.605 ;
        RECT -253.800 -177.870 -253.525 -177.605 ;
        RECT -243.880 -177.870 -243.605 -177.605 ;
        RECT -233.960 -177.870 -233.685 -177.605 ;
        RECT -224.040 -177.870 -223.765 -177.605 ;
        RECT -214.120 -177.870 -213.845 -177.605 ;
        RECT -204.200 -177.870 -203.925 -177.605 ;
        RECT -194.280 -177.870 -194.005 -177.605 ;
        RECT -184.360 -177.870 -184.085 -177.605 ;
        RECT -174.440 -177.870 -174.165 -177.605 ;
        RECT -164.520 -177.870 -164.245 -177.605 ;
        RECT -154.600 -177.870 -154.325 -177.605 ;
        RECT -144.680 -177.870 -144.405 -177.605 ;
        RECT -134.760 -177.870 -134.485 -177.605 ;
        RECT -124.840 -177.870 -124.565 -177.605 ;
        RECT -114.920 -177.870 -114.645 -177.605 ;
        RECT -105.000 -177.870 -104.725 -177.605 ;
        RECT -95.080 -177.870 -94.805 -177.605 ;
        RECT -85.160 -177.870 -84.885 -177.605 ;
        RECT -75.240 -177.870 -74.965 -177.605 ;
        RECT -65.320 -177.870 -65.045 -177.605 ;
        RECT -55.400 -177.870 -55.125 -177.605 ;
        RECT -45.480 -177.870 -45.205 -177.605 ;
        RECT -35.560 -177.870 -35.285 -177.605 ;
        RECT -25.640 -177.870 -25.365 -177.605 ;
        RECT -15.720 -177.870 -15.445 -177.605 ;
        RECT -5.800 -177.870 -5.525 -177.605 ;
        RECT 4.120 -177.870 4.395 -177.605 ;
        RECT 14.040 -177.870 14.315 -177.605 ;
      LAYER met2 ;
        RECT -288.280 93.760 -287.110 94.560 ;
        RECT -278.360 93.760 -277.190 94.560 ;
        RECT -268.440 93.760 -267.270 94.560 ;
        RECT -258.520 93.760 -257.350 94.560 ;
        RECT -248.600 93.760 -247.430 94.560 ;
        RECT -238.680 93.760 -237.510 94.560 ;
        RECT -228.760 93.760 -227.590 94.560 ;
        RECT -218.840 93.760 -217.670 94.560 ;
        RECT -208.920 93.760 -207.750 94.560 ;
        RECT -199.000 93.760 -197.830 94.560 ;
        RECT -189.080 93.760 -187.910 94.560 ;
        RECT -179.160 93.760 -177.990 94.560 ;
        RECT -169.240 93.760 -168.070 94.560 ;
        RECT -159.320 93.760 -158.150 94.560 ;
        RECT -149.400 93.760 -148.230 94.560 ;
        RECT -139.480 93.760 -138.310 94.560 ;
        RECT -129.560 93.760 -128.390 94.560 ;
        RECT -119.640 93.760 -118.470 94.560 ;
        RECT -109.720 93.760 -108.550 94.560 ;
        RECT -99.800 93.760 -98.630 94.560 ;
        RECT -89.880 93.760 -88.710 94.560 ;
        RECT -79.960 93.760 -78.790 94.560 ;
        RECT -70.040 93.760 -68.870 94.560 ;
        RECT -60.120 93.760 -58.950 94.560 ;
        RECT -50.200 93.760 -49.030 94.560 ;
        RECT -40.280 93.760 -39.110 94.560 ;
        RECT -30.360 93.760 -29.190 94.560 ;
        RECT -20.440 93.760 -19.270 94.560 ;
        RECT -10.520 93.760 -9.350 94.560 ;
        RECT -0.600 93.760 0.570 94.560 ;
        RECT 9.320 93.760 10.490 94.560 ;
        RECT 19.240 93.760 20.410 94.560 ;
        RECT -280.620 93.090 -279.700 93.570 ;
        RECT -270.700 93.090 -269.780 93.570 ;
        RECT -260.780 93.090 -259.860 93.570 ;
        RECT -250.860 93.090 -249.940 93.570 ;
        RECT -240.940 93.090 -240.020 93.570 ;
        RECT -231.020 93.090 -230.100 93.570 ;
        RECT -221.100 93.090 -220.180 93.570 ;
        RECT -211.180 93.090 -210.260 93.570 ;
        RECT -201.260 93.090 -200.340 93.570 ;
        RECT -191.340 93.090 -190.420 93.570 ;
        RECT -181.420 93.090 -180.500 93.570 ;
        RECT -171.500 93.090 -170.580 93.570 ;
        RECT -161.580 93.090 -160.660 93.570 ;
        RECT -151.660 93.090 -150.740 93.570 ;
        RECT -141.740 93.090 -140.820 93.570 ;
        RECT -131.820 93.090 -130.900 93.570 ;
        RECT -121.900 93.090 -120.980 93.570 ;
        RECT -111.980 93.090 -111.060 93.570 ;
        RECT -102.060 93.090 -101.140 93.570 ;
        RECT -92.140 93.090 -91.220 93.570 ;
        RECT -82.220 93.090 -81.300 93.570 ;
        RECT -72.300 93.090 -71.380 93.570 ;
        RECT -62.380 93.090 -61.460 93.570 ;
        RECT -52.460 93.090 -51.540 93.570 ;
        RECT -42.540 93.090 -41.620 93.570 ;
        RECT -32.620 93.090 -31.700 93.570 ;
        RECT -22.700 93.090 -21.780 93.570 ;
        RECT -12.780 93.090 -11.860 93.570 ;
        RECT -2.860 93.090 -1.940 93.570 ;
        RECT 7.060 93.090 7.980 93.570 ;
        RECT 16.980 93.090 17.900 93.570 ;
        RECT -287.880 90.370 -286.960 90.850 ;
        RECT -277.960 90.370 -277.040 90.850 ;
        RECT -268.040 90.370 -267.120 90.850 ;
        RECT -258.120 90.370 -257.200 90.850 ;
        RECT -248.200 90.370 -247.280 90.850 ;
        RECT -238.280 90.370 -237.360 90.850 ;
        RECT -228.360 90.370 -227.440 90.850 ;
        RECT -218.440 90.370 -217.520 90.850 ;
        RECT -208.520 90.370 -207.600 90.850 ;
        RECT -198.600 90.370 -197.680 90.850 ;
        RECT -188.680 90.370 -187.760 90.850 ;
        RECT -178.760 90.370 -177.840 90.850 ;
        RECT -168.840 90.370 -167.920 90.850 ;
        RECT -158.920 90.370 -158.000 90.850 ;
        RECT -149.000 90.370 -148.080 90.850 ;
        RECT -139.080 90.370 -138.160 90.850 ;
        RECT -129.160 90.370 -128.240 90.850 ;
        RECT -119.240 90.370 -118.320 90.850 ;
        RECT -109.320 90.370 -108.400 90.850 ;
        RECT -99.400 90.370 -98.480 90.850 ;
        RECT -89.480 90.370 -88.560 90.850 ;
        RECT -79.560 90.370 -78.640 90.850 ;
        RECT -69.640 90.370 -68.720 90.850 ;
        RECT -59.720 90.370 -58.800 90.850 ;
        RECT -49.800 90.370 -48.880 90.850 ;
        RECT -39.880 90.370 -38.960 90.850 ;
        RECT -29.960 90.370 -29.040 90.850 ;
        RECT -20.040 90.370 -19.120 90.850 ;
        RECT -10.120 90.370 -9.200 90.850 ;
        RECT -0.200 90.370 0.720 90.850 ;
        RECT 9.720 90.370 10.640 90.850 ;
        RECT 19.640 90.370 20.560 90.850 ;
        RECT -280.460 89.390 -279.290 90.190 ;
        RECT -270.540 89.390 -269.370 90.190 ;
        RECT -260.620 89.390 -259.450 90.190 ;
        RECT -250.700 89.390 -249.530 90.190 ;
        RECT -240.780 89.390 -239.610 90.190 ;
        RECT -230.860 89.390 -229.690 90.190 ;
        RECT -220.940 89.390 -219.770 90.190 ;
        RECT -211.020 89.390 -209.850 90.190 ;
        RECT -201.100 89.390 -199.930 90.190 ;
        RECT -191.180 89.390 -190.010 90.190 ;
        RECT -181.260 89.390 -180.090 90.190 ;
        RECT -171.340 89.390 -170.170 90.190 ;
        RECT -161.420 89.390 -160.250 90.190 ;
        RECT -151.500 89.390 -150.330 90.190 ;
        RECT -141.580 89.390 -140.410 90.190 ;
        RECT -131.660 89.390 -130.490 90.190 ;
        RECT -121.740 89.390 -120.570 90.190 ;
        RECT -111.820 89.390 -110.650 90.190 ;
        RECT -101.900 89.390 -100.730 90.190 ;
        RECT -91.980 89.390 -90.810 90.190 ;
        RECT -82.060 89.390 -80.890 90.190 ;
        RECT -72.140 89.390 -70.970 90.190 ;
        RECT -62.220 89.390 -61.050 90.190 ;
        RECT -52.300 89.390 -51.130 90.190 ;
        RECT -42.380 89.390 -41.210 90.190 ;
        RECT -32.460 89.390 -31.290 90.190 ;
        RECT -22.540 89.390 -21.370 90.190 ;
        RECT -12.620 89.390 -11.450 90.190 ;
        RECT -2.700 89.390 -1.530 90.190 ;
        RECT 7.220 89.390 8.390 90.190 ;
        RECT 17.140 89.390 18.310 90.190 ;
        RECT -290.300 9.710 -289.130 10.510 ;
        RECT -280.380 9.710 -279.210 10.510 ;
        RECT -270.460 9.710 -269.290 10.510 ;
        RECT -260.540 9.710 -259.370 10.510 ;
        RECT -250.620 9.710 -249.450 10.510 ;
        RECT -240.700 9.710 -239.530 10.510 ;
        RECT -230.780 9.710 -229.610 10.510 ;
        RECT -220.860 9.710 -219.690 10.510 ;
        RECT -210.940 9.710 -209.770 10.510 ;
        RECT -201.020 9.710 -199.850 10.510 ;
        RECT -191.100 9.710 -189.930 10.510 ;
        RECT -181.180 9.710 -180.010 10.510 ;
        RECT -171.260 9.710 -170.090 10.510 ;
        RECT -161.340 9.710 -160.170 10.510 ;
        RECT -151.420 9.710 -150.250 10.510 ;
        RECT -141.500 9.710 -140.330 10.510 ;
        RECT -131.580 9.710 -130.410 10.510 ;
        RECT -121.660 9.710 -120.490 10.510 ;
        RECT -111.740 9.710 -110.570 10.510 ;
        RECT -101.820 9.710 -100.650 10.510 ;
        RECT -91.900 9.710 -90.730 10.510 ;
        RECT -81.980 9.710 -80.810 10.510 ;
        RECT -72.060 9.710 -70.890 10.510 ;
        RECT -62.140 9.710 -60.970 10.510 ;
        RECT -52.220 9.710 -51.050 10.510 ;
        RECT -42.300 9.710 -41.130 10.510 ;
        RECT -32.380 9.710 -31.210 10.510 ;
        RECT -22.460 9.710 -21.290 10.510 ;
        RECT -12.540 9.710 -11.370 10.510 ;
        RECT -2.620 9.710 -1.450 10.510 ;
        RECT 7.300 9.710 8.470 10.510 ;
        RECT 17.220 9.710 18.390 10.510 ;
        RECT -282.640 9.040 -281.720 9.520 ;
        RECT -272.720 9.040 -271.800 9.520 ;
        RECT -262.800 9.040 -261.880 9.520 ;
        RECT -252.880 9.040 -251.960 9.520 ;
        RECT -242.960 9.040 -242.040 9.520 ;
        RECT -233.040 9.040 -232.120 9.520 ;
        RECT -223.120 9.040 -222.200 9.520 ;
        RECT -213.200 9.040 -212.280 9.520 ;
        RECT -203.280 9.040 -202.360 9.520 ;
        RECT -193.360 9.040 -192.440 9.520 ;
        RECT -183.440 9.040 -182.520 9.520 ;
        RECT -173.520 9.040 -172.600 9.520 ;
        RECT -163.600 9.040 -162.680 9.520 ;
        RECT -153.680 9.040 -152.760 9.520 ;
        RECT -143.760 9.040 -142.840 9.520 ;
        RECT -133.840 9.040 -132.920 9.520 ;
        RECT -123.920 9.040 -123.000 9.520 ;
        RECT -114.000 9.040 -113.080 9.520 ;
        RECT -104.080 9.040 -103.160 9.520 ;
        RECT -94.160 9.040 -93.240 9.520 ;
        RECT -84.240 9.040 -83.320 9.520 ;
        RECT -74.320 9.040 -73.400 9.520 ;
        RECT -64.400 9.040 -63.480 9.520 ;
        RECT -54.480 9.040 -53.560 9.520 ;
        RECT -44.560 9.040 -43.640 9.520 ;
        RECT -34.640 9.040 -33.720 9.520 ;
        RECT -24.720 9.040 -23.800 9.520 ;
        RECT -14.800 9.040 -13.880 9.520 ;
        RECT -4.880 9.040 -3.960 9.520 ;
        RECT 5.040 9.040 5.960 9.520 ;
        RECT 14.960 9.040 15.880 9.520 ;
        RECT -289.900 6.320 -288.980 6.800 ;
        RECT -279.980 6.320 -279.060 6.800 ;
        RECT -270.060 6.320 -269.140 6.800 ;
        RECT -260.140 6.320 -259.220 6.800 ;
        RECT -250.220 6.320 -249.300 6.800 ;
        RECT -240.300 6.320 -239.380 6.800 ;
        RECT -230.380 6.320 -229.460 6.800 ;
        RECT -220.460 6.320 -219.540 6.800 ;
        RECT -210.540 6.320 -209.620 6.800 ;
        RECT -200.620 6.320 -199.700 6.800 ;
        RECT -190.700 6.320 -189.780 6.800 ;
        RECT -180.780 6.320 -179.860 6.800 ;
        RECT -170.860 6.320 -169.940 6.800 ;
        RECT -160.940 6.320 -160.020 6.800 ;
        RECT -151.020 6.320 -150.100 6.800 ;
        RECT -141.100 6.320 -140.180 6.800 ;
        RECT -131.180 6.320 -130.260 6.800 ;
        RECT -121.260 6.320 -120.340 6.800 ;
        RECT -111.340 6.320 -110.420 6.800 ;
        RECT -101.420 6.320 -100.500 6.800 ;
        RECT -91.500 6.320 -90.580 6.800 ;
        RECT -81.580 6.320 -80.660 6.800 ;
        RECT -71.660 6.320 -70.740 6.800 ;
        RECT -61.740 6.320 -60.820 6.800 ;
        RECT -51.820 6.320 -50.900 6.800 ;
        RECT -41.900 6.320 -40.980 6.800 ;
        RECT -31.980 6.320 -31.060 6.800 ;
        RECT -22.060 6.320 -21.140 6.800 ;
        RECT -12.140 6.320 -11.220 6.800 ;
        RECT -2.220 6.320 -1.300 6.800 ;
        RECT 7.700 6.320 8.620 6.800 ;
        RECT 17.620 6.320 18.540 6.800 ;
        RECT -282.480 5.340 -281.310 6.140 ;
        RECT -272.560 5.340 -271.390 6.140 ;
        RECT -262.640 5.340 -261.470 6.140 ;
        RECT -252.720 5.340 -251.550 6.140 ;
        RECT -242.800 5.340 -241.630 6.140 ;
        RECT -232.880 5.340 -231.710 6.140 ;
        RECT -222.960 5.340 -221.790 6.140 ;
        RECT -213.040 5.340 -211.870 6.140 ;
        RECT -203.120 5.340 -201.950 6.140 ;
        RECT -193.200 5.340 -192.030 6.140 ;
        RECT -183.280 5.340 -182.110 6.140 ;
        RECT -173.360 5.340 -172.190 6.140 ;
        RECT -163.440 5.340 -162.270 6.140 ;
        RECT -153.520 5.340 -152.350 6.140 ;
        RECT -143.600 5.340 -142.430 6.140 ;
        RECT -133.680 5.340 -132.510 6.140 ;
        RECT -123.760 5.340 -122.590 6.140 ;
        RECT -113.840 5.340 -112.670 6.140 ;
        RECT -103.920 5.340 -102.750 6.140 ;
        RECT -94.000 5.340 -92.830 6.140 ;
        RECT -84.080 5.340 -82.910 6.140 ;
        RECT -74.160 5.340 -72.990 6.140 ;
        RECT -64.240 5.340 -63.070 6.140 ;
        RECT -54.320 5.340 -53.150 6.140 ;
        RECT -44.400 5.340 -43.230 6.140 ;
        RECT -34.480 5.340 -33.310 6.140 ;
        RECT -24.560 5.340 -23.390 6.140 ;
        RECT -14.640 5.340 -13.470 6.140 ;
        RECT -4.720 5.340 -3.550 6.140 ;
        RECT 5.200 5.340 6.370 6.140 ;
        RECT 15.120 5.340 16.290 6.140 ;
        RECT -289.940 -79.240 -288.770 -78.440 ;
        RECT -280.020 -79.240 -278.850 -78.440 ;
        RECT -270.100 -79.240 -268.930 -78.440 ;
        RECT -260.180 -79.240 -259.010 -78.440 ;
        RECT -250.260 -79.240 -249.090 -78.440 ;
        RECT -240.340 -79.240 -239.170 -78.440 ;
        RECT -230.420 -79.240 -229.250 -78.440 ;
        RECT -220.500 -79.240 -219.330 -78.440 ;
        RECT -210.580 -79.240 -209.410 -78.440 ;
        RECT -200.660 -79.240 -199.490 -78.440 ;
        RECT -190.740 -79.240 -189.570 -78.440 ;
        RECT -180.820 -79.240 -179.650 -78.440 ;
        RECT -170.900 -79.240 -169.730 -78.440 ;
        RECT -160.980 -79.240 -159.810 -78.440 ;
        RECT -151.060 -79.240 -149.890 -78.440 ;
        RECT -141.140 -79.240 -139.970 -78.440 ;
        RECT -131.220 -79.240 -130.050 -78.440 ;
        RECT -121.300 -79.240 -120.130 -78.440 ;
        RECT -111.380 -79.240 -110.210 -78.440 ;
        RECT -101.460 -79.240 -100.290 -78.440 ;
        RECT -91.540 -79.240 -90.370 -78.440 ;
        RECT -81.620 -79.240 -80.450 -78.440 ;
        RECT -71.700 -79.240 -70.530 -78.440 ;
        RECT -61.780 -79.240 -60.610 -78.440 ;
        RECT -51.860 -79.240 -50.690 -78.440 ;
        RECT -41.940 -79.240 -40.770 -78.440 ;
        RECT -32.020 -79.240 -30.850 -78.440 ;
        RECT -22.100 -79.240 -20.930 -78.440 ;
        RECT -12.180 -79.240 -11.010 -78.440 ;
        RECT -2.260 -79.240 -1.090 -78.440 ;
        RECT 7.660 -79.240 8.830 -78.440 ;
        RECT 17.580 -79.240 18.750 -78.440 ;
        RECT -282.280 -79.910 -281.360 -79.430 ;
        RECT -272.360 -79.910 -271.440 -79.430 ;
        RECT -262.440 -79.910 -261.520 -79.430 ;
        RECT -252.520 -79.910 -251.600 -79.430 ;
        RECT -242.600 -79.910 -241.680 -79.430 ;
        RECT -232.680 -79.910 -231.760 -79.430 ;
        RECT -222.760 -79.910 -221.840 -79.430 ;
        RECT -212.840 -79.910 -211.920 -79.430 ;
        RECT -202.920 -79.910 -202.000 -79.430 ;
        RECT -193.000 -79.910 -192.080 -79.430 ;
        RECT -183.080 -79.910 -182.160 -79.430 ;
        RECT -173.160 -79.910 -172.240 -79.430 ;
        RECT -163.240 -79.910 -162.320 -79.430 ;
        RECT -153.320 -79.910 -152.400 -79.430 ;
        RECT -143.400 -79.910 -142.480 -79.430 ;
        RECT -133.480 -79.910 -132.560 -79.430 ;
        RECT -123.560 -79.910 -122.640 -79.430 ;
        RECT -113.640 -79.910 -112.720 -79.430 ;
        RECT -103.720 -79.910 -102.800 -79.430 ;
        RECT -93.800 -79.910 -92.880 -79.430 ;
        RECT -83.880 -79.910 -82.960 -79.430 ;
        RECT -73.960 -79.910 -73.040 -79.430 ;
        RECT -64.040 -79.910 -63.120 -79.430 ;
        RECT -54.120 -79.910 -53.200 -79.430 ;
        RECT -44.200 -79.910 -43.280 -79.430 ;
        RECT -34.280 -79.910 -33.360 -79.430 ;
        RECT -24.360 -79.910 -23.440 -79.430 ;
        RECT -14.440 -79.910 -13.520 -79.430 ;
        RECT -4.520 -79.910 -3.600 -79.430 ;
        RECT 5.400 -79.910 6.320 -79.430 ;
        RECT 15.320 -79.910 16.240 -79.430 ;
        RECT -289.540 -82.630 -288.620 -82.150 ;
        RECT -279.620 -82.630 -278.700 -82.150 ;
        RECT -269.700 -82.630 -268.780 -82.150 ;
        RECT -259.780 -82.630 -258.860 -82.150 ;
        RECT -249.860 -82.630 -248.940 -82.150 ;
        RECT -239.940 -82.630 -239.020 -82.150 ;
        RECT -230.020 -82.630 -229.100 -82.150 ;
        RECT -220.100 -82.630 -219.180 -82.150 ;
        RECT -210.180 -82.630 -209.260 -82.150 ;
        RECT -200.260 -82.630 -199.340 -82.150 ;
        RECT -190.340 -82.630 -189.420 -82.150 ;
        RECT -180.420 -82.630 -179.500 -82.150 ;
        RECT -170.500 -82.630 -169.580 -82.150 ;
        RECT -160.580 -82.630 -159.660 -82.150 ;
        RECT -150.660 -82.630 -149.740 -82.150 ;
        RECT -140.740 -82.630 -139.820 -82.150 ;
        RECT -130.820 -82.630 -129.900 -82.150 ;
        RECT -120.900 -82.630 -119.980 -82.150 ;
        RECT -110.980 -82.630 -110.060 -82.150 ;
        RECT -101.060 -82.630 -100.140 -82.150 ;
        RECT -91.140 -82.630 -90.220 -82.150 ;
        RECT -81.220 -82.630 -80.300 -82.150 ;
        RECT -71.300 -82.630 -70.380 -82.150 ;
        RECT -61.380 -82.630 -60.460 -82.150 ;
        RECT -51.460 -82.630 -50.540 -82.150 ;
        RECT -41.540 -82.630 -40.620 -82.150 ;
        RECT -31.620 -82.630 -30.700 -82.150 ;
        RECT -21.700 -82.630 -20.780 -82.150 ;
        RECT -11.780 -82.630 -10.860 -82.150 ;
        RECT -1.860 -82.630 -0.940 -82.150 ;
        RECT 8.060 -82.630 8.980 -82.150 ;
        RECT 17.980 -82.630 18.900 -82.150 ;
        RECT -282.120 -83.610 -280.950 -82.810 ;
        RECT -272.200 -83.610 -271.030 -82.810 ;
        RECT -262.280 -83.610 -261.110 -82.810 ;
        RECT -252.360 -83.610 -251.190 -82.810 ;
        RECT -242.440 -83.610 -241.270 -82.810 ;
        RECT -232.520 -83.610 -231.350 -82.810 ;
        RECT -222.600 -83.610 -221.430 -82.810 ;
        RECT -212.680 -83.610 -211.510 -82.810 ;
        RECT -202.760 -83.610 -201.590 -82.810 ;
        RECT -192.840 -83.610 -191.670 -82.810 ;
        RECT -182.920 -83.610 -181.750 -82.810 ;
        RECT -173.000 -83.610 -171.830 -82.810 ;
        RECT -163.080 -83.610 -161.910 -82.810 ;
        RECT -153.160 -83.610 -151.990 -82.810 ;
        RECT -143.240 -83.610 -142.070 -82.810 ;
        RECT -133.320 -83.610 -132.150 -82.810 ;
        RECT -123.400 -83.610 -122.230 -82.810 ;
        RECT -113.480 -83.610 -112.310 -82.810 ;
        RECT -103.560 -83.610 -102.390 -82.810 ;
        RECT -93.640 -83.610 -92.470 -82.810 ;
        RECT -83.720 -83.610 -82.550 -82.810 ;
        RECT -73.800 -83.610 -72.630 -82.810 ;
        RECT -63.880 -83.610 -62.710 -82.810 ;
        RECT -53.960 -83.610 -52.790 -82.810 ;
        RECT -44.040 -83.610 -42.870 -82.810 ;
        RECT -34.120 -83.610 -32.950 -82.810 ;
        RECT -24.200 -83.610 -23.030 -82.810 ;
        RECT -14.280 -83.610 -13.110 -82.810 ;
        RECT -4.360 -83.610 -3.190 -82.810 ;
        RECT 5.560 -83.610 6.730 -82.810 ;
        RECT 15.480 -83.610 16.650 -82.810 ;
        RECT -291.700 -173.820 -290.530 -173.020 ;
        RECT -281.780 -173.820 -280.610 -173.020 ;
        RECT -271.860 -173.820 -270.690 -173.020 ;
        RECT -261.940 -173.820 -260.770 -173.020 ;
        RECT -252.020 -173.820 -250.850 -173.020 ;
        RECT -242.100 -173.820 -240.930 -173.020 ;
        RECT -232.180 -173.820 -231.010 -173.020 ;
        RECT -222.260 -173.820 -221.090 -173.020 ;
        RECT -212.340 -173.820 -211.170 -173.020 ;
        RECT -202.420 -173.820 -201.250 -173.020 ;
        RECT -192.500 -173.820 -191.330 -173.020 ;
        RECT -182.580 -173.820 -181.410 -173.020 ;
        RECT -172.660 -173.820 -171.490 -173.020 ;
        RECT -162.740 -173.820 -161.570 -173.020 ;
        RECT -152.820 -173.820 -151.650 -173.020 ;
        RECT -142.900 -173.820 -141.730 -173.020 ;
        RECT -132.980 -173.820 -131.810 -173.020 ;
        RECT -123.060 -173.820 -121.890 -173.020 ;
        RECT -113.140 -173.820 -111.970 -173.020 ;
        RECT -103.220 -173.820 -102.050 -173.020 ;
        RECT -93.300 -173.820 -92.130 -173.020 ;
        RECT -83.380 -173.820 -82.210 -173.020 ;
        RECT -73.460 -173.820 -72.290 -173.020 ;
        RECT -63.540 -173.820 -62.370 -173.020 ;
        RECT -53.620 -173.820 -52.450 -173.020 ;
        RECT -43.700 -173.820 -42.530 -173.020 ;
        RECT -33.780 -173.820 -32.610 -173.020 ;
        RECT -23.860 -173.820 -22.690 -173.020 ;
        RECT -13.940 -173.820 -12.770 -173.020 ;
        RECT -4.020 -173.820 -2.850 -173.020 ;
        RECT 5.900 -173.820 7.070 -173.020 ;
        RECT 15.820 -173.820 16.990 -173.020 ;
        RECT -284.040 -174.490 -283.120 -174.010 ;
        RECT -274.120 -174.490 -273.200 -174.010 ;
        RECT -264.200 -174.490 -263.280 -174.010 ;
        RECT -254.280 -174.490 -253.360 -174.010 ;
        RECT -244.360 -174.490 -243.440 -174.010 ;
        RECT -234.440 -174.490 -233.520 -174.010 ;
        RECT -224.520 -174.490 -223.600 -174.010 ;
        RECT -214.600 -174.490 -213.680 -174.010 ;
        RECT -204.680 -174.490 -203.760 -174.010 ;
        RECT -194.760 -174.490 -193.840 -174.010 ;
        RECT -184.840 -174.490 -183.920 -174.010 ;
        RECT -174.920 -174.490 -174.000 -174.010 ;
        RECT -165.000 -174.490 -164.080 -174.010 ;
        RECT -155.080 -174.490 -154.160 -174.010 ;
        RECT -145.160 -174.490 -144.240 -174.010 ;
        RECT -135.240 -174.490 -134.320 -174.010 ;
        RECT -125.320 -174.490 -124.400 -174.010 ;
        RECT -115.400 -174.490 -114.480 -174.010 ;
        RECT -105.480 -174.490 -104.560 -174.010 ;
        RECT -95.560 -174.490 -94.640 -174.010 ;
        RECT -85.640 -174.490 -84.720 -174.010 ;
        RECT -75.720 -174.490 -74.800 -174.010 ;
        RECT -65.800 -174.490 -64.880 -174.010 ;
        RECT -55.880 -174.490 -54.960 -174.010 ;
        RECT -45.960 -174.490 -45.040 -174.010 ;
        RECT -36.040 -174.490 -35.120 -174.010 ;
        RECT -26.120 -174.490 -25.200 -174.010 ;
        RECT -16.200 -174.490 -15.280 -174.010 ;
        RECT -6.280 -174.490 -5.360 -174.010 ;
        RECT 3.640 -174.490 4.560 -174.010 ;
        RECT 13.560 -174.490 14.480 -174.010 ;
        RECT -291.300 -177.210 -290.380 -176.730 ;
        RECT -281.380 -177.210 -280.460 -176.730 ;
        RECT -271.460 -177.210 -270.540 -176.730 ;
        RECT -261.540 -177.210 -260.620 -176.730 ;
        RECT -251.620 -177.210 -250.700 -176.730 ;
        RECT -241.700 -177.210 -240.780 -176.730 ;
        RECT -231.780 -177.210 -230.860 -176.730 ;
        RECT -221.860 -177.210 -220.940 -176.730 ;
        RECT -211.940 -177.210 -211.020 -176.730 ;
        RECT -202.020 -177.210 -201.100 -176.730 ;
        RECT -192.100 -177.210 -191.180 -176.730 ;
        RECT -182.180 -177.210 -181.260 -176.730 ;
        RECT -172.260 -177.210 -171.340 -176.730 ;
        RECT -162.340 -177.210 -161.420 -176.730 ;
        RECT -152.420 -177.210 -151.500 -176.730 ;
        RECT -142.500 -177.210 -141.580 -176.730 ;
        RECT -132.580 -177.210 -131.660 -176.730 ;
        RECT -122.660 -177.210 -121.740 -176.730 ;
        RECT -112.740 -177.210 -111.820 -176.730 ;
        RECT -102.820 -177.210 -101.900 -176.730 ;
        RECT -92.900 -177.210 -91.980 -176.730 ;
        RECT -82.980 -177.210 -82.060 -176.730 ;
        RECT -73.060 -177.210 -72.140 -176.730 ;
        RECT -63.140 -177.210 -62.220 -176.730 ;
        RECT -53.220 -177.210 -52.300 -176.730 ;
        RECT -43.300 -177.210 -42.380 -176.730 ;
        RECT -33.380 -177.210 -32.460 -176.730 ;
        RECT -23.460 -177.210 -22.540 -176.730 ;
        RECT -13.540 -177.210 -12.620 -176.730 ;
        RECT -3.620 -177.210 -2.700 -176.730 ;
        RECT 6.300 -177.210 7.220 -176.730 ;
        RECT 16.220 -177.210 17.140 -176.730 ;
        RECT -283.880 -178.190 -282.710 -177.390 ;
        RECT -273.960 -178.190 -272.790 -177.390 ;
        RECT -264.040 -178.190 -262.870 -177.390 ;
        RECT -254.120 -178.190 -252.950 -177.390 ;
        RECT -244.200 -178.190 -243.030 -177.390 ;
        RECT -234.280 -178.190 -233.110 -177.390 ;
        RECT -224.360 -178.190 -223.190 -177.390 ;
        RECT -214.440 -178.190 -213.270 -177.390 ;
        RECT -204.520 -178.190 -203.350 -177.390 ;
        RECT -194.600 -178.190 -193.430 -177.390 ;
        RECT -184.680 -178.190 -183.510 -177.390 ;
        RECT -174.760 -178.190 -173.590 -177.390 ;
        RECT -164.840 -178.190 -163.670 -177.390 ;
        RECT -154.920 -178.190 -153.750 -177.390 ;
        RECT -145.000 -178.190 -143.830 -177.390 ;
        RECT -135.080 -178.190 -133.910 -177.390 ;
        RECT -125.160 -178.190 -123.990 -177.390 ;
        RECT -115.240 -178.190 -114.070 -177.390 ;
        RECT -105.320 -178.190 -104.150 -177.390 ;
        RECT -95.400 -178.190 -94.230 -177.390 ;
        RECT -85.480 -178.190 -84.310 -177.390 ;
        RECT -75.560 -178.190 -74.390 -177.390 ;
        RECT -65.640 -178.190 -64.470 -177.390 ;
        RECT -55.720 -178.190 -54.550 -177.390 ;
        RECT -45.800 -178.190 -44.630 -177.390 ;
        RECT -35.880 -178.190 -34.710 -177.390 ;
        RECT -25.960 -178.190 -24.790 -177.390 ;
        RECT -16.040 -178.190 -14.870 -177.390 ;
        RECT -6.120 -178.190 -4.950 -177.390 ;
        RECT 3.800 -178.190 4.970 -177.390 ;
        RECT 13.720 -178.190 14.890 -177.390 ;
      LAYER via2 ;
        RECT -287.710 94.060 -287.420 94.340 ;
        RECT -277.790 94.060 -277.500 94.340 ;
        RECT -267.870 94.060 -267.580 94.340 ;
        RECT -257.950 94.060 -257.660 94.340 ;
        RECT -248.030 94.060 -247.740 94.340 ;
        RECT -238.110 94.060 -237.820 94.340 ;
        RECT -228.190 94.060 -227.900 94.340 ;
        RECT -218.270 94.060 -217.980 94.340 ;
        RECT -208.350 94.060 -208.060 94.340 ;
        RECT -198.430 94.060 -198.140 94.340 ;
        RECT -188.510 94.060 -188.220 94.340 ;
        RECT -178.590 94.060 -178.300 94.340 ;
        RECT -168.670 94.060 -168.380 94.340 ;
        RECT -158.750 94.060 -158.460 94.340 ;
        RECT -148.830 94.060 -148.540 94.340 ;
        RECT -138.910 94.060 -138.620 94.340 ;
        RECT -128.990 94.060 -128.700 94.340 ;
        RECT -119.070 94.060 -118.780 94.340 ;
        RECT -109.150 94.060 -108.860 94.340 ;
        RECT -99.230 94.060 -98.940 94.340 ;
        RECT -89.310 94.060 -89.020 94.340 ;
        RECT -79.390 94.060 -79.100 94.340 ;
        RECT -69.470 94.060 -69.180 94.340 ;
        RECT -59.550 94.060 -59.260 94.340 ;
        RECT -49.630 94.060 -49.340 94.340 ;
        RECT -39.710 94.060 -39.420 94.340 ;
        RECT -29.790 94.060 -29.500 94.340 ;
        RECT -19.870 94.060 -19.580 94.340 ;
        RECT -9.950 94.060 -9.660 94.340 ;
        RECT -0.030 94.060 0.260 94.340 ;
        RECT 9.890 94.060 10.180 94.340 ;
        RECT 19.810 94.060 20.100 94.340 ;
        RECT -280.540 93.190 -280.250 93.470 ;
        RECT -280.070 93.190 -279.780 93.470 ;
        RECT -270.620 93.190 -270.330 93.470 ;
        RECT -270.150 93.190 -269.860 93.470 ;
        RECT -260.700 93.190 -260.410 93.470 ;
        RECT -260.230 93.190 -259.940 93.470 ;
        RECT -250.780 93.190 -250.490 93.470 ;
        RECT -250.310 93.190 -250.020 93.470 ;
        RECT -240.860 93.190 -240.570 93.470 ;
        RECT -240.390 93.190 -240.100 93.470 ;
        RECT -230.940 93.190 -230.650 93.470 ;
        RECT -230.470 93.190 -230.180 93.470 ;
        RECT -221.020 93.190 -220.730 93.470 ;
        RECT -220.550 93.190 -220.260 93.470 ;
        RECT -211.100 93.190 -210.810 93.470 ;
        RECT -210.630 93.190 -210.340 93.470 ;
        RECT -201.180 93.190 -200.890 93.470 ;
        RECT -200.710 93.190 -200.420 93.470 ;
        RECT -191.260 93.190 -190.970 93.470 ;
        RECT -190.790 93.190 -190.500 93.470 ;
        RECT -181.340 93.190 -181.050 93.470 ;
        RECT -180.870 93.190 -180.580 93.470 ;
        RECT -171.420 93.190 -171.130 93.470 ;
        RECT -170.950 93.190 -170.660 93.470 ;
        RECT -161.500 93.190 -161.210 93.470 ;
        RECT -161.030 93.190 -160.740 93.470 ;
        RECT -151.580 93.190 -151.290 93.470 ;
        RECT -151.110 93.190 -150.820 93.470 ;
        RECT -141.660 93.190 -141.370 93.470 ;
        RECT -141.190 93.190 -140.900 93.470 ;
        RECT -131.740 93.190 -131.450 93.470 ;
        RECT -131.270 93.190 -130.980 93.470 ;
        RECT -121.820 93.190 -121.530 93.470 ;
        RECT -121.350 93.190 -121.060 93.470 ;
        RECT -111.900 93.190 -111.610 93.470 ;
        RECT -111.430 93.190 -111.140 93.470 ;
        RECT -101.980 93.190 -101.690 93.470 ;
        RECT -101.510 93.190 -101.220 93.470 ;
        RECT -92.060 93.190 -91.770 93.470 ;
        RECT -91.590 93.190 -91.300 93.470 ;
        RECT -82.140 93.190 -81.850 93.470 ;
        RECT -81.670 93.190 -81.380 93.470 ;
        RECT -72.220 93.190 -71.930 93.470 ;
        RECT -71.750 93.190 -71.460 93.470 ;
        RECT -62.300 93.190 -62.010 93.470 ;
        RECT -61.830 93.190 -61.540 93.470 ;
        RECT -52.380 93.190 -52.090 93.470 ;
        RECT -51.910 93.190 -51.620 93.470 ;
        RECT -42.460 93.190 -42.170 93.470 ;
        RECT -41.990 93.190 -41.700 93.470 ;
        RECT -32.540 93.190 -32.250 93.470 ;
        RECT -32.070 93.190 -31.780 93.470 ;
        RECT -22.620 93.190 -22.330 93.470 ;
        RECT -22.150 93.190 -21.860 93.470 ;
        RECT -12.700 93.190 -12.410 93.470 ;
        RECT -12.230 93.190 -11.940 93.470 ;
        RECT -2.780 93.190 -2.490 93.470 ;
        RECT -2.310 93.190 -2.020 93.470 ;
        RECT 7.140 93.190 7.430 93.470 ;
        RECT 7.610 93.190 7.900 93.470 ;
        RECT 17.060 93.190 17.350 93.470 ;
        RECT 17.530 93.190 17.820 93.470 ;
        RECT -287.800 90.460 -287.510 90.740 ;
        RECT -287.340 90.470 -287.050 90.750 ;
        RECT -277.880 90.460 -277.590 90.740 ;
        RECT -277.420 90.470 -277.130 90.750 ;
        RECT -267.960 90.460 -267.670 90.740 ;
        RECT -267.500 90.470 -267.210 90.750 ;
        RECT -258.040 90.460 -257.750 90.740 ;
        RECT -257.580 90.470 -257.290 90.750 ;
        RECT -248.120 90.460 -247.830 90.740 ;
        RECT -247.660 90.470 -247.370 90.750 ;
        RECT -238.200 90.460 -237.910 90.740 ;
        RECT -237.740 90.470 -237.450 90.750 ;
        RECT -228.280 90.460 -227.990 90.740 ;
        RECT -227.820 90.470 -227.530 90.750 ;
        RECT -218.360 90.460 -218.070 90.740 ;
        RECT -217.900 90.470 -217.610 90.750 ;
        RECT -208.440 90.460 -208.150 90.740 ;
        RECT -207.980 90.470 -207.690 90.750 ;
        RECT -198.520 90.460 -198.230 90.740 ;
        RECT -198.060 90.470 -197.770 90.750 ;
        RECT -188.600 90.460 -188.310 90.740 ;
        RECT -188.140 90.470 -187.850 90.750 ;
        RECT -178.680 90.460 -178.390 90.740 ;
        RECT -178.220 90.470 -177.930 90.750 ;
        RECT -168.760 90.460 -168.470 90.740 ;
        RECT -168.300 90.470 -168.010 90.750 ;
        RECT -158.840 90.460 -158.550 90.740 ;
        RECT -158.380 90.470 -158.090 90.750 ;
        RECT -148.920 90.460 -148.630 90.740 ;
        RECT -148.460 90.470 -148.170 90.750 ;
        RECT -139.000 90.460 -138.710 90.740 ;
        RECT -138.540 90.470 -138.250 90.750 ;
        RECT -129.080 90.460 -128.790 90.740 ;
        RECT -128.620 90.470 -128.330 90.750 ;
        RECT -119.160 90.460 -118.870 90.740 ;
        RECT -118.700 90.470 -118.410 90.750 ;
        RECT -109.240 90.460 -108.950 90.740 ;
        RECT -108.780 90.470 -108.490 90.750 ;
        RECT -99.320 90.460 -99.030 90.740 ;
        RECT -98.860 90.470 -98.570 90.750 ;
        RECT -89.400 90.460 -89.110 90.740 ;
        RECT -88.940 90.470 -88.650 90.750 ;
        RECT -79.480 90.460 -79.190 90.740 ;
        RECT -79.020 90.470 -78.730 90.750 ;
        RECT -69.560 90.460 -69.270 90.740 ;
        RECT -69.100 90.470 -68.810 90.750 ;
        RECT -59.640 90.460 -59.350 90.740 ;
        RECT -59.180 90.470 -58.890 90.750 ;
        RECT -49.720 90.460 -49.430 90.740 ;
        RECT -49.260 90.470 -48.970 90.750 ;
        RECT -39.800 90.460 -39.510 90.740 ;
        RECT -39.340 90.470 -39.050 90.750 ;
        RECT -29.880 90.460 -29.590 90.740 ;
        RECT -29.420 90.470 -29.130 90.750 ;
        RECT -19.960 90.460 -19.670 90.740 ;
        RECT -19.500 90.470 -19.210 90.750 ;
        RECT -10.040 90.460 -9.750 90.740 ;
        RECT -9.580 90.470 -9.290 90.750 ;
        RECT -0.120 90.460 0.170 90.740 ;
        RECT 0.340 90.470 0.630 90.750 ;
        RECT 9.800 90.460 10.090 90.740 ;
        RECT 10.260 90.470 10.550 90.750 ;
        RECT 19.720 90.460 20.010 90.740 ;
        RECT 20.180 90.470 20.470 90.750 ;
        RECT -280.150 89.700 -279.860 89.980 ;
        RECT -270.230 89.700 -269.940 89.980 ;
        RECT -260.310 89.700 -260.020 89.980 ;
        RECT -250.390 89.700 -250.100 89.980 ;
        RECT -240.470 89.700 -240.180 89.980 ;
        RECT -230.550 89.700 -230.260 89.980 ;
        RECT -220.630 89.700 -220.340 89.980 ;
        RECT -210.710 89.700 -210.420 89.980 ;
        RECT -200.790 89.700 -200.500 89.980 ;
        RECT -190.870 89.700 -190.580 89.980 ;
        RECT -180.950 89.700 -180.660 89.980 ;
        RECT -171.030 89.700 -170.740 89.980 ;
        RECT -161.110 89.700 -160.820 89.980 ;
        RECT -151.190 89.700 -150.900 89.980 ;
        RECT -141.270 89.700 -140.980 89.980 ;
        RECT -131.350 89.700 -131.060 89.980 ;
        RECT -121.430 89.700 -121.140 89.980 ;
        RECT -111.510 89.700 -111.220 89.980 ;
        RECT -101.590 89.700 -101.300 89.980 ;
        RECT -91.670 89.700 -91.380 89.980 ;
        RECT -81.750 89.700 -81.460 89.980 ;
        RECT -71.830 89.700 -71.540 89.980 ;
        RECT -61.910 89.700 -61.620 89.980 ;
        RECT -51.990 89.700 -51.700 89.980 ;
        RECT -42.070 89.700 -41.780 89.980 ;
        RECT -32.150 89.700 -31.860 89.980 ;
        RECT -22.230 89.700 -21.940 89.980 ;
        RECT -12.310 89.700 -12.020 89.980 ;
        RECT -2.390 89.700 -2.100 89.980 ;
        RECT 7.530 89.700 7.820 89.980 ;
        RECT 17.450 89.700 17.740 89.980 ;
        RECT -289.730 10.010 -289.440 10.290 ;
        RECT -279.810 10.010 -279.520 10.290 ;
        RECT -269.890 10.010 -269.600 10.290 ;
        RECT -259.970 10.010 -259.680 10.290 ;
        RECT -250.050 10.010 -249.760 10.290 ;
        RECT -240.130 10.010 -239.840 10.290 ;
        RECT -230.210 10.010 -229.920 10.290 ;
        RECT -220.290 10.010 -220.000 10.290 ;
        RECT -210.370 10.010 -210.080 10.290 ;
        RECT -200.450 10.010 -200.160 10.290 ;
        RECT -190.530 10.010 -190.240 10.290 ;
        RECT -180.610 10.010 -180.320 10.290 ;
        RECT -170.690 10.010 -170.400 10.290 ;
        RECT -160.770 10.010 -160.480 10.290 ;
        RECT -150.850 10.010 -150.560 10.290 ;
        RECT -140.930 10.010 -140.640 10.290 ;
        RECT -131.010 10.010 -130.720 10.290 ;
        RECT -121.090 10.010 -120.800 10.290 ;
        RECT -111.170 10.010 -110.880 10.290 ;
        RECT -101.250 10.010 -100.960 10.290 ;
        RECT -91.330 10.010 -91.040 10.290 ;
        RECT -81.410 10.010 -81.120 10.290 ;
        RECT -71.490 10.010 -71.200 10.290 ;
        RECT -61.570 10.010 -61.280 10.290 ;
        RECT -51.650 10.010 -51.360 10.290 ;
        RECT -41.730 10.010 -41.440 10.290 ;
        RECT -31.810 10.010 -31.520 10.290 ;
        RECT -21.890 10.010 -21.600 10.290 ;
        RECT -11.970 10.010 -11.680 10.290 ;
        RECT -2.050 10.010 -1.760 10.290 ;
        RECT 7.870 10.010 8.160 10.290 ;
        RECT 17.790 10.010 18.080 10.290 ;
        RECT -282.560 9.140 -282.270 9.420 ;
        RECT -282.090 9.140 -281.800 9.420 ;
        RECT -272.640 9.140 -272.350 9.420 ;
        RECT -272.170 9.140 -271.880 9.420 ;
        RECT -262.720 9.140 -262.430 9.420 ;
        RECT -262.250 9.140 -261.960 9.420 ;
        RECT -252.800 9.140 -252.510 9.420 ;
        RECT -252.330 9.140 -252.040 9.420 ;
        RECT -242.880 9.140 -242.590 9.420 ;
        RECT -242.410 9.140 -242.120 9.420 ;
        RECT -232.960 9.140 -232.670 9.420 ;
        RECT -232.490 9.140 -232.200 9.420 ;
        RECT -223.040 9.140 -222.750 9.420 ;
        RECT -222.570 9.140 -222.280 9.420 ;
        RECT -213.120 9.140 -212.830 9.420 ;
        RECT -212.650 9.140 -212.360 9.420 ;
        RECT -203.200 9.140 -202.910 9.420 ;
        RECT -202.730 9.140 -202.440 9.420 ;
        RECT -193.280 9.140 -192.990 9.420 ;
        RECT -192.810 9.140 -192.520 9.420 ;
        RECT -183.360 9.140 -183.070 9.420 ;
        RECT -182.890 9.140 -182.600 9.420 ;
        RECT -173.440 9.140 -173.150 9.420 ;
        RECT -172.970 9.140 -172.680 9.420 ;
        RECT -163.520 9.140 -163.230 9.420 ;
        RECT -163.050 9.140 -162.760 9.420 ;
        RECT -153.600 9.140 -153.310 9.420 ;
        RECT -153.130 9.140 -152.840 9.420 ;
        RECT -143.680 9.140 -143.390 9.420 ;
        RECT -143.210 9.140 -142.920 9.420 ;
        RECT -133.760 9.140 -133.470 9.420 ;
        RECT -133.290 9.140 -133.000 9.420 ;
        RECT -123.840 9.140 -123.550 9.420 ;
        RECT -123.370 9.140 -123.080 9.420 ;
        RECT -113.920 9.140 -113.630 9.420 ;
        RECT -113.450 9.140 -113.160 9.420 ;
        RECT -104.000 9.140 -103.710 9.420 ;
        RECT -103.530 9.140 -103.240 9.420 ;
        RECT -94.080 9.140 -93.790 9.420 ;
        RECT -93.610 9.140 -93.320 9.420 ;
        RECT -84.160 9.140 -83.870 9.420 ;
        RECT -83.690 9.140 -83.400 9.420 ;
        RECT -74.240 9.140 -73.950 9.420 ;
        RECT -73.770 9.140 -73.480 9.420 ;
        RECT -64.320 9.140 -64.030 9.420 ;
        RECT -63.850 9.140 -63.560 9.420 ;
        RECT -54.400 9.140 -54.110 9.420 ;
        RECT -53.930 9.140 -53.640 9.420 ;
        RECT -44.480 9.140 -44.190 9.420 ;
        RECT -44.010 9.140 -43.720 9.420 ;
        RECT -34.560 9.140 -34.270 9.420 ;
        RECT -34.090 9.140 -33.800 9.420 ;
        RECT -24.640 9.140 -24.350 9.420 ;
        RECT -24.170 9.140 -23.880 9.420 ;
        RECT -14.720 9.140 -14.430 9.420 ;
        RECT -14.250 9.140 -13.960 9.420 ;
        RECT -4.800 9.140 -4.510 9.420 ;
        RECT -4.330 9.140 -4.040 9.420 ;
        RECT 5.120 9.140 5.410 9.420 ;
        RECT 5.590 9.140 5.880 9.420 ;
        RECT 15.040 9.140 15.330 9.420 ;
        RECT 15.510 9.140 15.800 9.420 ;
        RECT -289.820 6.410 -289.530 6.690 ;
        RECT -289.360 6.420 -289.070 6.700 ;
        RECT -279.900 6.410 -279.610 6.690 ;
        RECT -279.440 6.420 -279.150 6.700 ;
        RECT -269.980 6.410 -269.690 6.690 ;
        RECT -269.520 6.420 -269.230 6.700 ;
        RECT -260.060 6.410 -259.770 6.690 ;
        RECT -259.600 6.420 -259.310 6.700 ;
        RECT -250.140 6.410 -249.850 6.690 ;
        RECT -249.680 6.420 -249.390 6.700 ;
        RECT -240.220 6.410 -239.930 6.690 ;
        RECT -239.760 6.420 -239.470 6.700 ;
        RECT -230.300 6.410 -230.010 6.690 ;
        RECT -229.840 6.420 -229.550 6.700 ;
        RECT -220.380 6.410 -220.090 6.690 ;
        RECT -219.920 6.420 -219.630 6.700 ;
        RECT -210.460 6.410 -210.170 6.690 ;
        RECT -210.000 6.420 -209.710 6.700 ;
        RECT -200.540 6.410 -200.250 6.690 ;
        RECT -200.080 6.420 -199.790 6.700 ;
        RECT -190.620 6.410 -190.330 6.690 ;
        RECT -190.160 6.420 -189.870 6.700 ;
        RECT -180.700 6.410 -180.410 6.690 ;
        RECT -180.240 6.420 -179.950 6.700 ;
        RECT -170.780 6.410 -170.490 6.690 ;
        RECT -170.320 6.420 -170.030 6.700 ;
        RECT -160.860 6.410 -160.570 6.690 ;
        RECT -160.400 6.420 -160.110 6.700 ;
        RECT -150.940 6.410 -150.650 6.690 ;
        RECT -150.480 6.420 -150.190 6.700 ;
        RECT -141.020 6.410 -140.730 6.690 ;
        RECT -140.560 6.420 -140.270 6.700 ;
        RECT -131.100 6.410 -130.810 6.690 ;
        RECT -130.640 6.420 -130.350 6.700 ;
        RECT -121.180 6.410 -120.890 6.690 ;
        RECT -120.720 6.420 -120.430 6.700 ;
        RECT -111.260 6.410 -110.970 6.690 ;
        RECT -110.800 6.420 -110.510 6.700 ;
        RECT -101.340 6.410 -101.050 6.690 ;
        RECT -100.880 6.420 -100.590 6.700 ;
        RECT -91.420 6.410 -91.130 6.690 ;
        RECT -90.960 6.420 -90.670 6.700 ;
        RECT -81.500 6.410 -81.210 6.690 ;
        RECT -81.040 6.420 -80.750 6.700 ;
        RECT -71.580 6.410 -71.290 6.690 ;
        RECT -71.120 6.420 -70.830 6.700 ;
        RECT -61.660 6.410 -61.370 6.690 ;
        RECT -61.200 6.420 -60.910 6.700 ;
        RECT -51.740 6.410 -51.450 6.690 ;
        RECT -51.280 6.420 -50.990 6.700 ;
        RECT -41.820 6.410 -41.530 6.690 ;
        RECT -41.360 6.420 -41.070 6.700 ;
        RECT -31.900 6.410 -31.610 6.690 ;
        RECT -31.440 6.420 -31.150 6.700 ;
        RECT -21.980 6.410 -21.690 6.690 ;
        RECT -21.520 6.420 -21.230 6.700 ;
        RECT -12.060 6.410 -11.770 6.690 ;
        RECT -11.600 6.420 -11.310 6.700 ;
        RECT -2.140 6.410 -1.850 6.690 ;
        RECT -1.680 6.420 -1.390 6.700 ;
        RECT 7.780 6.410 8.070 6.690 ;
        RECT 8.240 6.420 8.530 6.700 ;
        RECT 17.700 6.410 17.990 6.690 ;
        RECT 18.160 6.420 18.450 6.700 ;
        RECT -282.170 5.650 -281.880 5.930 ;
        RECT -272.250 5.650 -271.960 5.930 ;
        RECT -262.330 5.650 -262.040 5.930 ;
        RECT -252.410 5.650 -252.120 5.930 ;
        RECT -242.490 5.650 -242.200 5.930 ;
        RECT -232.570 5.650 -232.280 5.930 ;
        RECT -222.650 5.650 -222.360 5.930 ;
        RECT -212.730 5.650 -212.440 5.930 ;
        RECT -202.810 5.650 -202.520 5.930 ;
        RECT -192.890 5.650 -192.600 5.930 ;
        RECT -182.970 5.650 -182.680 5.930 ;
        RECT -173.050 5.650 -172.760 5.930 ;
        RECT -163.130 5.650 -162.840 5.930 ;
        RECT -153.210 5.650 -152.920 5.930 ;
        RECT -143.290 5.650 -143.000 5.930 ;
        RECT -133.370 5.650 -133.080 5.930 ;
        RECT -123.450 5.650 -123.160 5.930 ;
        RECT -113.530 5.650 -113.240 5.930 ;
        RECT -103.610 5.650 -103.320 5.930 ;
        RECT -93.690 5.650 -93.400 5.930 ;
        RECT -83.770 5.650 -83.480 5.930 ;
        RECT -73.850 5.650 -73.560 5.930 ;
        RECT -63.930 5.650 -63.640 5.930 ;
        RECT -54.010 5.650 -53.720 5.930 ;
        RECT -44.090 5.650 -43.800 5.930 ;
        RECT -34.170 5.650 -33.880 5.930 ;
        RECT -24.250 5.650 -23.960 5.930 ;
        RECT -14.330 5.650 -14.040 5.930 ;
        RECT -4.410 5.650 -4.120 5.930 ;
        RECT 5.510 5.650 5.800 5.930 ;
        RECT 15.430 5.650 15.720 5.930 ;
        RECT -289.370 -78.940 -289.080 -78.660 ;
        RECT -279.450 -78.940 -279.160 -78.660 ;
        RECT -269.530 -78.940 -269.240 -78.660 ;
        RECT -259.610 -78.940 -259.320 -78.660 ;
        RECT -249.690 -78.940 -249.400 -78.660 ;
        RECT -239.770 -78.940 -239.480 -78.660 ;
        RECT -229.850 -78.940 -229.560 -78.660 ;
        RECT -219.930 -78.940 -219.640 -78.660 ;
        RECT -210.010 -78.940 -209.720 -78.660 ;
        RECT -200.090 -78.940 -199.800 -78.660 ;
        RECT -190.170 -78.940 -189.880 -78.660 ;
        RECT -180.250 -78.940 -179.960 -78.660 ;
        RECT -170.330 -78.940 -170.040 -78.660 ;
        RECT -160.410 -78.940 -160.120 -78.660 ;
        RECT -150.490 -78.940 -150.200 -78.660 ;
        RECT -140.570 -78.940 -140.280 -78.660 ;
        RECT -130.650 -78.940 -130.360 -78.660 ;
        RECT -120.730 -78.940 -120.440 -78.660 ;
        RECT -110.810 -78.940 -110.520 -78.660 ;
        RECT -100.890 -78.940 -100.600 -78.660 ;
        RECT -90.970 -78.940 -90.680 -78.660 ;
        RECT -81.050 -78.940 -80.760 -78.660 ;
        RECT -71.130 -78.940 -70.840 -78.660 ;
        RECT -61.210 -78.940 -60.920 -78.660 ;
        RECT -51.290 -78.940 -51.000 -78.660 ;
        RECT -41.370 -78.940 -41.080 -78.660 ;
        RECT -31.450 -78.940 -31.160 -78.660 ;
        RECT -21.530 -78.940 -21.240 -78.660 ;
        RECT -11.610 -78.940 -11.320 -78.660 ;
        RECT -1.690 -78.940 -1.400 -78.660 ;
        RECT 8.230 -78.940 8.520 -78.660 ;
        RECT 18.150 -78.940 18.440 -78.660 ;
        RECT -282.200 -79.810 -281.910 -79.530 ;
        RECT -281.730 -79.810 -281.440 -79.530 ;
        RECT -272.280 -79.810 -271.990 -79.530 ;
        RECT -271.810 -79.810 -271.520 -79.530 ;
        RECT -262.360 -79.810 -262.070 -79.530 ;
        RECT -261.890 -79.810 -261.600 -79.530 ;
        RECT -252.440 -79.810 -252.150 -79.530 ;
        RECT -251.970 -79.810 -251.680 -79.530 ;
        RECT -242.520 -79.810 -242.230 -79.530 ;
        RECT -242.050 -79.810 -241.760 -79.530 ;
        RECT -232.600 -79.810 -232.310 -79.530 ;
        RECT -232.130 -79.810 -231.840 -79.530 ;
        RECT -222.680 -79.810 -222.390 -79.530 ;
        RECT -222.210 -79.810 -221.920 -79.530 ;
        RECT -212.760 -79.810 -212.470 -79.530 ;
        RECT -212.290 -79.810 -212.000 -79.530 ;
        RECT -202.840 -79.810 -202.550 -79.530 ;
        RECT -202.370 -79.810 -202.080 -79.530 ;
        RECT -192.920 -79.810 -192.630 -79.530 ;
        RECT -192.450 -79.810 -192.160 -79.530 ;
        RECT -183.000 -79.810 -182.710 -79.530 ;
        RECT -182.530 -79.810 -182.240 -79.530 ;
        RECT -173.080 -79.810 -172.790 -79.530 ;
        RECT -172.610 -79.810 -172.320 -79.530 ;
        RECT -163.160 -79.810 -162.870 -79.530 ;
        RECT -162.690 -79.810 -162.400 -79.530 ;
        RECT -153.240 -79.810 -152.950 -79.530 ;
        RECT -152.770 -79.810 -152.480 -79.530 ;
        RECT -143.320 -79.810 -143.030 -79.530 ;
        RECT -142.850 -79.810 -142.560 -79.530 ;
        RECT -133.400 -79.810 -133.110 -79.530 ;
        RECT -132.930 -79.810 -132.640 -79.530 ;
        RECT -123.480 -79.810 -123.190 -79.530 ;
        RECT -123.010 -79.810 -122.720 -79.530 ;
        RECT -113.560 -79.810 -113.270 -79.530 ;
        RECT -113.090 -79.810 -112.800 -79.530 ;
        RECT -103.640 -79.810 -103.350 -79.530 ;
        RECT -103.170 -79.810 -102.880 -79.530 ;
        RECT -93.720 -79.810 -93.430 -79.530 ;
        RECT -93.250 -79.810 -92.960 -79.530 ;
        RECT -83.800 -79.810 -83.510 -79.530 ;
        RECT -83.330 -79.810 -83.040 -79.530 ;
        RECT -73.880 -79.810 -73.590 -79.530 ;
        RECT -73.410 -79.810 -73.120 -79.530 ;
        RECT -63.960 -79.810 -63.670 -79.530 ;
        RECT -63.490 -79.810 -63.200 -79.530 ;
        RECT -54.040 -79.810 -53.750 -79.530 ;
        RECT -53.570 -79.810 -53.280 -79.530 ;
        RECT -44.120 -79.810 -43.830 -79.530 ;
        RECT -43.650 -79.810 -43.360 -79.530 ;
        RECT -34.200 -79.810 -33.910 -79.530 ;
        RECT -33.730 -79.810 -33.440 -79.530 ;
        RECT -24.280 -79.810 -23.990 -79.530 ;
        RECT -23.810 -79.810 -23.520 -79.530 ;
        RECT -14.360 -79.810 -14.070 -79.530 ;
        RECT -13.890 -79.810 -13.600 -79.530 ;
        RECT -4.440 -79.810 -4.150 -79.530 ;
        RECT -3.970 -79.810 -3.680 -79.530 ;
        RECT 5.480 -79.810 5.770 -79.530 ;
        RECT 5.950 -79.810 6.240 -79.530 ;
        RECT 15.400 -79.810 15.690 -79.530 ;
        RECT 15.870 -79.810 16.160 -79.530 ;
        RECT -289.460 -82.540 -289.170 -82.260 ;
        RECT -289.000 -82.530 -288.710 -82.250 ;
        RECT -279.540 -82.540 -279.250 -82.260 ;
        RECT -279.080 -82.530 -278.790 -82.250 ;
        RECT -269.620 -82.540 -269.330 -82.260 ;
        RECT -269.160 -82.530 -268.870 -82.250 ;
        RECT -259.700 -82.540 -259.410 -82.260 ;
        RECT -259.240 -82.530 -258.950 -82.250 ;
        RECT -249.780 -82.540 -249.490 -82.260 ;
        RECT -249.320 -82.530 -249.030 -82.250 ;
        RECT -239.860 -82.540 -239.570 -82.260 ;
        RECT -239.400 -82.530 -239.110 -82.250 ;
        RECT -229.940 -82.540 -229.650 -82.260 ;
        RECT -229.480 -82.530 -229.190 -82.250 ;
        RECT -220.020 -82.540 -219.730 -82.260 ;
        RECT -219.560 -82.530 -219.270 -82.250 ;
        RECT -210.100 -82.540 -209.810 -82.260 ;
        RECT -209.640 -82.530 -209.350 -82.250 ;
        RECT -200.180 -82.540 -199.890 -82.260 ;
        RECT -199.720 -82.530 -199.430 -82.250 ;
        RECT -190.260 -82.540 -189.970 -82.260 ;
        RECT -189.800 -82.530 -189.510 -82.250 ;
        RECT -180.340 -82.540 -180.050 -82.260 ;
        RECT -179.880 -82.530 -179.590 -82.250 ;
        RECT -170.420 -82.540 -170.130 -82.260 ;
        RECT -169.960 -82.530 -169.670 -82.250 ;
        RECT -160.500 -82.540 -160.210 -82.260 ;
        RECT -160.040 -82.530 -159.750 -82.250 ;
        RECT -150.580 -82.540 -150.290 -82.260 ;
        RECT -150.120 -82.530 -149.830 -82.250 ;
        RECT -140.660 -82.540 -140.370 -82.260 ;
        RECT -140.200 -82.530 -139.910 -82.250 ;
        RECT -130.740 -82.540 -130.450 -82.260 ;
        RECT -130.280 -82.530 -129.990 -82.250 ;
        RECT -120.820 -82.540 -120.530 -82.260 ;
        RECT -120.360 -82.530 -120.070 -82.250 ;
        RECT -110.900 -82.540 -110.610 -82.260 ;
        RECT -110.440 -82.530 -110.150 -82.250 ;
        RECT -100.980 -82.540 -100.690 -82.260 ;
        RECT -100.520 -82.530 -100.230 -82.250 ;
        RECT -91.060 -82.540 -90.770 -82.260 ;
        RECT -90.600 -82.530 -90.310 -82.250 ;
        RECT -81.140 -82.540 -80.850 -82.260 ;
        RECT -80.680 -82.530 -80.390 -82.250 ;
        RECT -71.220 -82.540 -70.930 -82.260 ;
        RECT -70.760 -82.530 -70.470 -82.250 ;
        RECT -61.300 -82.540 -61.010 -82.260 ;
        RECT -60.840 -82.530 -60.550 -82.250 ;
        RECT -51.380 -82.540 -51.090 -82.260 ;
        RECT -50.920 -82.530 -50.630 -82.250 ;
        RECT -41.460 -82.540 -41.170 -82.260 ;
        RECT -41.000 -82.530 -40.710 -82.250 ;
        RECT -31.540 -82.540 -31.250 -82.260 ;
        RECT -31.080 -82.530 -30.790 -82.250 ;
        RECT -21.620 -82.540 -21.330 -82.260 ;
        RECT -21.160 -82.530 -20.870 -82.250 ;
        RECT -11.700 -82.540 -11.410 -82.260 ;
        RECT -11.240 -82.530 -10.950 -82.250 ;
        RECT -1.780 -82.540 -1.490 -82.260 ;
        RECT -1.320 -82.530 -1.030 -82.250 ;
        RECT 8.140 -82.540 8.430 -82.260 ;
        RECT 8.600 -82.530 8.890 -82.250 ;
        RECT 18.060 -82.540 18.350 -82.260 ;
        RECT 18.520 -82.530 18.810 -82.250 ;
        RECT -281.810 -83.300 -281.520 -83.020 ;
        RECT -271.890 -83.300 -271.600 -83.020 ;
        RECT -261.970 -83.300 -261.680 -83.020 ;
        RECT -252.050 -83.300 -251.760 -83.020 ;
        RECT -242.130 -83.300 -241.840 -83.020 ;
        RECT -232.210 -83.300 -231.920 -83.020 ;
        RECT -222.290 -83.300 -222.000 -83.020 ;
        RECT -212.370 -83.300 -212.080 -83.020 ;
        RECT -202.450 -83.300 -202.160 -83.020 ;
        RECT -192.530 -83.300 -192.240 -83.020 ;
        RECT -182.610 -83.300 -182.320 -83.020 ;
        RECT -172.690 -83.300 -172.400 -83.020 ;
        RECT -162.770 -83.300 -162.480 -83.020 ;
        RECT -152.850 -83.300 -152.560 -83.020 ;
        RECT -142.930 -83.300 -142.640 -83.020 ;
        RECT -133.010 -83.300 -132.720 -83.020 ;
        RECT -123.090 -83.300 -122.800 -83.020 ;
        RECT -113.170 -83.300 -112.880 -83.020 ;
        RECT -103.250 -83.300 -102.960 -83.020 ;
        RECT -93.330 -83.300 -93.040 -83.020 ;
        RECT -83.410 -83.300 -83.120 -83.020 ;
        RECT -73.490 -83.300 -73.200 -83.020 ;
        RECT -63.570 -83.300 -63.280 -83.020 ;
        RECT -53.650 -83.300 -53.360 -83.020 ;
        RECT -43.730 -83.300 -43.440 -83.020 ;
        RECT -33.810 -83.300 -33.520 -83.020 ;
        RECT -23.890 -83.300 -23.600 -83.020 ;
        RECT -13.970 -83.300 -13.680 -83.020 ;
        RECT -4.050 -83.300 -3.760 -83.020 ;
        RECT 5.870 -83.300 6.160 -83.020 ;
        RECT 15.790 -83.300 16.080 -83.020 ;
        RECT -291.130 -173.520 -290.840 -173.240 ;
        RECT -281.210 -173.520 -280.920 -173.240 ;
        RECT -271.290 -173.520 -271.000 -173.240 ;
        RECT -261.370 -173.520 -261.080 -173.240 ;
        RECT -251.450 -173.520 -251.160 -173.240 ;
        RECT -241.530 -173.520 -241.240 -173.240 ;
        RECT -231.610 -173.520 -231.320 -173.240 ;
        RECT -221.690 -173.520 -221.400 -173.240 ;
        RECT -211.770 -173.520 -211.480 -173.240 ;
        RECT -201.850 -173.520 -201.560 -173.240 ;
        RECT -191.930 -173.520 -191.640 -173.240 ;
        RECT -182.010 -173.520 -181.720 -173.240 ;
        RECT -172.090 -173.520 -171.800 -173.240 ;
        RECT -162.170 -173.520 -161.880 -173.240 ;
        RECT -152.250 -173.520 -151.960 -173.240 ;
        RECT -142.330 -173.520 -142.040 -173.240 ;
        RECT -132.410 -173.520 -132.120 -173.240 ;
        RECT -122.490 -173.520 -122.200 -173.240 ;
        RECT -112.570 -173.520 -112.280 -173.240 ;
        RECT -102.650 -173.520 -102.360 -173.240 ;
        RECT -92.730 -173.520 -92.440 -173.240 ;
        RECT -82.810 -173.520 -82.520 -173.240 ;
        RECT -72.890 -173.520 -72.600 -173.240 ;
        RECT -62.970 -173.520 -62.680 -173.240 ;
        RECT -53.050 -173.520 -52.760 -173.240 ;
        RECT -43.130 -173.520 -42.840 -173.240 ;
        RECT -33.210 -173.520 -32.920 -173.240 ;
        RECT -23.290 -173.520 -23.000 -173.240 ;
        RECT -13.370 -173.520 -13.080 -173.240 ;
        RECT -3.450 -173.520 -3.160 -173.240 ;
        RECT 6.470 -173.520 6.760 -173.240 ;
        RECT 16.390 -173.520 16.680 -173.240 ;
        RECT -283.960 -174.390 -283.670 -174.110 ;
        RECT -283.490 -174.390 -283.200 -174.110 ;
        RECT -274.040 -174.390 -273.750 -174.110 ;
        RECT -273.570 -174.390 -273.280 -174.110 ;
        RECT -264.120 -174.390 -263.830 -174.110 ;
        RECT -263.650 -174.390 -263.360 -174.110 ;
        RECT -254.200 -174.390 -253.910 -174.110 ;
        RECT -253.730 -174.390 -253.440 -174.110 ;
        RECT -244.280 -174.390 -243.990 -174.110 ;
        RECT -243.810 -174.390 -243.520 -174.110 ;
        RECT -234.360 -174.390 -234.070 -174.110 ;
        RECT -233.890 -174.390 -233.600 -174.110 ;
        RECT -224.440 -174.390 -224.150 -174.110 ;
        RECT -223.970 -174.390 -223.680 -174.110 ;
        RECT -214.520 -174.390 -214.230 -174.110 ;
        RECT -214.050 -174.390 -213.760 -174.110 ;
        RECT -204.600 -174.390 -204.310 -174.110 ;
        RECT -204.130 -174.390 -203.840 -174.110 ;
        RECT -194.680 -174.390 -194.390 -174.110 ;
        RECT -194.210 -174.390 -193.920 -174.110 ;
        RECT -184.760 -174.390 -184.470 -174.110 ;
        RECT -184.290 -174.390 -184.000 -174.110 ;
        RECT -174.840 -174.390 -174.550 -174.110 ;
        RECT -174.370 -174.390 -174.080 -174.110 ;
        RECT -164.920 -174.390 -164.630 -174.110 ;
        RECT -164.450 -174.390 -164.160 -174.110 ;
        RECT -155.000 -174.390 -154.710 -174.110 ;
        RECT -154.530 -174.390 -154.240 -174.110 ;
        RECT -145.080 -174.390 -144.790 -174.110 ;
        RECT -144.610 -174.390 -144.320 -174.110 ;
        RECT -135.160 -174.390 -134.870 -174.110 ;
        RECT -134.690 -174.390 -134.400 -174.110 ;
        RECT -125.240 -174.390 -124.950 -174.110 ;
        RECT -124.770 -174.390 -124.480 -174.110 ;
        RECT -115.320 -174.390 -115.030 -174.110 ;
        RECT -114.850 -174.390 -114.560 -174.110 ;
        RECT -105.400 -174.390 -105.110 -174.110 ;
        RECT -104.930 -174.390 -104.640 -174.110 ;
        RECT -95.480 -174.390 -95.190 -174.110 ;
        RECT -95.010 -174.390 -94.720 -174.110 ;
        RECT -85.560 -174.390 -85.270 -174.110 ;
        RECT -85.090 -174.390 -84.800 -174.110 ;
        RECT -75.640 -174.390 -75.350 -174.110 ;
        RECT -75.170 -174.390 -74.880 -174.110 ;
        RECT -65.720 -174.390 -65.430 -174.110 ;
        RECT -65.250 -174.390 -64.960 -174.110 ;
        RECT -55.800 -174.390 -55.510 -174.110 ;
        RECT -55.330 -174.390 -55.040 -174.110 ;
        RECT -45.880 -174.390 -45.590 -174.110 ;
        RECT -45.410 -174.390 -45.120 -174.110 ;
        RECT -35.960 -174.390 -35.670 -174.110 ;
        RECT -35.490 -174.390 -35.200 -174.110 ;
        RECT -26.040 -174.390 -25.750 -174.110 ;
        RECT -25.570 -174.390 -25.280 -174.110 ;
        RECT -16.120 -174.390 -15.830 -174.110 ;
        RECT -15.650 -174.390 -15.360 -174.110 ;
        RECT -6.200 -174.390 -5.910 -174.110 ;
        RECT -5.730 -174.390 -5.440 -174.110 ;
        RECT 3.720 -174.390 4.010 -174.110 ;
        RECT 4.190 -174.390 4.480 -174.110 ;
        RECT 13.640 -174.390 13.930 -174.110 ;
        RECT 14.110 -174.390 14.400 -174.110 ;
        RECT -291.220 -177.120 -290.930 -176.840 ;
        RECT -290.760 -177.110 -290.470 -176.830 ;
        RECT -281.300 -177.120 -281.010 -176.840 ;
        RECT -280.840 -177.110 -280.550 -176.830 ;
        RECT -271.380 -177.120 -271.090 -176.840 ;
        RECT -270.920 -177.110 -270.630 -176.830 ;
        RECT -261.460 -177.120 -261.170 -176.840 ;
        RECT -261.000 -177.110 -260.710 -176.830 ;
        RECT -251.540 -177.120 -251.250 -176.840 ;
        RECT -251.080 -177.110 -250.790 -176.830 ;
        RECT -241.620 -177.120 -241.330 -176.840 ;
        RECT -241.160 -177.110 -240.870 -176.830 ;
        RECT -231.700 -177.120 -231.410 -176.840 ;
        RECT -231.240 -177.110 -230.950 -176.830 ;
        RECT -221.780 -177.120 -221.490 -176.840 ;
        RECT -221.320 -177.110 -221.030 -176.830 ;
        RECT -211.860 -177.120 -211.570 -176.840 ;
        RECT -211.400 -177.110 -211.110 -176.830 ;
        RECT -201.940 -177.120 -201.650 -176.840 ;
        RECT -201.480 -177.110 -201.190 -176.830 ;
        RECT -192.020 -177.120 -191.730 -176.840 ;
        RECT -191.560 -177.110 -191.270 -176.830 ;
        RECT -182.100 -177.120 -181.810 -176.840 ;
        RECT -181.640 -177.110 -181.350 -176.830 ;
        RECT -172.180 -177.120 -171.890 -176.840 ;
        RECT -171.720 -177.110 -171.430 -176.830 ;
        RECT -162.260 -177.120 -161.970 -176.840 ;
        RECT -161.800 -177.110 -161.510 -176.830 ;
        RECT -152.340 -177.120 -152.050 -176.840 ;
        RECT -151.880 -177.110 -151.590 -176.830 ;
        RECT -142.420 -177.120 -142.130 -176.840 ;
        RECT -141.960 -177.110 -141.670 -176.830 ;
        RECT -132.500 -177.120 -132.210 -176.840 ;
        RECT -132.040 -177.110 -131.750 -176.830 ;
        RECT -122.580 -177.120 -122.290 -176.840 ;
        RECT -122.120 -177.110 -121.830 -176.830 ;
        RECT -112.660 -177.120 -112.370 -176.840 ;
        RECT -112.200 -177.110 -111.910 -176.830 ;
        RECT -102.740 -177.120 -102.450 -176.840 ;
        RECT -102.280 -177.110 -101.990 -176.830 ;
        RECT -92.820 -177.120 -92.530 -176.840 ;
        RECT -92.360 -177.110 -92.070 -176.830 ;
        RECT -82.900 -177.120 -82.610 -176.840 ;
        RECT -82.440 -177.110 -82.150 -176.830 ;
        RECT -72.980 -177.120 -72.690 -176.840 ;
        RECT -72.520 -177.110 -72.230 -176.830 ;
        RECT -63.060 -177.120 -62.770 -176.840 ;
        RECT -62.600 -177.110 -62.310 -176.830 ;
        RECT -53.140 -177.120 -52.850 -176.840 ;
        RECT -52.680 -177.110 -52.390 -176.830 ;
        RECT -43.220 -177.120 -42.930 -176.840 ;
        RECT -42.760 -177.110 -42.470 -176.830 ;
        RECT -33.300 -177.120 -33.010 -176.840 ;
        RECT -32.840 -177.110 -32.550 -176.830 ;
        RECT -23.380 -177.120 -23.090 -176.840 ;
        RECT -22.920 -177.110 -22.630 -176.830 ;
        RECT -13.460 -177.120 -13.170 -176.840 ;
        RECT -13.000 -177.110 -12.710 -176.830 ;
        RECT -3.540 -177.120 -3.250 -176.840 ;
        RECT -3.080 -177.110 -2.790 -176.830 ;
        RECT 6.380 -177.120 6.670 -176.840 ;
        RECT 6.840 -177.110 7.130 -176.830 ;
        RECT 16.300 -177.120 16.590 -176.840 ;
        RECT 16.760 -177.110 17.050 -176.830 ;
        RECT -283.570 -177.880 -283.280 -177.600 ;
        RECT -273.650 -177.880 -273.360 -177.600 ;
        RECT -263.730 -177.880 -263.440 -177.600 ;
        RECT -253.810 -177.880 -253.520 -177.600 ;
        RECT -243.890 -177.880 -243.600 -177.600 ;
        RECT -233.970 -177.880 -233.680 -177.600 ;
        RECT -224.050 -177.880 -223.760 -177.600 ;
        RECT -214.130 -177.880 -213.840 -177.600 ;
        RECT -204.210 -177.880 -203.920 -177.600 ;
        RECT -194.290 -177.880 -194.000 -177.600 ;
        RECT -184.370 -177.880 -184.080 -177.600 ;
        RECT -174.450 -177.880 -174.160 -177.600 ;
        RECT -164.530 -177.880 -164.240 -177.600 ;
        RECT -154.610 -177.880 -154.320 -177.600 ;
        RECT -144.690 -177.880 -144.400 -177.600 ;
        RECT -134.770 -177.880 -134.480 -177.600 ;
        RECT -124.850 -177.880 -124.560 -177.600 ;
        RECT -114.930 -177.880 -114.640 -177.600 ;
        RECT -105.010 -177.880 -104.720 -177.600 ;
        RECT -95.090 -177.880 -94.800 -177.600 ;
        RECT -85.170 -177.880 -84.880 -177.600 ;
        RECT -75.250 -177.880 -74.960 -177.600 ;
        RECT -65.330 -177.880 -65.040 -177.600 ;
        RECT -55.410 -177.880 -55.120 -177.600 ;
        RECT -45.490 -177.880 -45.200 -177.600 ;
        RECT -35.570 -177.880 -35.280 -177.600 ;
        RECT -25.650 -177.880 -25.360 -177.600 ;
        RECT -15.730 -177.880 -15.440 -177.600 ;
        RECT -5.810 -177.880 -5.520 -177.600 ;
        RECT 4.110 -177.880 4.400 -177.600 ;
        RECT 14.030 -177.880 14.320 -177.600 ;
      LAYER met3 ;
        RECT -288.280 93.760 -287.110 94.560 ;
        RECT -278.360 93.760 -277.190 94.560 ;
        RECT -268.440 93.760 -267.270 94.560 ;
        RECT -258.520 93.760 -257.350 94.560 ;
        RECT -248.600 93.760 -247.430 94.560 ;
        RECT -238.680 93.760 -237.510 94.560 ;
        RECT -228.760 93.760 -227.590 94.560 ;
        RECT -218.840 93.760 -217.670 94.560 ;
        RECT -208.920 93.760 -207.750 94.560 ;
        RECT -199.000 93.760 -197.830 94.560 ;
        RECT -189.080 93.760 -187.910 94.560 ;
        RECT -179.160 93.760 -177.990 94.560 ;
        RECT -169.240 93.760 -168.070 94.560 ;
        RECT -159.320 93.760 -158.150 94.560 ;
        RECT -149.400 93.760 -148.230 94.560 ;
        RECT -139.480 93.760 -138.310 94.560 ;
        RECT -129.560 93.760 -128.390 94.560 ;
        RECT -119.640 93.760 -118.470 94.560 ;
        RECT -109.720 93.760 -108.550 94.560 ;
        RECT -99.800 93.760 -98.630 94.560 ;
        RECT -89.880 93.760 -88.710 94.560 ;
        RECT -79.960 93.760 -78.790 94.560 ;
        RECT -70.040 93.760 -68.870 94.560 ;
        RECT -60.120 93.760 -58.950 94.560 ;
        RECT -50.200 93.760 -49.030 94.560 ;
        RECT -40.280 93.760 -39.110 94.560 ;
        RECT -30.360 93.760 -29.190 94.560 ;
        RECT -20.440 93.760 -19.270 94.560 ;
        RECT -10.520 93.760 -9.350 94.560 ;
        RECT -0.600 93.760 0.570 94.560 ;
        RECT 9.320 93.760 10.490 94.560 ;
        RECT 19.240 93.760 20.410 94.560 ;
        RECT -280.620 93.090 -279.700 93.570 ;
        RECT -270.700 93.090 -269.780 93.570 ;
        RECT -260.780 93.090 -259.860 93.570 ;
        RECT -250.860 93.090 -249.940 93.570 ;
        RECT -240.940 93.090 -240.020 93.570 ;
        RECT -231.020 93.090 -230.100 93.570 ;
        RECT -221.100 93.090 -220.180 93.570 ;
        RECT -211.180 93.090 -210.260 93.570 ;
        RECT -201.260 93.090 -200.340 93.570 ;
        RECT -191.340 93.090 -190.420 93.570 ;
        RECT -181.420 93.090 -180.500 93.570 ;
        RECT -171.500 93.090 -170.580 93.570 ;
        RECT -161.580 93.090 -160.660 93.570 ;
        RECT -151.660 93.090 -150.740 93.570 ;
        RECT -141.740 93.090 -140.820 93.570 ;
        RECT -131.820 93.090 -130.900 93.570 ;
        RECT -121.900 93.090 -120.980 93.570 ;
        RECT -111.980 93.090 -111.060 93.570 ;
        RECT -102.060 93.090 -101.140 93.570 ;
        RECT -92.140 93.090 -91.220 93.570 ;
        RECT -82.220 93.090 -81.300 93.570 ;
        RECT -72.300 93.090 -71.380 93.570 ;
        RECT -62.380 93.090 -61.460 93.570 ;
        RECT -52.460 93.090 -51.540 93.570 ;
        RECT -42.540 93.090 -41.620 93.570 ;
        RECT -32.620 93.090 -31.700 93.570 ;
        RECT -22.700 93.090 -21.780 93.570 ;
        RECT -12.780 93.090 -11.860 93.570 ;
        RECT -2.860 93.090 -1.940 93.570 ;
        RECT 7.060 93.090 7.980 93.570 ;
        RECT 16.980 93.090 17.900 93.570 ;
        RECT -287.880 90.370 -286.960 90.850 ;
        RECT -277.960 90.370 -277.060 90.850 ;
        RECT -268.040 90.370 -267.120 90.850 ;
        RECT -258.120 90.370 -257.200 90.850 ;
        RECT -248.200 90.370 -247.280 90.850 ;
        RECT -238.280 90.370 -237.360 90.850 ;
        RECT -228.360 90.370 -227.440 90.850 ;
        RECT -218.440 90.370 -217.520 90.850 ;
        RECT -208.520 90.370 -207.600 90.850 ;
        RECT -198.600 90.370 -197.680 90.850 ;
        RECT -188.680 90.370 -187.760 90.850 ;
        RECT -178.760 90.370 -177.840 90.850 ;
        RECT -168.840 90.370 -167.920 90.850 ;
        RECT -158.920 90.370 -158.000 90.850 ;
        RECT -149.000 90.370 -148.080 90.850 ;
        RECT -139.080 90.370 -138.160 90.850 ;
        RECT -129.160 90.370 -128.240 90.850 ;
        RECT -119.240 90.370 -118.320 90.850 ;
        RECT -109.320 90.370 -108.400 90.850 ;
        RECT -99.400 90.370 -98.480 90.850 ;
        RECT -89.480 90.370 -88.560 90.850 ;
        RECT -79.560 90.370 -78.640 90.850 ;
        RECT -69.640 90.370 -68.720 90.850 ;
        RECT -59.720 90.370 -58.800 90.850 ;
        RECT -49.800 90.370 -48.880 90.850 ;
        RECT -39.880 90.370 -38.960 90.850 ;
        RECT -29.960 90.370 -29.040 90.850 ;
        RECT -20.040 90.370 -19.120 90.850 ;
        RECT -10.120 90.370 -9.200 90.850 ;
        RECT -0.200 90.370 0.720 90.850 ;
        RECT 9.720 90.370 10.640 90.850 ;
        RECT 19.640 90.370 20.560 90.850 ;
        RECT -280.460 89.390 -279.290 90.190 ;
        RECT -270.540 89.390 -269.370 90.190 ;
        RECT -260.620 89.390 -259.450 90.190 ;
        RECT -250.700 89.390 -249.530 90.190 ;
        RECT -240.780 89.390 -239.610 90.190 ;
        RECT -230.860 89.390 -229.690 90.190 ;
        RECT -220.940 89.390 -219.770 90.190 ;
        RECT -211.020 89.390 -209.850 90.190 ;
        RECT -201.100 89.390 -199.930 90.190 ;
        RECT -191.180 89.390 -190.010 90.190 ;
        RECT -181.260 89.390 -180.090 90.190 ;
        RECT -171.340 89.390 -170.170 90.190 ;
        RECT -161.420 89.390 -160.250 90.190 ;
        RECT -151.500 89.390 -150.330 90.190 ;
        RECT -141.580 89.390 -140.410 90.190 ;
        RECT -131.660 89.390 -130.490 90.190 ;
        RECT -121.740 89.390 -120.570 90.190 ;
        RECT -111.820 89.390 -110.650 90.190 ;
        RECT -101.900 89.390 -100.730 90.190 ;
        RECT -91.980 89.390 -90.810 90.190 ;
        RECT -82.060 89.390 -80.890 90.190 ;
        RECT -72.140 89.390 -70.970 90.190 ;
        RECT -62.220 89.390 -61.050 90.190 ;
        RECT -52.300 89.390 -51.130 90.190 ;
        RECT -42.380 89.390 -41.210 90.190 ;
        RECT -32.460 89.390 -31.290 90.190 ;
        RECT -22.540 89.390 -21.370 90.190 ;
        RECT -12.620 89.390 -11.450 90.190 ;
        RECT -2.700 89.390 -1.530 90.190 ;
        RECT 7.220 89.390 8.390 90.190 ;
        RECT 17.140 89.390 18.310 90.190 ;
        RECT -290.300 9.710 -289.130 10.510 ;
        RECT -280.380 9.710 -279.210 10.510 ;
        RECT -270.460 9.710 -269.290 10.510 ;
        RECT -260.540 9.710 -259.370 10.510 ;
        RECT -250.620 9.710 -249.450 10.510 ;
        RECT -240.700 9.710 -239.530 10.510 ;
        RECT -230.780 9.710 -229.610 10.510 ;
        RECT -220.860 9.710 -219.690 10.510 ;
        RECT -210.940 9.710 -209.770 10.510 ;
        RECT -201.020 9.710 -199.850 10.510 ;
        RECT -191.100 9.710 -189.930 10.510 ;
        RECT -181.180 9.710 -180.010 10.510 ;
        RECT -171.260 9.710 -170.090 10.510 ;
        RECT -161.340 9.710 -160.170 10.510 ;
        RECT -151.420 9.710 -150.250 10.510 ;
        RECT -141.500 9.710 -140.330 10.510 ;
        RECT -131.580 9.710 -130.410 10.510 ;
        RECT -121.660 9.710 -120.490 10.510 ;
        RECT -111.740 9.710 -110.570 10.510 ;
        RECT -101.820 9.710 -100.650 10.510 ;
        RECT -91.900 9.710 -90.730 10.510 ;
        RECT -81.980 9.710 -80.810 10.510 ;
        RECT -72.060 9.710 -70.890 10.510 ;
        RECT -62.140 9.710 -60.970 10.510 ;
        RECT -52.220 9.710 -51.050 10.510 ;
        RECT -42.300 9.710 -41.130 10.510 ;
        RECT -32.380 9.710 -31.210 10.510 ;
        RECT -22.460 9.710 -21.290 10.510 ;
        RECT -12.540 9.710 -11.370 10.510 ;
        RECT -2.620 9.710 -1.450 10.510 ;
        RECT 7.300 9.710 8.470 10.510 ;
        RECT 17.220 9.710 18.390 10.510 ;
        RECT -282.640 9.040 -281.720 9.520 ;
        RECT -272.720 9.040 -271.800 9.520 ;
        RECT -262.800 9.040 -261.880 9.520 ;
        RECT -252.880 9.040 -251.960 9.520 ;
        RECT -242.960 9.040 -242.040 9.520 ;
        RECT -233.040 9.040 -232.120 9.520 ;
        RECT -223.120 9.040 -222.200 9.520 ;
        RECT -213.200 9.040 -212.280 9.520 ;
        RECT -203.280 9.040 -202.360 9.520 ;
        RECT -193.360 9.040 -192.440 9.520 ;
        RECT -183.440 9.040 -182.520 9.520 ;
        RECT -173.520 9.040 -172.600 9.520 ;
        RECT -163.600 9.040 -162.680 9.520 ;
        RECT -153.680 9.040 -152.760 9.520 ;
        RECT -143.760 9.040 -142.840 9.520 ;
        RECT -133.840 9.040 -132.920 9.520 ;
        RECT -123.920 9.040 -123.000 9.520 ;
        RECT -114.000 9.040 -113.080 9.520 ;
        RECT -104.080 9.040 -103.160 9.520 ;
        RECT -94.160 9.040 -93.240 9.520 ;
        RECT -84.240 9.040 -83.320 9.520 ;
        RECT -74.320 9.040 -73.400 9.520 ;
        RECT -64.400 9.040 -63.480 9.520 ;
        RECT -54.480 9.040 -53.560 9.520 ;
        RECT -44.560 9.040 -43.640 9.520 ;
        RECT -34.640 9.040 -33.720 9.520 ;
        RECT -24.720 9.040 -23.800 9.520 ;
        RECT -14.800 9.040 -13.880 9.520 ;
        RECT -4.880 9.040 -3.960 9.520 ;
        RECT 5.040 9.040 5.960 9.520 ;
        RECT 14.960 9.040 15.880 9.520 ;
        RECT -289.900 6.320 -288.980 6.800 ;
        RECT -279.980 6.320 -279.080 6.800 ;
        RECT -270.060 6.320 -269.140 6.800 ;
        RECT -260.140 6.320 -259.220 6.800 ;
        RECT -250.220 6.320 -249.300 6.800 ;
        RECT -240.300 6.320 -239.380 6.800 ;
        RECT -230.380 6.320 -229.460 6.800 ;
        RECT -220.460 6.320 -219.540 6.800 ;
        RECT -210.540 6.320 -209.620 6.800 ;
        RECT -200.620 6.320 -199.700 6.800 ;
        RECT -190.700 6.320 -189.780 6.800 ;
        RECT -180.780 6.320 -179.860 6.800 ;
        RECT -170.860 6.320 -169.940 6.800 ;
        RECT -160.940 6.320 -160.020 6.800 ;
        RECT -151.020 6.320 -150.100 6.800 ;
        RECT -141.100 6.320 -140.180 6.800 ;
        RECT -131.180 6.320 -130.260 6.800 ;
        RECT -121.260 6.320 -120.340 6.800 ;
        RECT -111.340 6.320 -110.420 6.800 ;
        RECT -101.420 6.320 -100.500 6.800 ;
        RECT -91.500 6.320 -90.580 6.800 ;
        RECT -81.580 6.320 -80.660 6.800 ;
        RECT -71.660 6.320 -70.740 6.800 ;
        RECT -61.740 6.320 -60.820 6.800 ;
        RECT -51.820 6.320 -50.900 6.800 ;
        RECT -41.900 6.320 -40.980 6.800 ;
        RECT -31.980 6.320 -31.060 6.800 ;
        RECT -22.060 6.320 -21.140 6.800 ;
        RECT -12.140 6.320 -11.220 6.800 ;
        RECT -2.220 6.320 -1.300 6.800 ;
        RECT 7.700 6.320 8.620 6.800 ;
        RECT 17.620 6.320 18.540 6.800 ;
        RECT -282.480 5.340 -281.310 6.140 ;
        RECT -272.560 5.340 -271.390 6.140 ;
        RECT -262.640 5.340 -261.470 6.140 ;
        RECT -252.720 5.340 -251.550 6.140 ;
        RECT -242.800 5.340 -241.630 6.140 ;
        RECT -232.880 5.340 -231.710 6.140 ;
        RECT -222.960 5.340 -221.790 6.140 ;
        RECT -213.040 5.340 -211.870 6.140 ;
        RECT -203.120 5.340 -201.950 6.140 ;
        RECT -193.200 5.340 -192.030 6.140 ;
        RECT -183.280 5.340 -182.110 6.140 ;
        RECT -173.360 5.340 -172.190 6.140 ;
        RECT -163.440 5.340 -162.270 6.140 ;
        RECT -153.520 5.340 -152.350 6.140 ;
        RECT -143.600 5.340 -142.430 6.140 ;
        RECT -133.680 5.340 -132.510 6.140 ;
        RECT -123.760 5.340 -122.590 6.140 ;
        RECT -113.840 5.340 -112.670 6.140 ;
        RECT -103.920 5.340 -102.750 6.140 ;
        RECT -94.000 5.340 -92.830 6.140 ;
        RECT -84.080 5.340 -82.910 6.140 ;
        RECT -74.160 5.340 -72.990 6.140 ;
        RECT -64.240 5.340 -63.070 6.140 ;
        RECT -54.320 5.340 -53.150 6.140 ;
        RECT -44.400 5.340 -43.230 6.140 ;
        RECT -34.480 5.340 -33.310 6.140 ;
        RECT -24.560 5.340 -23.390 6.140 ;
        RECT -14.640 5.340 -13.470 6.140 ;
        RECT -4.720 5.340 -3.550 6.140 ;
        RECT 5.200 5.340 6.370 6.140 ;
        RECT 15.120 5.340 16.290 6.140 ;
        RECT -289.940 -79.240 -288.770 -78.440 ;
        RECT -280.020 -79.240 -278.850 -78.440 ;
        RECT -270.100 -79.240 -268.930 -78.440 ;
        RECT -260.180 -79.240 -259.010 -78.440 ;
        RECT -250.260 -79.240 -249.090 -78.440 ;
        RECT -240.340 -79.240 -239.170 -78.440 ;
        RECT -230.420 -79.240 -229.250 -78.440 ;
        RECT -220.500 -79.240 -219.330 -78.440 ;
        RECT -210.580 -79.240 -209.410 -78.440 ;
        RECT -200.660 -79.240 -199.490 -78.440 ;
        RECT -190.740 -79.240 -189.570 -78.440 ;
        RECT -180.820 -79.240 -179.650 -78.440 ;
        RECT -170.900 -79.240 -169.730 -78.440 ;
        RECT -160.980 -79.240 -159.810 -78.440 ;
        RECT -151.060 -79.240 -149.890 -78.440 ;
        RECT -141.140 -79.240 -139.970 -78.440 ;
        RECT -131.220 -79.240 -130.050 -78.440 ;
        RECT -121.300 -79.240 -120.130 -78.440 ;
        RECT -111.380 -79.240 -110.210 -78.440 ;
        RECT -101.460 -79.240 -100.290 -78.440 ;
        RECT -91.540 -79.240 -90.370 -78.440 ;
        RECT -81.620 -79.240 -80.450 -78.440 ;
        RECT -71.700 -79.240 -70.530 -78.440 ;
        RECT -61.780 -79.240 -60.610 -78.440 ;
        RECT -51.860 -79.240 -50.690 -78.440 ;
        RECT -41.940 -79.240 -40.770 -78.440 ;
        RECT -32.020 -79.240 -30.850 -78.440 ;
        RECT -22.100 -79.240 -20.930 -78.440 ;
        RECT -12.180 -79.240 -11.010 -78.440 ;
        RECT -2.260 -79.240 -1.090 -78.440 ;
        RECT 7.660 -79.240 8.830 -78.440 ;
        RECT 17.580 -79.240 18.750 -78.440 ;
        RECT -282.280 -79.910 -281.360 -79.430 ;
        RECT -272.360 -79.910 -271.440 -79.430 ;
        RECT -262.440 -79.910 -261.520 -79.430 ;
        RECT -252.520 -79.910 -251.600 -79.430 ;
        RECT -242.600 -79.910 -241.680 -79.430 ;
        RECT -232.680 -79.910 -231.760 -79.430 ;
        RECT -222.760 -79.910 -221.840 -79.430 ;
        RECT -212.840 -79.910 -211.920 -79.430 ;
        RECT -202.920 -79.910 -202.000 -79.430 ;
        RECT -193.000 -79.910 -192.080 -79.430 ;
        RECT -183.080 -79.910 -182.160 -79.430 ;
        RECT -173.160 -79.910 -172.240 -79.430 ;
        RECT -163.240 -79.910 -162.320 -79.430 ;
        RECT -153.320 -79.910 -152.400 -79.430 ;
        RECT -143.400 -79.910 -142.480 -79.430 ;
        RECT -133.480 -79.910 -132.560 -79.430 ;
        RECT -123.560 -79.910 -122.640 -79.430 ;
        RECT -113.640 -79.910 -112.720 -79.430 ;
        RECT -103.720 -79.910 -102.800 -79.430 ;
        RECT -93.800 -79.910 -92.880 -79.430 ;
        RECT -83.880 -79.910 -82.960 -79.430 ;
        RECT -73.960 -79.910 -73.040 -79.430 ;
        RECT -64.040 -79.910 -63.120 -79.430 ;
        RECT -54.120 -79.910 -53.200 -79.430 ;
        RECT -44.200 -79.910 -43.280 -79.430 ;
        RECT -34.280 -79.910 -33.360 -79.430 ;
        RECT -24.360 -79.910 -23.440 -79.430 ;
        RECT -14.440 -79.910 -13.520 -79.430 ;
        RECT -4.520 -79.910 -3.600 -79.430 ;
        RECT 5.400 -79.910 6.320 -79.430 ;
        RECT 15.320 -79.910 16.240 -79.430 ;
        RECT -289.540 -82.630 -288.620 -82.150 ;
        RECT -279.620 -82.630 -278.720 -82.150 ;
        RECT -269.700 -82.630 -268.780 -82.150 ;
        RECT -259.780 -82.630 -258.860 -82.150 ;
        RECT -249.860 -82.630 -248.940 -82.150 ;
        RECT -239.940 -82.630 -239.020 -82.150 ;
        RECT -230.020 -82.630 -229.100 -82.150 ;
        RECT -220.100 -82.630 -219.180 -82.150 ;
        RECT -210.180 -82.630 -209.260 -82.150 ;
        RECT -200.260 -82.630 -199.340 -82.150 ;
        RECT -190.340 -82.630 -189.420 -82.150 ;
        RECT -180.420 -82.630 -179.500 -82.150 ;
        RECT -170.500 -82.630 -169.580 -82.150 ;
        RECT -160.580 -82.630 -159.660 -82.150 ;
        RECT -150.660 -82.630 -149.740 -82.150 ;
        RECT -140.740 -82.630 -139.820 -82.150 ;
        RECT -130.820 -82.630 -129.900 -82.150 ;
        RECT -120.900 -82.630 -119.980 -82.150 ;
        RECT -110.980 -82.630 -110.060 -82.150 ;
        RECT -101.060 -82.630 -100.140 -82.150 ;
        RECT -91.140 -82.630 -90.220 -82.150 ;
        RECT -81.220 -82.630 -80.300 -82.150 ;
        RECT -71.300 -82.630 -70.380 -82.150 ;
        RECT -61.380 -82.630 -60.460 -82.150 ;
        RECT -51.460 -82.630 -50.540 -82.150 ;
        RECT -41.540 -82.630 -40.620 -82.150 ;
        RECT -31.620 -82.630 -30.700 -82.150 ;
        RECT -21.700 -82.630 -20.780 -82.150 ;
        RECT -11.780 -82.630 -10.860 -82.150 ;
        RECT -1.860 -82.630 -0.940 -82.150 ;
        RECT 8.060 -82.630 8.980 -82.150 ;
        RECT 17.980 -82.630 18.900 -82.150 ;
        RECT -282.120 -83.610 -280.950 -82.810 ;
        RECT -272.200 -83.610 -271.030 -82.810 ;
        RECT -262.280 -83.610 -261.110 -82.810 ;
        RECT -252.360 -83.610 -251.190 -82.810 ;
        RECT -242.440 -83.610 -241.270 -82.810 ;
        RECT -232.520 -83.610 -231.350 -82.810 ;
        RECT -222.600 -83.610 -221.430 -82.810 ;
        RECT -212.680 -83.610 -211.510 -82.810 ;
        RECT -202.760 -83.610 -201.590 -82.810 ;
        RECT -192.840 -83.610 -191.670 -82.810 ;
        RECT -182.920 -83.610 -181.750 -82.810 ;
        RECT -173.000 -83.610 -171.830 -82.810 ;
        RECT -163.080 -83.610 -161.910 -82.810 ;
        RECT -153.160 -83.610 -151.990 -82.810 ;
        RECT -143.240 -83.610 -142.070 -82.810 ;
        RECT -133.320 -83.610 -132.150 -82.810 ;
        RECT -123.400 -83.610 -122.230 -82.810 ;
        RECT -113.480 -83.610 -112.310 -82.810 ;
        RECT -103.560 -83.610 -102.390 -82.810 ;
        RECT -93.640 -83.610 -92.470 -82.810 ;
        RECT -83.720 -83.610 -82.550 -82.810 ;
        RECT -73.800 -83.610 -72.630 -82.810 ;
        RECT -63.880 -83.610 -62.710 -82.810 ;
        RECT -53.960 -83.610 -52.790 -82.810 ;
        RECT -44.040 -83.610 -42.870 -82.810 ;
        RECT -34.120 -83.610 -32.950 -82.810 ;
        RECT -24.200 -83.610 -23.030 -82.810 ;
        RECT -14.280 -83.610 -13.110 -82.810 ;
        RECT -4.360 -83.610 -3.190 -82.810 ;
        RECT 5.560 -83.610 6.730 -82.810 ;
        RECT 15.480 -83.610 16.650 -82.810 ;
        RECT -291.700 -173.820 -290.530 -173.020 ;
        RECT -281.780 -173.820 -280.610 -173.020 ;
        RECT -271.860 -173.820 -270.690 -173.020 ;
        RECT -261.940 -173.820 -260.770 -173.020 ;
        RECT -252.020 -173.820 -250.850 -173.020 ;
        RECT -242.100 -173.820 -240.930 -173.020 ;
        RECT -232.180 -173.820 -231.010 -173.020 ;
        RECT -222.260 -173.820 -221.090 -173.020 ;
        RECT -212.340 -173.820 -211.170 -173.020 ;
        RECT -202.420 -173.820 -201.250 -173.020 ;
        RECT -192.500 -173.820 -191.330 -173.020 ;
        RECT -182.580 -173.820 -181.410 -173.020 ;
        RECT -172.660 -173.820 -171.490 -173.020 ;
        RECT -162.740 -173.820 -161.570 -173.020 ;
        RECT -152.820 -173.820 -151.650 -173.020 ;
        RECT -142.900 -173.820 -141.730 -173.020 ;
        RECT -132.980 -173.820 -131.810 -173.020 ;
        RECT -123.060 -173.820 -121.890 -173.020 ;
        RECT -113.140 -173.820 -111.970 -173.020 ;
        RECT -103.220 -173.820 -102.050 -173.020 ;
        RECT -93.300 -173.820 -92.130 -173.020 ;
        RECT -83.380 -173.820 -82.210 -173.020 ;
        RECT -73.460 -173.820 -72.290 -173.020 ;
        RECT -63.540 -173.820 -62.370 -173.020 ;
        RECT -53.620 -173.820 -52.450 -173.020 ;
        RECT -43.700 -173.820 -42.530 -173.020 ;
        RECT -33.780 -173.820 -32.610 -173.020 ;
        RECT -23.860 -173.820 -22.690 -173.020 ;
        RECT -13.940 -173.820 -12.770 -173.020 ;
        RECT -4.020 -173.820 -2.850 -173.020 ;
        RECT 5.900 -173.820 7.070 -173.020 ;
        RECT 15.820 -173.820 16.990 -173.020 ;
        RECT -284.040 -174.490 -283.120 -174.010 ;
        RECT -274.120 -174.490 -273.200 -174.010 ;
        RECT -264.200 -174.490 -263.280 -174.010 ;
        RECT -254.280 -174.490 -253.360 -174.010 ;
        RECT -244.360 -174.490 -243.440 -174.010 ;
        RECT -234.440 -174.490 -233.520 -174.010 ;
        RECT -224.520 -174.490 -223.600 -174.010 ;
        RECT -214.600 -174.490 -213.680 -174.010 ;
        RECT -204.680 -174.490 -203.760 -174.010 ;
        RECT -194.760 -174.490 -193.840 -174.010 ;
        RECT -184.840 -174.490 -183.920 -174.010 ;
        RECT -174.920 -174.490 -174.000 -174.010 ;
        RECT -165.000 -174.490 -164.080 -174.010 ;
        RECT -155.080 -174.490 -154.160 -174.010 ;
        RECT -145.160 -174.490 -144.240 -174.010 ;
        RECT -135.240 -174.490 -134.320 -174.010 ;
        RECT -125.320 -174.490 -124.400 -174.010 ;
        RECT -115.400 -174.490 -114.480 -174.010 ;
        RECT -105.480 -174.490 -104.560 -174.010 ;
        RECT -95.560 -174.490 -94.640 -174.010 ;
        RECT -85.640 -174.490 -84.720 -174.010 ;
        RECT -75.720 -174.490 -74.800 -174.010 ;
        RECT -65.800 -174.490 -64.880 -174.010 ;
        RECT -55.880 -174.490 -54.960 -174.010 ;
        RECT -45.960 -174.490 -45.040 -174.010 ;
        RECT -36.040 -174.490 -35.120 -174.010 ;
        RECT -26.120 -174.490 -25.200 -174.010 ;
        RECT -16.200 -174.490 -15.280 -174.010 ;
        RECT -6.280 -174.490 -5.360 -174.010 ;
        RECT 3.640 -174.490 4.560 -174.010 ;
        RECT 13.560 -174.490 14.480 -174.010 ;
        RECT -291.300 -177.210 -290.380 -176.730 ;
        RECT -281.380 -177.210 -280.480 -176.730 ;
        RECT -271.460 -177.210 -270.540 -176.730 ;
        RECT -261.540 -177.210 -260.620 -176.730 ;
        RECT -251.620 -177.210 -250.700 -176.730 ;
        RECT -241.700 -177.210 -240.780 -176.730 ;
        RECT -231.780 -177.210 -230.860 -176.730 ;
        RECT -221.860 -177.210 -220.940 -176.730 ;
        RECT -211.940 -177.210 -211.020 -176.730 ;
        RECT -202.020 -177.210 -201.100 -176.730 ;
        RECT -192.100 -177.210 -191.180 -176.730 ;
        RECT -182.180 -177.210 -181.260 -176.730 ;
        RECT -172.260 -177.210 -171.340 -176.730 ;
        RECT -162.340 -177.210 -161.420 -176.730 ;
        RECT -152.420 -177.210 -151.500 -176.730 ;
        RECT -142.500 -177.210 -141.580 -176.730 ;
        RECT -132.580 -177.210 -131.660 -176.730 ;
        RECT -122.660 -177.210 -121.740 -176.730 ;
        RECT -112.740 -177.210 -111.820 -176.730 ;
        RECT -102.820 -177.210 -101.900 -176.730 ;
        RECT -92.900 -177.210 -91.980 -176.730 ;
        RECT -82.980 -177.210 -82.060 -176.730 ;
        RECT -73.060 -177.210 -72.140 -176.730 ;
        RECT -63.140 -177.210 -62.220 -176.730 ;
        RECT -53.220 -177.210 -52.300 -176.730 ;
        RECT -43.300 -177.210 -42.380 -176.730 ;
        RECT -33.380 -177.210 -32.460 -176.730 ;
        RECT -23.460 -177.210 -22.540 -176.730 ;
        RECT -13.540 -177.210 -12.620 -176.730 ;
        RECT -3.620 -177.210 -2.700 -176.730 ;
        RECT 6.300 -177.210 7.220 -176.730 ;
        RECT 16.220 -177.210 17.140 -176.730 ;
        RECT -283.880 -178.190 -282.710 -177.390 ;
        RECT -273.960 -178.190 -272.790 -177.390 ;
        RECT -264.040 -178.190 -262.870 -177.390 ;
        RECT -254.120 -178.190 -252.950 -177.390 ;
        RECT -244.200 -178.190 -243.030 -177.390 ;
        RECT -234.280 -178.190 -233.110 -177.390 ;
        RECT -224.360 -178.190 -223.190 -177.390 ;
        RECT -214.440 -178.190 -213.270 -177.390 ;
        RECT -204.520 -178.190 -203.350 -177.390 ;
        RECT -194.600 -178.190 -193.430 -177.390 ;
        RECT -184.680 -178.190 -183.510 -177.390 ;
        RECT -174.760 -178.190 -173.590 -177.390 ;
        RECT -164.840 -178.190 -163.670 -177.390 ;
        RECT -154.920 -178.190 -153.750 -177.390 ;
        RECT -145.000 -178.190 -143.830 -177.390 ;
        RECT -135.080 -178.190 -133.910 -177.390 ;
        RECT -125.160 -178.190 -123.990 -177.390 ;
        RECT -115.240 -178.190 -114.070 -177.390 ;
        RECT -105.320 -178.190 -104.150 -177.390 ;
        RECT -95.400 -178.190 -94.230 -177.390 ;
        RECT -85.480 -178.190 -84.310 -177.390 ;
        RECT -75.560 -178.190 -74.390 -177.390 ;
        RECT -65.640 -178.190 -64.470 -177.390 ;
        RECT -55.720 -178.190 -54.550 -177.390 ;
        RECT -45.800 -178.190 -44.630 -177.390 ;
        RECT -35.880 -178.190 -34.710 -177.390 ;
        RECT -25.960 -178.190 -24.790 -177.390 ;
        RECT -16.040 -178.190 -14.870 -177.390 ;
        RECT -6.120 -178.190 -4.950 -177.390 ;
        RECT 3.800 -178.190 4.970 -177.390 ;
        RECT 13.720 -178.190 14.890 -177.390 ;
      LAYER via3 ;
        RECT -287.740 94.030 -287.400 94.360 ;
        RECT -277.820 94.030 -277.480 94.360 ;
        RECT -267.900 94.030 -267.560 94.360 ;
        RECT -257.980 94.030 -257.640 94.360 ;
        RECT -248.060 94.030 -247.720 94.360 ;
        RECT -238.140 94.030 -237.800 94.360 ;
        RECT -228.220 94.030 -227.880 94.360 ;
        RECT -218.300 94.030 -217.960 94.360 ;
        RECT -208.380 94.030 -208.040 94.360 ;
        RECT -198.460 94.030 -198.120 94.360 ;
        RECT -188.540 94.030 -188.200 94.360 ;
        RECT -178.620 94.030 -178.280 94.360 ;
        RECT -168.700 94.030 -168.360 94.360 ;
        RECT -158.780 94.030 -158.440 94.360 ;
        RECT -148.860 94.030 -148.520 94.360 ;
        RECT -138.940 94.030 -138.600 94.360 ;
        RECT -129.020 94.030 -128.680 94.360 ;
        RECT -119.100 94.030 -118.760 94.360 ;
        RECT -109.180 94.030 -108.840 94.360 ;
        RECT -99.260 94.030 -98.920 94.360 ;
        RECT -89.340 94.030 -89.000 94.360 ;
        RECT -79.420 94.030 -79.080 94.360 ;
        RECT -69.500 94.030 -69.160 94.360 ;
        RECT -59.580 94.030 -59.240 94.360 ;
        RECT -49.660 94.030 -49.320 94.360 ;
        RECT -39.740 94.030 -39.400 94.360 ;
        RECT -29.820 94.030 -29.480 94.360 ;
        RECT -19.900 94.030 -19.560 94.360 ;
        RECT -9.980 94.030 -9.640 94.360 ;
        RECT -0.060 94.030 0.280 94.360 ;
        RECT 9.860 94.030 10.200 94.360 ;
        RECT 19.780 94.030 20.120 94.360 ;
        RECT -280.560 93.160 -280.220 93.490 ;
        RECT -280.090 93.160 -279.750 93.490 ;
        RECT -270.640 93.160 -270.300 93.490 ;
        RECT -270.170 93.160 -269.830 93.490 ;
        RECT -260.720 93.160 -260.380 93.490 ;
        RECT -260.250 93.160 -259.910 93.490 ;
        RECT -250.800 93.160 -250.460 93.490 ;
        RECT -250.330 93.160 -249.990 93.490 ;
        RECT -240.880 93.160 -240.540 93.490 ;
        RECT -240.410 93.160 -240.070 93.490 ;
        RECT -230.960 93.160 -230.620 93.490 ;
        RECT -230.490 93.160 -230.150 93.490 ;
        RECT -221.040 93.160 -220.700 93.490 ;
        RECT -220.570 93.160 -220.230 93.490 ;
        RECT -211.120 93.160 -210.780 93.490 ;
        RECT -210.650 93.160 -210.310 93.490 ;
        RECT -201.200 93.160 -200.860 93.490 ;
        RECT -200.730 93.160 -200.390 93.490 ;
        RECT -191.280 93.160 -190.940 93.490 ;
        RECT -190.810 93.160 -190.470 93.490 ;
        RECT -181.360 93.160 -181.020 93.490 ;
        RECT -180.890 93.160 -180.550 93.490 ;
        RECT -171.440 93.160 -171.100 93.490 ;
        RECT -170.970 93.160 -170.630 93.490 ;
        RECT -161.520 93.160 -161.180 93.490 ;
        RECT -161.050 93.160 -160.710 93.490 ;
        RECT -151.600 93.160 -151.260 93.490 ;
        RECT -151.130 93.160 -150.790 93.490 ;
        RECT -141.680 93.160 -141.340 93.490 ;
        RECT -141.210 93.160 -140.870 93.490 ;
        RECT -131.760 93.160 -131.420 93.490 ;
        RECT -131.290 93.160 -130.950 93.490 ;
        RECT -121.840 93.160 -121.500 93.490 ;
        RECT -121.370 93.160 -121.030 93.490 ;
        RECT -111.920 93.160 -111.580 93.490 ;
        RECT -111.450 93.160 -111.110 93.490 ;
        RECT -102.000 93.160 -101.660 93.490 ;
        RECT -101.530 93.160 -101.190 93.490 ;
        RECT -92.080 93.160 -91.740 93.490 ;
        RECT -91.610 93.160 -91.270 93.490 ;
        RECT -82.160 93.160 -81.820 93.490 ;
        RECT -81.690 93.160 -81.350 93.490 ;
        RECT -72.240 93.160 -71.900 93.490 ;
        RECT -71.770 93.160 -71.430 93.490 ;
        RECT -62.320 93.160 -61.980 93.490 ;
        RECT -61.850 93.160 -61.510 93.490 ;
        RECT -52.400 93.160 -52.060 93.490 ;
        RECT -51.930 93.160 -51.590 93.490 ;
        RECT -42.480 93.160 -42.140 93.490 ;
        RECT -42.010 93.160 -41.670 93.490 ;
        RECT -32.560 93.160 -32.220 93.490 ;
        RECT -32.090 93.160 -31.750 93.490 ;
        RECT -22.640 93.160 -22.300 93.490 ;
        RECT -22.170 93.160 -21.830 93.490 ;
        RECT -12.720 93.160 -12.380 93.490 ;
        RECT -12.250 93.160 -11.910 93.490 ;
        RECT -2.800 93.160 -2.460 93.490 ;
        RECT -2.330 93.160 -1.990 93.490 ;
        RECT 7.120 93.160 7.460 93.490 ;
        RECT 7.590 93.160 7.930 93.490 ;
        RECT 17.040 93.160 17.380 93.490 ;
        RECT 17.510 93.160 17.850 93.490 ;
        RECT -287.820 90.440 -287.480 90.770 ;
        RECT -287.360 90.440 -287.020 90.770 ;
        RECT -277.900 90.440 -277.560 90.770 ;
        RECT -277.440 90.440 -277.100 90.770 ;
        RECT -267.980 90.440 -267.640 90.770 ;
        RECT -267.520 90.440 -267.180 90.770 ;
        RECT -258.060 90.440 -257.720 90.770 ;
        RECT -257.600 90.440 -257.260 90.770 ;
        RECT -248.140 90.440 -247.800 90.770 ;
        RECT -247.680 90.440 -247.340 90.770 ;
        RECT -238.220 90.440 -237.880 90.770 ;
        RECT -237.760 90.440 -237.420 90.770 ;
        RECT -228.300 90.440 -227.960 90.770 ;
        RECT -227.840 90.440 -227.500 90.770 ;
        RECT -218.380 90.440 -218.040 90.770 ;
        RECT -217.920 90.440 -217.580 90.770 ;
        RECT -208.460 90.440 -208.120 90.770 ;
        RECT -208.000 90.440 -207.660 90.770 ;
        RECT -198.540 90.440 -198.200 90.770 ;
        RECT -198.080 90.440 -197.740 90.770 ;
        RECT -188.620 90.440 -188.280 90.770 ;
        RECT -188.160 90.440 -187.820 90.770 ;
        RECT -178.700 90.440 -178.360 90.770 ;
        RECT -178.240 90.440 -177.900 90.770 ;
        RECT -168.780 90.440 -168.440 90.770 ;
        RECT -168.320 90.440 -167.980 90.770 ;
        RECT -158.860 90.440 -158.520 90.770 ;
        RECT -158.400 90.440 -158.060 90.770 ;
        RECT -148.940 90.440 -148.600 90.770 ;
        RECT -148.480 90.440 -148.140 90.770 ;
        RECT -139.020 90.440 -138.680 90.770 ;
        RECT -138.560 90.440 -138.220 90.770 ;
        RECT -129.100 90.440 -128.760 90.770 ;
        RECT -128.640 90.440 -128.300 90.770 ;
        RECT -119.180 90.440 -118.840 90.770 ;
        RECT -118.720 90.440 -118.380 90.770 ;
        RECT -109.260 90.440 -108.920 90.770 ;
        RECT -108.800 90.440 -108.460 90.770 ;
        RECT -99.340 90.440 -99.000 90.770 ;
        RECT -98.880 90.440 -98.540 90.770 ;
        RECT -89.420 90.440 -89.080 90.770 ;
        RECT -88.960 90.440 -88.620 90.770 ;
        RECT -79.500 90.440 -79.160 90.770 ;
        RECT -79.040 90.440 -78.700 90.770 ;
        RECT -69.580 90.440 -69.240 90.770 ;
        RECT -69.120 90.440 -68.780 90.770 ;
        RECT -59.660 90.440 -59.320 90.770 ;
        RECT -59.200 90.440 -58.860 90.770 ;
        RECT -49.740 90.440 -49.400 90.770 ;
        RECT -49.280 90.440 -48.940 90.770 ;
        RECT -39.820 90.440 -39.480 90.770 ;
        RECT -39.360 90.440 -39.020 90.770 ;
        RECT -29.900 90.440 -29.560 90.770 ;
        RECT -29.440 90.440 -29.100 90.770 ;
        RECT -19.980 90.440 -19.640 90.770 ;
        RECT -19.520 90.440 -19.180 90.770 ;
        RECT -10.060 90.440 -9.720 90.770 ;
        RECT -9.600 90.440 -9.260 90.770 ;
        RECT -0.140 90.440 0.200 90.770 ;
        RECT 0.320 90.440 0.660 90.770 ;
        RECT 9.780 90.440 10.120 90.770 ;
        RECT 10.240 90.440 10.580 90.770 ;
        RECT 19.700 90.440 20.040 90.770 ;
        RECT 20.160 90.440 20.500 90.770 ;
        RECT -280.170 89.680 -279.830 90.010 ;
        RECT -270.250 89.680 -269.910 90.010 ;
        RECT -260.330 89.680 -259.990 90.010 ;
        RECT -250.410 89.680 -250.070 90.010 ;
        RECT -240.490 89.680 -240.150 90.010 ;
        RECT -230.570 89.680 -230.230 90.010 ;
        RECT -220.650 89.680 -220.310 90.010 ;
        RECT -210.730 89.680 -210.390 90.010 ;
        RECT -200.810 89.680 -200.470 90.010 ;
        RECT -190.890 89.680 -190.550 90.010 ;
        RECT -180.970 89.680 -180.630 90.010 ;
        RECT -171.050 89.680 -170.710 90.010 ;
        RECT -161.130 89.680 -160.790 90.010 ;
        RECT -151.210 89.680 -150.870 90.010 ;
        RECT -141.290 89.680 -140.950 90.010 ;
        RECT -131.370 89.680 -131.030 90.010 ;
        RECT -121.450 89.680 -121.110 90.010 ;
        RECT -111.530 89.680 -111.190 90.010 ;
        RECT -101.610 89.680 -101.270 90.010 ;
        RECT -91.690 89.680 -91.350 90.010 ;
        RECT -81.770 89.680 -81.430 90.010 ;
        RECT -71.850 89.680 -71.510 90.010 ;
        RECT -61.930 89.680 -61.590 90.010 ;
        RECT -52.010 89.680 -51.670 90.010 ;
        RECT -42.090 89.680 -41.750 90.010 ;
        RECT -32.170 89.680 -31.830 90.010 ;
        RECT -22.250 89.680 -21.910 90.010 ;
        RECT -12.330 89.680 -11.990 90.010 ;
        RECT -2.410 89.680 -2.070 90.010 ;
        RECT 7.510 89.680 7.850 90.010 ;
        RECT 17.430 89.680 17.770 90.010 ;
        RECT -289.760 9.980 -289.420 10.310 ;
        RECT -279.840 9.980 -279.500 10.310 ;
        RECT -269.920 9.980 -269.580 10.310 ;
        RECT -260.000 9.980 -259.660 10.310 ;
        RECT -250.080 9.980 -249.740 10.310 ;
        RECT -240.160 9.980 -239.820 10.310 ;
        RECT -230.240 9.980 -229.900 10.310 ;
        RECT -220.320 9.980 -219.980 10.310 ;
        RECT -210.400 9.980 -210.060 10.310 ;
        RECT -200.480 9.980 -200.140 10.310 ;
        RECT -190.560 9.980 -190.220 10.310 ;
        RECT -180.640 9.980 -180.300 10.310 ;
        RECT -170.720 9.980 -170.380 10.310 ;
        RECT -160.800 9.980 -160.460 10.310 ;
        RECT -150.880 9.980 -150.540 10.310 ;
        RECT -140.960 9.980 -140.620 10.310 ;
        RECT -131.040 9.980 -130.700 10.310 ;
        RECT -121.120 9.980 -120.780 10.310 ;
        RECT -111.200 9.980 -110.860 10.310 ;
        RECT -101.280 9.980 -100.940 10.310 ;
        RECT -91.360 9.980 -91.020 10.310 ;
        RECT -81.440 9.980 -81.100 10.310 ;
        RECT -71.520 9.980 -71.180 10.310 ;
        RECT -61.600 9.980 -61.260 10.310 ;
        RECT -51.680 9.980 -51.340 10.310 ;
        RECT -41.760 9.980 -41.420 10.310 ;
        RECT -31.840 9.980 -31.500 10.310 ;
        RECT -21.920 9.980 -21.580 10.310 ;
        RECT -12.000 9.980 -11.660 10.310 ;
        RECT -2.080 9.980 -1.740 10.310 ;
        RECT 7.840 9.980 8.180 10.310 ;
        RECT 17.760 9.980 18.100 10.310 ;
        RECT -282.580 9.110 -282.240 9.440 ;
        RECT -282.110 9.110 -281.770 9.440 ;
        RECT -272.660 9.110 -272.320 9.440 ;
        RECT -272.190 9.110 -271.850 9.440 ;
        RECT -262.740 9.110 -262.400 9.440 ;
        RECT -262.270 9.110 -261.930 9.440 ;
        RECT -252.820 9.110 -252.480 9.440 ;
        RECT -252.350 9.110 -252.010 9.440 ;
        RECT -242.900 9.110 -242.560 9.440 ;
        RECT -242.430 9.110 -242.090 9.440 ;
        RECT -232.980 9.110 -232.640 9.440 ;
        RECT -232.510 9.110 -232.170 9.440 ;
        RECT -223.060 9.110 -222.720 9.440 ;
        RECT -222.590 9.110 -222.250 9.440 ;
        RECT -213.140 9.110 -212.800 9.440 ;
        RECT -212.670 9.110 -212.330 9.440 ;
        RECT -203.220 9.110 -202.880 9.440 ;
        RECT -202.750 9.110 -202.410 9.440 ;
        RECT -193.300 9.110 -192.960 9.440 ;
        RECT -192.830 9.110 -192.490 9.440 ;
        RECT -183.380 9.110 -183.040 9.440 ;
        RECT -182.910 9.110 -182.570 9.440 ;
        RECT -173.460 9.110 -173.120 9.440 ;
        RECT -172.990 9.110 -172.650 9.440 ;
        RECT -163.540 9.110 -163.200 9.440 ;
        RECT -163.070 9.110 -162.730 9.440 ;
        RECT -153.620 9.110 -153.280 9.440 ;
        RECT -153.150 9.110 -152.810 9.440 ;
        RECT -143.700 9.110 -143.360 9.440 ;
        RECT -143.230 9.110 -142.890 9.440 ;
        RECT -133.780 9.110 -133.440 9.440 ;
        RECT -133.310 9.110 -132.970 9.440 ;
        RECT -123.860 9.110 -123.520 9.440 ;
        RECT -123.390 9.110 -123.050 9.440 ;
        RECT -113.940 9.110 -113.600 9.440 ;
        RECT -113.470 9.110 -113.130 9.440 ;
        RECT -104.020 9.110 -103.680 9.440 ;
        RECT -103.550 9.110 -103.210 9.440 ;
        RECT -94.100 9.110 -93.760 9.440 ;
        RECT -93.630 9.110 -93.290 9.440 ;
        RECT -84.180 9.110 -83.840 9.440 ;
        RECT -83.710 9.110 -83.370 9.440 ;
        RECT -74.260 9.110 -73.920 9.440 ;
        RECT -73.790 9.110 -73.450 9.440 ;
        RECT -64.340 9.110 -64.000 9.440 ;
        RECT -63.870 9.110 -63.530 9.440 ;
        RECT -54.420 9.110 -54.080 9.440 ;
        RECT -53.950 9.110 -53.610 9.440 ;
        RECT -44.500 9.110 -44.160 9.440 ;
        RECT -44.030 9.110 -43.690 9.440 ;
        RECT -34.580 9.110 -34.240 9.440 ;
        RECT -34.110 9.110 -33.770 9.440 ;
        RECT -24.660 9.110 -24.320 9.440 ;
        RECT -24.190 9.110 -23.850 9.440 ;
        RECT -14.740 9.110 -14.400 9.440 ;
        RECT -14.270 9.110 -13.930 9.440 ;
        RECT -4.820 9.110 -4.480 9.440 ;
        RECT -4.350 9.110 -4.010 9.440 ;
        RECT 5.100 9.110 5.440 9.440 ;
        RECT 5.570 9.110 5.910 9.440 ;
        RECT 15.020 9.110 15.360 9.440 ;
        RECT 15.490 9.110 15.830 9.440 ;
        RECT -289.840 6.390 -289.500 6.720 ;
        RECT -289.380 6.390 -289.040 6.720 ;
        RECT -279.920 6.390 -279.580 6.720 ;
        RECT -279.460 6.390 -279.120 6.720 ;
        RECT -270.000 6.390 -269.660 6.720 ;
        RECT -269.540 6.390 -269.200 6.720 ;
        RECT -260.080 6.390 -259.740 6.720 ;
        RECT -259.620 6.390 -259.280 6.720 ;
        RECT -250.160 6.390 -249.820 6.720 ;
        RECT -249.700 6.390 -249.360 6.720 ;
        RECT -240.240 6.390 -239.900 6.720 ;
        RECT -239.780 6.390 -239.440 6.720 ;
        RECT -230.320 6.390 -229.980 6.720 ;
        RECT -229.860 6.390 -229.520 6.720 ;
        RECT -220.400 6.390 -220.060 6.720 ;
        RECT -219.940 6.390 -219.600 6.720 ;
        RECT -210.480 6.390 -210.140 6.720 ;
        RECT -210.020 6.390 -209.680 6.720 ;
        RECT -200.560 6.390 -200.220 6.720 ;
        RECT -200.100 6.390 -199.760 6.720 ;
        RECT -190.640 6.390 -190.300 6.720 ;
        RECT -190.180 6.390 -189.840 6.720 ;
        RECT -180.720 6.390 -180.380 6.720 ;
        RECT -180.260 6.390 -179.920 6.720 ;
        RECT -170.800 6.390 -170.460 6.720 ;
        RECT -170.340 6.390 -170.000 6.720 ;
        RECT -160.880 6.390 -160.540 6.720 ;
        RECT -160.420 6.390 -160.080 6.720 ;
        RECT -150.960 6.390 -150.620 6.720 ;
        RECT -150.500 6.390 -150.160 6.720 ;
        RECT -141.040 6.390 -140.700 6.720 ;
        RECT -140.580 6.390 -140.240 6.720 ;
        RECT -131.120 6.390 -130.780 6.720 ;
        RECT -130.660 6.390 -130.320 6.720 ;
        RECT -121.200 6.390 -120.860 6.720 ;
        RECT -120.740 6.390 -120.400 6.720 ;
        RECT -111.280 6.390 -110.940 6.720 ;
        RECT -110.820 6.390 -110.480 6.720 ;
        RECT -101.360 6.390 -101.020 6.720 ;
        RECT -100.900 6.390 -100.560 6.720 ;
        RECT -91.440 6.390 -91.100 6.720 ;
        RECT -90.980 6.390 -90.640 6.720 ;
        RECT -81.520 6.390 -81.180 6.720 ;
        RECT -81.060 6.390 -80.720 6.720 ;
        RECT -71.600 6.390 -71.260 6.720 ;
        RECT -71.140 6.390 -70.800 6.720 ;
        RECT -61.680 6.390 -61.340 6.720 ;
        RECT -61.220 6.390 -60.880 6.720 ;
        RECT -51.760 6.390 -51.420 6.720 ;
        RECT -51.300 6.390 -50.960 6.720 ;
        RECT -41.840 6.390 -41.500 6.720 ;
        RECT -41.380 6.390 -41.040 6.720 ;
        RECT -31.920 6.390 -31.580 6.720 ;
        RECT -31.460 6.390 -31.120 6.720 ;
        RECT -22.000 6.390 -21.660 6.720 ;
        RECT -21.540 6.390 -21.200 6.720 ;
        RECT -12.080 6.390 -11.740 6.720 ;
        RECT -11.620 6.390 -11.280 6.720 ;
        RECT -2.160 6.390 -1.820 6.720 ;
        RECT -1.700 6.390 -1.360 6.720 ;
        RECT 7.760 6.390 8.100 6.720 ;
        RECT 8.220 6.390 8.560 6.720 ;
        RECT 17.680 6.390 18.020 6.720 ;
        RECT 18.140 6.390 18.480 6.720 ;
        RECT -282.190 5.630 -281.850 5.960 ;
        RECT -272.270 5.630 -271.930 5.960 ;
        RECT -262.350 5.630 -262.010 5.960 ;
        RECT -252.430 5.630 -252.090 5.960 ;
        RECT -242.510 5.630 -242.170 5.960 ;
        RECT -232.590 5.630 -232.250 5.960 ;
        RECT -222.670 5.630 -222.330 5.960 ;
        RECT -212.750 5.630 -212.410 5.960 ;
        RECT -202.830 5.630 -202.490 5.960 ;
        RECT -192.910 5.630 -192.570 5.960 ;
        RECT -182.990 5.630 -182.650 5.960 ;
        RECT -173.070 5.630 -172.730 5.960 ;
        RECT -163.150 5.630 -162.810 5.960 ;
        RECT -153.230 5.630 -152.890 5.960 ;
        RECT -143.310 5.630 -142.970 5.960 ;
        RECT -133.390 5.630 -133.050 5.960 ;
        RECT -123.470 5.630 -123.130 5.960 ;
        RECT -113.550 5.630 -113.210 5.960 ;
        RECT -103.630 5.630 -103.290 5.960 ;
        RECT -93.710 5.630 -93.370 5.960 ;
        RECT -83.790 5.630 -83.450 5.960 ;
        RECT -73.870 5.630 -73.530 5.960 ;
        RECT -63.950 5.630 -63.610 5.960 ;
        RECT -54.030 5.630 -53.690 5.960 ;
        RECT -44.110 5.630 -43.770 5.960 ;
        RECT -34.190 5.630 -33.850 5.960 ;
        RECT -24.270 5.630 -23.930 5.960 ;
        RECT -14.350 5.630 -14.010 5.960 ;
        RECT -4.430 5.630 -4.090 5.960 ;
        RECT 5.490 5.630 5.830 5.960 ;
        RECT 15.410 5.630 15.750 5.960 ;
        RECT -289.400 -78.970 -289.060 -78.640 ;
        RECT -279.480 -78.970 -279.140 -78.640 ;
        RECT -269.560 -78.970 -269.220 -78.640 ;
        RECT -259.640 -78.970 -259.300 -78.640 ;
        RECT -249.720 -78.970 -249.380 -78.640 ;
        RECT -239.800 -78.970 -239.460 -78.640 ;
        RECT -229.880 -78.970 -229.540 -78.640 ;
        RECT -219.960 -78.970 -219.620 -78.640 ;
        RECT -210.040 -78.970 -209.700 -78.640 ;
        RECT -200.120 -78.970 -199.780 -78.640 ;
        RECT -190.200 -78.970 -189.860 -78.640 ;
        RECT -180.280 -78.970 -179.940 -78.640 ;
        RECT -170.360 -78.970 -170.020 -78.640 ;
        RECT -160.440 -78.970 -160.100 -78.640 ;
        RECT -150.520 -78.970 -150.180 -78.640 ;
        RECT -140.600 -78.970 -140.260 -78.640 ;
        RECT -130.680 -78.970 -130.340 -78.640 ;
        RECT -120.760 -78.970 -120.420 -78.640 ;
        RECT -110.840 -78.970 -110.500 -78.640 ;
        RECT -100.920 -78.970 -100.580 -78.640 ;
        RECT -91.000 -78.970 -90.660 -78.640 ;
        RECT -81.080 -78.970 -80.740 -78.640 ;
        RECT -71.160 -78.970 -70.820 -78.640 ;
        RECT -61.240 -78.970 -60.900 -78.640 ;
        RECT -51.320 -78.970 -50.980 -78.640 ;
        RECT -41.400 -78.970 -41.060 -78.640 ;
        RECT -31.480 -78.970 -31.140 -78.640 ;
        RECT -21.560 -78.970 -21.220 -78.640 ;
        RECT -11.640 -78.970 -11.300 -78.640 ;
        RECT -1.720 -78.970 -1.380 -78.640 ;
        RECT 8.200 -78.970 8.540 -78.640 ;
        RECT 18.120 -78.970 18.460 -78.640 ;
        RECT -282.220 -79.840 -281.880 -79.510 ;
        RECT -281.750 -79.840 -281.410 -79.510 ;
        RECT -272.300 -79.840 -271.960 -79.510 ;
        RECT -271.830 -79.840 -271.490 -79.510 ;
        RECT -262.380 -79.840 -262.040 -79.510 ;
        RECT -261.910 -79.840 -261.570 -79.510 ;
        RECT -252.460 -79.840 -252.120 -79.510 ;
        RECT -251.990 -79.840 -251.650 -79.510 ;
        RECT -242.540 -79.840 -242.200 -79.510 ;
        RECT -242.070 -79.840 -241.730 -79.510 ;
        RECT -232.620 -79.840 -232.280 -79.510 ;
        RECT -232.150 -79.840 -231.810 -79.510 ;
        RECT -222.700 -79.840 -222.360 -79.510 ;
        RECT -222.230 -79.840 -221.890 -79.510 ;
        RECT -212.780 -79.840 -212.440 -79.510 ;
        RECT -212.310 -79.840 -211.970 -79.510 ;
        RECT -202.860 -79.840 -202.520 -79.510 ;
        RECT -202.390 -79.840 -202.050 -79.510 ;
        RECT -192.940 -79.840 -192.600 -79.510 ;
        RECT -192.470 -79.840 -192.130 -79.510 ;
        RECT -183.020 -79.840 -182.680 -79.510 ;
        RECT -182.550 -79.840 -182.210 -79.510 ;
        RECT -173.100 -79.840 -172.760 -79.510 ;
        RECT -172.630 -79.840 -172.290 -79.510 ;
        RECT -163.180 -79.840 -162.840 -79.510 ;
        RECT -162.710 -79.840 -162.370 -79.510 ;
        RECT -153.260 -79.840 -152.920 -79.510 ;
        RECT -152.790 -79.840 -152.450 -79.510 ;
        RECT -143.340 -79.840 -143.000 -79.510 ;
        RECT -142.870 -79.840 -142.530 -79.510 ;
        RECT -133.420 -79.840 -133.080 -79.510 ;
        RECT -132.950 -79.840 -132.610 -79.510 ;
        RECT -123.500 -79.840 -123.160 -79.510 ;
        RECT -123.030 -79.840 -122.690 -79.510 ;
        RECT -113.580 -79.840 -113.240 -79.510 ;
        RECT -113.110 -79.840 -112.770 -79.510 ;
        RECT -103.660 -79.840 -103.320 -79.510 ;
        RECT -103.190 -79.840 -102.850 -79.510 ;
        RECT -93.740 -79.840 -93.400 -79.510 ;
        RECT -93.270 -79.840 -92.930 -79.510 ;
        RECT -83.820 -79.840 -83.480 -79.510 ;
        RECT -83.350 -79.840 -83.010 -79.510 ;
        RECT -73.900 -79.840 -73.560 -79.510 ;
        RECT -73.430 -79.840 -73.090 -79.510 ;
        RECT -63.980 -79.840 -63.640 -79.510 ;
        RECT -63.510 -79.840 -63.170 -79.510 ;
        RECT -54.060 -79.840 -53.720 -79.510 ;
        RECT -53.590 -79.840 -53.250 -79.510 ;
        RECT -44.140 -79.840 -43.800 -79.510 ;
        RECT -43.670 -79.840 -43.330 -79.510 ;
        RECT -34.220 -79.840 -33.880 -79.510 ;
        RECT -33.750 -79.840 -33.410 -79.510 ;
        RECT -24.300 -79.840 -23.960 -79.510 ;
        RECT -23.830 -79.840 -23.490 -79.510 ;
        RECT -14.380 -79.840 -14.040 -79.510 ;
        RECT -13.910 -79.840 -13.570 -79.510 ;
        RECT -4.460 -79.840 -4.120 -79.510 ;
        RECT -3.990 -79.840 -3.650 -79.510 ;
        RECT 5.460 -79.840 5.800 -79.510 ;
        RECT 5.930 -79.840 6.270 -79.510 ;
        RECT 15.380 -79.840 15.720 -79.510 ;
        RECT 15.850 -79.840 16.190 -79.510 ;
        RECT -289.480 -82.560 -289.140 -82.230 ;
        RECT -289.020 -82.560 -288.680 -82.230 ;
        RECT -279.560 -82.560 -279.220 -82.230 ;
        RECT -279.100 -82.560 -278.760 -82.230 ;
        RECT -269.640 -82.560 -269.300 -82.230 ;
        RECT -269.180 -82.560 -268.840 -82.230 ;
        RECT -259.720 -82.560 -259.380 -82.230 ;
        RECT -259.260 -82.560 -258.920 -82.230 ;
        RECT -249.800 -82.560 -249.460 -82.230 ;
        RECT -249.340 -82.560 -249.000 -82.230 ;
        RECT -239.880 -82.560 -239.540 -82.230 ;
        RECT -239.420 -82.560 -239.080 -82.230 ;
        RECT -229.960 -82.560 -229.620 -82.230 ;
        RECT -229.500 -82.560 -229.160 -82.230 ;
        RECT -220.040 -82.560 -219.700 -82.230 ;
        RECT -219.580 -82.560 -219.240 -82.230 ;
        RECT -210.120 -82.560 -209.780 -82.230 ;
        RECT -209.660 -82.560 -209.320 -82.230 ;
        RECT -200.200 -82.560 -199.860 -82.230 ;
        RECT -199.740 -82.560 -199.400 -82.230 ;
        RECT -190.280 -82.560 -189.940 -82.230 ;
        RECT -189.820 -82.560 -189.480 -82.230 ;
        RECT -180.360 -82.560 -180.020 -82.230 ;
        RECT -179.900 -82.560 -179.560 -82.230 ;
        RECT -170.440 -82.560 -170.100 -82.230 ;
        RECT -169.980 -82.560 -169.640 -82.230 ;
        RECT -160.520 -82.560 -160.180 -82.230 ;
        RECT -160.060 -82.560 -159.720 -82.230 ;
        RECT -150.600 -82.560 -150.260 -82.230 ;
        RECT -150.140 -82.560 -149.800 -82.230 ;
        RECT -140.680 -82.560 -140.340 -82.230 ;
        RECT -140.220 -82.560 -139.880 -82.230 ;
        RECT -130.760 -82.560 -130.420 -82.230 ;
        RECT -130.300 -82.560 -129.960 -82.230 ;
        RECT -120.840 -82.560 -120.500 -82.230 ;
        RECT -120.380 -82.560 -120.040 -82.230 ;
        RECT -110.920 -82.560 -110.580 -82.230 ;
        RECT -110.460 -82.560 -110.120 -82.230 ;
        RECT -101.000 -82.560 -100.660 -82.230 ;
        RECT -100.540 -82.560 -100.200 -82.230 ;
        RECT -91.080 -82.560 -90.740 -82.230 ;
        RECT -90.620 -82.560 -90.280 -82.230 ;
        RECT -81.160 -82.560 -80.820 -82.230 ;
        RECT -80.700 -82.560 -80.360 -82.230 ;
        RECT -71.240 -82.560 -70.900 -82.230 ;
        RECT -70.780 -82.560 -70.440 -82.230 ;
        RECT -61.320 -82.560 -60.980 -82.230 ;
        RECT -60.860 -82.560 -60.520 -82.230 ;
        RECT -51.400 -82.560 -51.060 -82.230 ;
        RECT -50.940 -82.560 -50.600 -82.230 ;
        RECT -41.480 -82.560 -41.140 -82.230 ;
        RECT -41.020 -82.560 -40.680 -82.230 ;
        RECT -31.560 -82.560 -31.220 -82.230 ;
        RECT -31.100 -82.560 -30.760 -82.230 ;
        RECT -21.640 -82.560 -21.300 -82.230 ;
        RECT -21.180 -82.560 -20.840 -82.230 ;
        RECT -11.720 -82.560 -11.380 -82.230 ;
        RECT -11.260 -82.560 -10.920 -82.230 ;
        RECT -1.800 -82.560 -1.460 -82.230 ;
        RECT -1.340 -82.560 -1.000 -82.230 ;
        RECT 8.120 -82.560 8.460 -82.230 ;
        RECT 8.580 -82.560 8.920 -82.230 ;
        RECT 18.040 -82.560 18.380 -82.230 ;
        RECT 18.500 -82.560 18.840 -82.230 ;
        RECT -281.830 -83.320 -281.490 -82.990 ;
        RECT -271.910 -83.320 -271.570 -82.990 ;
        RECT -261.990 -83.320 -261.650 -82.990 ;
        RECT -252.070 -83.320 -251.730 -82.990 ;
        RECT -242.150 -83.320 -241.810 -82.990 ;
        RECT -232.230 -83.320 -231.890 -82.990 ;
        RECT -222.310 -83.320 -221.970 -82.990 ;
        RECT -212.390 -83.320 -212.050 -82.990 ;
        RECT -202.470 -83.320 -202.130 -82.990 ;
        RECT -192.550 -83.320 -192.210 -82.990 ;
        RECT -182.630 -83.320 -182.290 -82.990 ;
        RECT -172.710 -83.320 -172.370 -82.990 ;
        RECT -162.790 -83.320 -162.450 -82.990 ;
        RECT -152.870 -83.320 -152.530 -82.990 ;
        RECT -142.950 -83.320 -142.610 -82.990 ;
        RECT -133.030 -83.320 -132.690 -82.990 ;
        RECT -123.110 -83.320 -122.770 -82.990 ;
        RECT -113.190 -83.320 -112.850 -82.990 ;
        RECT -103.270 -83.320 -102.930 -82.990 ;
        RECT -93.350 -83.320 -93.010 -82.990 ;
        RECT -83.430 -83.320 -83.090 -82.990 ;
        RECT -73.510 -83.320 -73.170 -82.990 ;
        RECT -63.590 -83.320 -63.250 -82.990 ;
        RECT -53.670 -83.320 -53.330 -82.990 ;
        RECT -43.750 -83.320 -43.410 -82.990 ;
        RECT -33.830 -83.320 -33.490 -82.990 ;
        RECT -23.910 -83.320 -23.570 -82.990 ;
        RECT -13.990 -83.320 -13.650 -82.990 ;
        RECT -4.070 -83.320 -3.730 -82.990 ;
        RECT 5.850 -83.320 6.190 -82.990 ;
        RECT 15.770 -83.320 16.110 -82.990 ;
        RECT -291.160 -173.550 -290.820 -173.220 ;
        RECT -281.240 -173.550 -280.900 -173.220 ;
        RECT -271.320 -173.550 -270.980 -173.220 ;
        RECT -261.400 -173.550 -261.060 -173.220 ;
        RECT -251.480 -173.550 -251.140 -173.220 ;
        RECT -241.560 -173.550 -241.220 -173.220 ;
        RECT -231.640 -173.550 -231.300 -173.220 ;
        RECT -221.720 -173.550 -221.380 -173.220 ;
        RECT -211.800 -173.550 -211.460 -173.220 ;
        RECT -201.880 -173.550 -201.540 -173.220 ;
        RECT -191.960 -173.550 -191.620 -173.220 ;
        RECT -182.040 -173.550 -181.700 -173.220 ;
        RECT -172.120 -173.550 -171.780 -173.220 ;
        RECT -162.200 -173.550 -161.860 -173.220 ;
        RECT -152.280 -173.550 -151.940 -173.220 ;
        RECT -142.360 -173.550 -142.020 -173.220 ;
        RECT -132.440 -173.550 -132.100 -173.220 ;
        RECT -122.520 -173.550 -122.180 -173.220 ;
        RECT -112.600 -173.550 -112.260 -173.220 ;
        RECT -102.680 -173.550 -102.340 -173.220 ;
        RECT -92.760 -173.550 -92.420 -173.220 ;
        RECT -82.840 -173.550 -82.500 -173.220 ;
        RECT -72.920 -173.550 -72.580 -173.220 ;
        RECT -63.000 -173.550 -62.660 -173.220 ;
        RECT -53.080 -173.550 -52.740 -173.220 ;
        RECT -43.160 -173.550 -42.820 -173.220 ;
        RECT -33.240 -173.550 -32.900 -173.220 ;
        RECT -23.320 -173.550 -22.980 -173.220 ;
        RECT -13.400 -173.550 -13.060 -173.220 ;
        RECT -3.480 -173.550 -3.140 -173.220 ;
        RECT 6.440 -173.550 6.780 -173.220 ;
        RECT 16.360 -173.550 16.700 -173.220 ;
        RECT -283.980 -174.420 -283.640 -174.090 ;
        RECT -283.510 -174.420 -283.170 -174.090 ;
        RECT -274.060 -174.420 -273.720 -174.090 ;
        RECT -273.590 -174.420 -273.250 -174.090 ;
        RECT -264.140 -174.420 -263.800 -174.090 ;
        RECT -263.670 -174.420 -263.330 -174.090 ;
        RECT -254.220 -174.420 -253.880 -174.090 ;
        RECT -253.750 -174.420 -253.410 -174.090 ;
        RECT -244.300 -174.420 -243.960 -174.090 ;
        RECT -243.830 -174.420 -243.490 -174.090 ;
        RECT -234.380 -174.420 -234.040 -174.090 ;
        RECT -233.910 -174.420 -233.570 -174.090 ;
        RECT -224.460 -174.420 -224.120 -174.090 ;
        RECT -223.990 -174.420 -223.650 -174.090 ;
        RECT -214.540 -174.420 -214.200 -174.090 ;
        RECT -214.070 -174.420 -213.730 -174.090 ;
        RECT -204.620 -174.420 -204.280 -174.090 ;
        RECT -204.150 -174.420 -203.810 -174.090 ;
        RECT -194.700 -174.420 -194.360 -174.090 ;
        RECT -194.230 -174.420 -193.890 -174.090 ;
        RECT -184.780 -174.420 -184.440 -174.090 ;
        RECT -184.310 -174.420 -183.970 -174.090 ;
        RECT -174.860 -174.420 -174.520 -174.090 ;
        RECT -174.390 -174.420 -174.050 -174.090 ;
        RECT -164.940 -174.420 -164.600 -174.090 ;
        RECT -164.470 -174.420 -164.130 -174.090 ;
        RECT -155.020 -174.420 -154.680 -174.090 ;
        RECT -154.550 -174.420 -154.210 -174.090 ;
        RECT -145.100 -174.420 -144.760 -174.090 ;
        RECT -144.630 -174.420 -144.290 -174.090 ;
        RECT -135.180 -174.420 -134.840 -174.090 ;
        RECT -134.710 -174.420 -134.370 -174.090 ;
        RECT -125.260 -174.420 -124.920 -174.090 ;
        RECT -124.790 -174.420 -124.450 -174.090 ;
        RECT -115.340 -174.420 -115.000 -174.090 ;
        RECT -114.870 -174.420 -114.530 -174.090 ;
        RECT -105.420 -174.420 -105.080 -174.090 ;
        RECT -104.950 -174.420 -104.610 -174.090 ;
        RECT -95.500 -174.420 -95.160 -174.090 ;
        RECT -95.030 -174.420 -94.690 -174.090 ;
        RECT -85.580 -174.420 -85.240 -174.090 ;
        RECT -85.110 -174.420 -84.770 -174.090 ;
        RECT -75.660 -174.420 -75.320 -174.090 ;
        RECT -75.190 -174.420 -74.850 -174.090 ;
        RECT -65.740 -174.420 -65.400 -174.090 ;
        RECT -65.270 -174.420 -64.930 -174.090 ;
        RECT -55.820 -174.420 -55.480 -174.090 ;
        RECT -55.350 -174.420 -55.010 -174.090 ;
        RECT -45.900 -174.420 -45.560 -174.090 ;
        RECT -45.430 -174.420 -45.090 -174.090 ;
        RECT -35.980 -174.420 -35.640 -174.090 ;
        RECT -35.510 -174.420 -35.170 -174.090 ;
        RECT -26.060 -174.420 -25.720 -174.090 ;
        RECT -25.590 -174.420 -25.250 -174.090 ;
        RECT -16.140 -174.420 -15.800 -174.090 ;
        RECT -15.670 -174.420 -15.330 -174.090 ;
        RECT -6.220 -174.420 -5.880 -174.090 ;
        RECT -5.750 -174.420 -5.410 -174.090 ;
        RECT 3.700 -174.420 4.040 -174.090 ;
        RECT 4.170 -174.420 4.510 -174.090 ;
        RECT 13.620 -174.420 13.960 -174.090 ;
        RECT 14.090 -174.420 14.430 -174.090 ;
        RECT -291.240 -177.140 -290.900 -176.810 ;
        RECT -290.780 -177.140 -290.440 -176.810 ;
        RECT -281.320 -177.140 -280.980 -176.810 ;
        RECT -280.860 -177.140 -280.520 -176.810 ;
        RECT -271.400 -177.140 -271.060 -176.810 ;
        RECT -270.940 -177.140 -270.600 -176.810 ;
        RECT -261.480 -177.140 -261.140 -176.810 ;
        RECT -261.020 -177.140 -260.680 -176.810 ;
        RECT -251.560 -177.140 -251.220 -176.810 ;
        RECT -251.100 -177.140 -250.760 -176.810 ;
        RECT -241.640 -177.140 -241.300 -176.810 ;
        RECT -241.180 -177.140 -240.840 -176.810 ;
        RECT -231.720 -177.140 -231.380 -176.810 ;
        RECT -231.260 -177.140 -230.920 -176.810 ;
        RECT -221.800 -177.140 -221.460 -176.810 ;
        RECT -221.340 -177.140 -221.000 -176.810 ;
        RECT -211.880 -177.140 -211.540 -176.810 ;
        RECT -211.420 -177.140 -211.080 -176.810 ;
        RECT -201.960 -177.140 -201.620 -176.810 ;
        RECT -201.500 -177.140 -201.160 -176.810 ;
        RECT -192.040 -177.140 -191.700 -176.810 ;
        RECT -191.580 -177.140 -191.240 -176.810 ;
        RECT -182.120 -177.140 -181.780 -176.810 ;
        RECT -181.660 -177.140 -181.320 -176.810 ;
        RECT -172.200 -177.140 -171.860 -176.810 ;
        RECT -171.740 -177.140 -171.400 -176.810 ;
        RECT -162.280 -177.140 -161.940 -176.810 ;
        RECT -161.820 -177.140 -161.480 -176.810 ;
        RECT -152.360 -177.140 -152.020 -176.810 ;
        RECT -151.900 -177.140 -151.560 -176.810 ;
        RECT -142.440 -177.140 -142.100 -176.810 ;
        RECT -141.980 -177.140 -141.640 -176.810 ;
        RECT -132.520 -177.140 -132.180 -176.810 ;
        RECT -132.060 -177.140 -131.720 -176.810 ;
        RECT -122.600 -177.140 -122.260 -176.810 ;
        RECT -122.140 -177.140 -121.800 -176.810 ;
        RECT -112.680 -177.140 -112.340 -176.810 ;
        RECT -112.220 -177.140 -111.880 -176.810 ;
        RECT -102.760 -177.140 -102.420 -176.810 ;
        RECT -102.300 -177.140 -101.960 -176.810 ;
        RECT -92.840 -177.140 -92.500 -176.810 ;
        RECT -92.380 -177.140 -92.040 -176.810 ;
        RECT -82.920 -177.140 -82.580 -176.810 ;
        RECT -82.460 -177.140 -82.120 -176.810 ;
        RECT -73.000 -177.140 -72.660 -176.810 ;
        RECT -72.540 -177.140 -72.200 -176.810 ;
        RECT -63.080 -177.140 -62.740 -176.810 ;
        RECT -62.620 -177.140 -62.280 -176.810 ;
        RECT -53.160 -177.140 -52.820 -176.810 ;
        RECT -52.700 -177.140 -52.360 -176.810 ;
        RECT -43.240 -177.140 -42.900 -176.810 ;
        RECT -42.780 -177.140 -42.440 -176.810 ;
        RECT -33.320 -177.140 -32.980 -176.810 ;
        RECT -32.860 -177.140 -32.520 -176.810 ;
        RECT -23.400 -177.140 -23.060 -176.810 ;
        RECT -22.940 -177.140 -22.600 -176.810 ;
        RECT -13.480 -177.140 -13.140 -176.810 ;
        RECT -13.020 -177.140 -12.680 -176.810 ;
        RECT -3.560 -177.140 -3.220 -176.810 ;
        RECT -3.100 -177.140 -2.760 -176.810 ;
        RECT 6.360 -177.140 6.700 -176.810 ;
        RECT 6.820 -177.140 7.160 -176.810 ;
        RECT 16.280 -177.140 16.620 -176.810 ;
        RECT 16.740 -177.140 17.080 -176.810 ;
        RECT -283.590 -177.900 -283.250 -177.570 ;
        RECT -273.670 -177.900 -273.330 -177.570 ;
        RECT -263.750 -177.900 -263.410 -177.570 ;
        RECT -253.830 -177.900 -253.490 -177.570 ;
        RECT -243.910 -177.900 -243.570 -177.570 ;
        RECT -233.990 -177.900 -233.650 -177.570 ;
        RECT -224.070 -177.900 -223.730 -177.570 ;
        RECT -214.150 -177.900 -213.810 -177.570 ;
        RECT -204.230 -177.900 -203.890 -177.570 ;
        RECT -194.310 -177.900 -193.970 -177.570 ;
        RECT -184.390 -177.900 -184.050 -177.570 ;
        RECT -174.470 -177.900 -174.130 -177.570 ;
        RECT -164.550 -177.900 -164.210 -177.570 ;
        RECT -154.630 -177.900 -154.290 -177.570 ;
        RECT -144.710 -177.900 -144.370 -177.570 ;
        RECT -134.790 -177.900 -134.450 -177.570 ;
        RECT -124.870 -177.900 -124.530 -177.570 ;
        RECT -114.950 -177.900 -114.610 -177.570 ;
        RECT -105.030 -177.900 -104.690 -177.570 ;
        RECT -95.110 -177.900 -94.770 -177.570 ;
        RECT -85.190 -177.900 -84.850 -177.570 ;
        RECT -75.270 -177.900 -74.930 -177.570 ;
        RECT -65.350 -177.900 -65.010 -177.570 ;
        RECT -55.430 -177.900 -55.090 -177.570 ;
        RECT -45.510 -177.900 -45.170 -177.570 ;
        RECT -35.590 -177.900 -35.250 -177.570 ;
        RECT -25.670 -177.900 -25.330 -177.570 ;
        RECT -15.750 -177.900 -15.410 -177.570 ;
        RECT -5.830 -177.900 -5.490 -177.570 ;
        RECT 4.090 -177.900 4.430 -177.570 ;
        RECT 14.010 -177.900 14.350 -177.570 ;
      LAYER met4 ;
        RECT -336.410 94.600 -323.960 94.660 ;
        RECT -336.500 94.560 -299.580 94.600 ;
        RECT 68.120 94.560 119.650 94.590 ;
        RECT -336.500 89.420 119.650 94.560 ;
        RECT -336.500 89.390 72.030 89.420 ;
        RECT -336.500 89.380 -299.580 89.390 ;
        RECT -336.410 10.550 -323.960 89.380 ;
        RECT -338.520 10.510 -301.600 10.550 ;
        RECT 66.100 10.510 117.630 10.540 ;
        RECT -338.520 5.370 117.630 10.510 ;
        RECT -338.520 5.340 70.010 5.370 ;
        RECT -338.520 5.330 -301.600 5.340 ;
        RECT -336.410 -78.400 -323.960 5.330 ;
        RECT -338.160 -78.440 -301.240 -78.400 ;
        RECT 66.460 -78.440 117.990 -78.410 ;
        RECT -338.160 -83.580 117.990 -78.440 ;
        RECT -338.160 -83.610 70.370 -83.580 ;
        RECT -338.160 -83.620 -301.240 -83.610 ;
        RECT -336.410 -172.980 -323.960 -83.620 ;
        RECT -339.920 -173.020 -303.000 -172.980 ;
        RECT 64.700 -173.020 116.230 -172.990 ;
        RECT -339.920 -178.160 116.230 -173.020 ;
        RECT -339.920 -178.190 68.610 -178.160 ;
        RECT -339.920 -178.200 -303.000 -178.190 ;
        RECT -336.410 -178.710 -323.960 -178.200 ;
    END
  END vssd1
  PIN o_ranQ[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 16.295 5.015 16.800 5.095 ;
        RECT 17.600 5.015 18.505 5.105 ;
        RECT 16.295 4.835 18.505 5.015 ;
      LAYER mcon ;
        RECT 16.485 4.925 16.655 5.095 ;
        RECT 17.850 4.925 18.020 5.095 ;
      LAYER met1 ;
        RECT 16.420 4.830 18.110 5.130 ;
        RECT 16.600 4.130 17.600 4.830 ;
    END
  END o_ranQ[65]
  PIN o_ranQ[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 11.335 10.825 13.545 11.005 ;
        RECT 11.335 10.745 11.840 10.825 ;
        RECT 12.640 10.735 13.545 10.825 ;
      LAYER mcon ;
        RECT 11.525 10.745 11.695 10.915 ;
        RECT 12.890 10.745 13.060 10.915 ;
      LAYER met1 ;
        RECT 11.640 11.010 12.640 11.710 ;
        RECT 11.460 10.710 13.150 11.010 ;
    END
  END o_ranQ[66]
  PIN o_ranQ[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 6.375 5.015 6.880 5.095 ;
        RECT 7.680 5.015 8.585 5.105 ;
        RECT 6.375 4.835 8.585 5.015 ;
      LAYER mcon ;
        RECT 6.565 4.925 6.735 5.095 ;
        RECT 7.930 4.925 8.100 5.095 ;
      LAYER met1 ;
        RECT 6.500 4.830 8.190 5.130 ;
        RECT 6.680 4.130 7.680 4.830 ;
    END
  END o_ranQ[67]
  PIN o_ranQ[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 21.255 10.825 23.465 11.005 ;
        RECT 21.255 10.745 21.760 10.825 ;
        RECT 22.560 10.735 23.465 10.825 ;
      LAYER mcon ;
        RECT 21.445 10.745 21.615 10.915 ;
        RECT 22.810 10.745 22.980 10.915 ;
      LAYER met1 ;
        RECT 21.560 11.010 22.560 11.710 ;
        RECT 21.380 10.710 23.070 11.010 ;
    END
  END o_ranQ[64]
  PIN o_ranQ[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 1.415 10.825 3.625 11.005 ;
        RECT 1.415 10.745 1.920 10.825 ;
        RECT 2.720 10.735 3.625 10.825 ;
      LAYER mcon ;
        RECT 1.605 10.745 1.775 10.915 ;
        RECT 2.970 10.745 3.140 10.915 ;
      LAYER met1 ;
        RECT 1.720 11.010 2.720 11.710 ;
        RECT 1.540 10.710 3.230 11.010 ;
    END
  END o_ranQ[68]
  PIN o_ranQ[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -3.545 5.015 -3.040 5.095 ;
        RECT -2.240 5.015 -1.335 5.105 ;
        RECT -3.545 4.835 -1.335 5.015 ;
      LAYER mcon ;
        RECT -3.355 4.925 -3.185 5.095 ;
        RECT -1.990 4.925 -1.820 5.095 ;
      LAYER met1 ;
        RECT -3.420 4.830 -1.730 5.130 ;
        RECT -3.240 4.130 -2.240 4.830 ;
    END
  END o_ranQ[69]
  PIN o_ranQ[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -8.505 10.825 -6.295 11.005 ;
        RECT -8.505 10.745 -8.000 10.825 ;
        RECT -7.200 10.735 -6.295 10.825 ;
      LAYER mcon ;
        RECT -8.315 10.745 -8.145 10.915 ;
        RECT -6.950 10.745 -6.780 10.915 ;
      LAYER met1 ;
        RECT -8.200 11.010 -7.200 11.710 ;
        RECT -8.380 10.710 -6.690 11.010 ;
    END
  END o_ranQ[70]
  PIN o_ranQ[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -13.465 5.015 -12.960 5.095 ;
        RECT -12.160 5.015 -11.255 5.105 ;
        RECT -13.465 4.835 -11.255 5.015 ;
      LAYER mcon ;
        RECT -13.275 4.925 -13.105 5.095 ;
        RECT -11.910 4.925 -11.740 5.095 ;
      LAYER met1 ;
        RECT -13.340 4.830 -11.650 5.130 ;
        RECT -13.160 4.130 -12.160 4.830 ;
    END
  END o_ranQ[71]
  PIN o_ranQ[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -18.425 10.825 -16.215 11.005 ;
        RECT -18.425 10.745 -17.920 10.825 ;
        RECT -17.120 10.735 -16.215 10.825 ;
      LAYER mcon ;
        RECT -18.235 10.745 -18.065 10.915 ;
        RECT -16.870 10.745 -16.700 10.915 ;
      LAYER met1 ;
        RECT -18.120 11.010 -17.120 11.710 ;
        RECT -18.300 10.710 -16.610 11.010 ;
    END
  END o_ranQ[72]
  PIN o_ranQ[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -23.385 5.015 -22.880 5.095 ;
        RECT -22.080 5.015 -21.175 5.105 ;
        RECT -23.385 4.835 -21.175 5.015 ;
      LAYER mcon ;
        RECT -23.195 4.925 -23.025 5.095 ;
        RECT -21.830 4.925 -21.660 5.095 ;
      LAYER met1 ;
        RECT -23.260 4.830 -21.570 5.130 ;
        RECT -23.080 4.130 -22.080 4.830 ;
    END
  END o_ranQ[73]
  PIN o_ranQ[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -28.345 10.825 -26.135 11.005 ;
        RECT -28.345 10.745 -27.840 10.825 ;
        RECT -27.040 10.735 -26.135 10.825 ;
      LAYER mcon ;
        RECT -28.155 10.745 -27.985 10.915 ;
        RECT -26.790 10.745 -26.620 10.915 ;
      LAYER met1 ;
        RECT -28.040 11.010 -27.040 11.710 ;
        RECT -28.220 10.710 -26.530 11.010 ;
    END
  END o_ranQ[74]
  PIN o_ranQ[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -33.305 5.015 -32.800 5.095 ;
        RECT -32.000 5.015 -31.095 5.105 ;
        RECT -33.305 4.835 -31.095 5.015 ;
      LAYER mcon ;
        RECT -33.115 4.925 -32.945 5.095 ;
        RECT -31.750 4.925 -31.580 5.095 ;
      LAYER met1 ;
        RECT -33.180 4.830 -31.490 5.130 ;
        RECT -33.000 4.130 -32.000 4.830 ;
    END
  END o_ranQ[75]
  PIN o_ranQ[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -38.265 10.825 -36.055 11.005 ;
        RECT -38.265 10.745 -37.760 10.825 ;
        RECT -36.960 10.735 -36.055 10.825 ;
      LAYER mcon ;
        RECT -38.075 10.745 -37.905 10.915 ;
        RECT -36.710 10.745 -36.540 10.915 ;
      LAYER met1 ;
        RECT -37.960 11.010 -36.960 11.710 ;
        RECT -38.140 10.710 -36.450 11.010 ;
    END
  END o_ranQ[76]
  PIN o_ranQ[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -43.225 5.015 -42.720 5.095 ;
        RECT -41.920 5.015 -41.015 5.105 ;
        RECT -43.225 4.835 -41.015 5.015 ;
      LAYER mcon ;
        RECT -43.035 4.925 -42.865 5.095 ;
        RECT -41.670 4.925 -41.500 5.095 ;
      LAYER met1 ;
        RECT -43.100 4.830 -41.410 5.130 ;
        RECT -42.920 4.130 -41.920 4.830 ;
    END
  END o_ranQ[77]
  PIN o_ranQ[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -48.185 10.825 -45.975 11.005 ;
        RECT -48.185 10.745 -47.680 10.825 ;
        RECT -46.880 10.735 -45.975 10.825 ;
      LAYER mcon ;
        RECT -47.995 10.745 -47.825 10.915 ;
        RECT -46.630 10.745 -46.460 10.915 ;
      LAYER met1 ;
        RECT -47.880 11.010 -46.880 11.710 ;
        RECT -48.060 10.710 -46.370 11.010 ;
    END
  END o_ranQ[78]
  PIN o_ranQ[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -53.145 5.015 -52.640 5.095 ;
        RECT -51.840 5.015 -50.935 5.105 ;
        RECT -53.145 4.835 -50.935 5.015 ;
      LAYER mcon ;
        RECT -52.955 4.925 -52.785 5.095 ;
        RECT -51.590 4.925 -51.420 5.095 ;
      LAYER met1 ;
        RECT -53.020 4.830 -51.330 5.130 ;
        RECT -52.840 4.130 -51.840 4.830 ;
    END
  END o_ranQ[79]
  PIN o_ranQ[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -63.065 5.015 -62.560 5.095 ;
        RECT -61.760 5.015 -60.855 5.105 ;
        RECT -63.065 4.835 -60.855 5.015 ;
      LAYER mcon ;
        RECT -62.875 4.925 -62.705 5.095 ;
        RECT -61.510 4.925 -61.340 5.095 ;
      LAYER met1 ;
        RECT -62.940 4.830 -61.250 5.130 ;
        RECT -62.760 4.130 -61.760 4.830 ;
    END
  END o_ranQ[81]
  PIN o_ranQ[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -68.025 10.825 -65.815 11.005 ;
        RECT -68.025 10.745 -67.520 10.825 ;
        RECT -66.720 10.735 -65.815 10.825 ;
      LAYER mcon ;
        RECT -67.835 10.745 -67.665 10.915 ;
        RECT -66.470 10.745 -66.300 10.915 ;
      LAYER met1 ;
        RECT -67.720 11.010 -66.720 11.710 ;
        RECT -67.900 10.710 -66.210 11.010 ;
    END
  END o_ranQ[82]
  PIN o_ranQ[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -72.985 5.015 -72.480 5.095 ;
        RECT -71.680 5.015 -70.775 5.105 ;
        RECT -72.985 4.835 -70.775 5.015 ;
      LAYER mcon ;
        RECT -72.795 4.925 -72.625 5.095 ;
        RECT -71.430 4.925 -71.260 5.095 ;
      LAYER met1 ;
        RECT -72.860 4.830 -71.170 5.130 ;
        RECT -72.680 4.130 -71.680 4.830 ;
    END
  END o_ranQ[83]
  PIN o_ranQ[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -58.105 10.825 -55.895 11.005 ;
        RECT -58.105 10.745 -57.600 10.825 ;
        RECT -56.800 10.735 -55.895 10.825 ;
      LAYER mcon ;
        RECT -57.915 10.745 -57.745 10.915 ;
        RECT -56.550 10.745 -56.380 10.915 ;
      LAYER met1 ;
        RECT -57.800 11.010 -56.800 11.710 ;
        RECT -57.980 10.710 -56.290 11.010 ;
    END
  END o_ranQ[80]
  PIN o_ranQ[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -77.945 10.825 -75.735 11.005 ;
        RECT -77.945 10.745 -77.440 10.825 ;
        RECT -76.640 10.735 -75.735 10.825 ;
      LAYER mcon ;
        RECT -77.755 10.745 -77.585 10.915 ;
        RECT -76.390 10.745 -76.220 10.915 ;
      LAYER met1 ;
        RECT -77.640 11.010 -76.640 11.710 ;
        RECT -77.820 10.710 -76.130 11.010 ;
    END
  END o_ranQ[84]
  PIN o_ranQ[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -82.905 5.015 -82.400 5.095 ;
        RECT -81.600 5.015 -80.695 5.105 ;
        RECT -82.905 4.835 -80.695 5.015 ;
      LAYER mcon ;
        RECT -82.715 4.925 -82.545 5.095 ;
        RECT -81.350 4.925 -81.180 5.095 ;
      LAYER met1 ;
        RECT -82.780 4.830 -81.090 5.130 ;
        RECT -82.600 4.130 -81.600 4.830 ;
    END
  END o_ranQ[85]
  PIN o_ranQ[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -87.865 10.825 -85.655 11.005 ;
        RECT -87.865 10.745 -87.360 10.825 ;
        RECT -86.560 10.735 -85.655 10.825 ;
      LAYER mcon ;
        RECT -87.675 10.745 -87.505 10.915 ;
        RECT -86.310 10.745 -86.140 10.915 ;
      LAYER met1 ;
        RECT -87.560 11.010 -86.560 11.710 ;
        RECT -87.740 10.710 -86.050 11.010 ;
    END
  END o_ranQ[86]
  PIN o_ranQ[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -92.825 5.015 -92.320 5.095 ;
        RECT -91.520 5.015 -90.615 5.105 ;
        RECT -92.825 4.835 -90.615 5.015 ;
      LAYER mcon ;
        RECT -92.635 4.925 -92.465 5.095 ;
        RECT -91.270 4.925 -91.100 5.095 ;
      LAYER met1 ;
        RECT -92.700 4.830 -91.010 5.130 ;
        RECT -92.520 4.130 -91.520 4.830 ;
    END
  END o_ranQ[87]
  PIN o_ranQ[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -97.785 10.825 -95.575 11.005 ;
        RECT -97.785 10.745 -97.280 10.825 ;
        RECT -96.480 10.735 -95.575 10.825 ;
      LAYER mcon ;
        RECT -97.595 10.745 -97.425 10.915 ;
        RECT -96.230 10.745 -96.060 10.915 ;
      LAYER met1 ;
        RECT -97.480 11.010 -96.480 11.710 ;
        RECT -97.660 10.710 -95.970 11.010 ;
    END
  END o_ranQ[88]
  PIN o_ranQ[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -102.745 5.015 -102.240 5.095 ;
        RECT -101.440 5.015 -100.535 5.105 ;
        RECT -102.745 4.835 -100.535 5.015 ;
      LAYER mcon ;
        RECT -102.555 4.925 -102.385 5.095 ;
        RECT -101.190 4.925 -101.020 5.095 ;
      LAYER met1 ;
        RECT -102.620 4.830 -100.930 5.130 ;
        RECT -102.440 4.130 -101.440 4.830 ;
    END
  END o_ranQ[89]
  PIN o_ranQ[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -107.705 10.825 -105.495 11.005 ;
        RECT -107.705 10.745 -107.200 10.825 ;
        RECT -106.400 10.735 -105.495 10.825 ;
      LAYER mcon ;
        RECT -107.515 10.745 -107.345 10.915 ;
        RECT -106.150 10.745 -105.980 10.915 ;
      LAYER met1 ;
        RECT -107.400 11.010 -106.400 11.710 ;
        RECT -107.580 10.710 -105.890 11.010 ;
    END
  END o_ranQ[90]
  PIN o_ranQ[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -112.665 5.015 -112.160 5.095 ;
        RECT -111.360 5.015 -110.455 5.105 ;
        RECT -112.665 4.835 -110.455 5.015 ;
      LAYER mcon ;
        RECT -112.475 4.925 -112.305 5.095 ;
        RECT -111.110 4.925 -110.940 5.095 ;
      LAYER met1 ;
        RECT -112.540 4.830 -110.850 5.130 ;
        RECT -112.360 4.130 -111.360 4.830 ;
    END
  END o_ranQ[91]
  PIN o_ranQ[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -117.625 10.825 -115.415 11.005 ;
        RECT -117.625 10.745 -117.120 10.825 ;
        RECT -116.320 10.735 -115.415 10.825 ;
      LAYER mcon ;
        RECT -117.435 10.745 -117.265 10.915 ;
        RECT -116.070 10.745 -115.900 10.915 ;
      LAYER met1 ;
        RECT -117.320 11.010 -116.320 11.710 ;
        RECT -117.500 10.710 -115.810 11.010 ;
    END
  END o_ranQ[92]
  PIN o_ranQ[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -122.585 5.015 -122.080 5.095 ;
        RECT -121.280 5.015 -120.375 5.105 ;
        RECT -122.585 4.835 -120.375 5.015 ;
      LAYER mcon ;
        RECT -122.395 4.925 -122.225 5.095 ;
        RECT -121.030 4.925 -120.860 5.095 ;
      LAYER met1 ;
        RECT -122.460 4.830 -120.770 5.130 ;
        RECT -122.280 4.130 -121.280 4.830 ;
    END
  END o_ranQ[93]
  PIN o_ranQ[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -127.545 10.825 -125.335 11.005 ;
        RECT -127.545 10.745 -127.040 10.825 ;
        RECT -126.240 10.735 -125.335 10.825 ;
      LAYER mcon ;
        RECT -127.355 10.745 -127.185 10.915 ;
        RECT -125.990 10.745 -125.820 10.915 ;
      LAYER met1 ;
        RECT -127.240 11.010 -126.240 11.710 ;
        RECT -127.420 10.710 -125.730 11.010 ;
    END
  END o_ranQ[94]
  PIN o_ranQ[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -132.505 5.015 -132.000 5.095 ;
        RECT -131.200 5.015 -130.295 5.105 ;
        RECT -132.505 4.835 -130.295 5.015 ;
      LAYER mcon ;
        RECT -132.315 4.925 -132.145 5.095 ;
        RECT -130.950 4.925 -130.780 5.095 ;
      LAYER met1 ;
        RECT -132.380 4.830 -130.690 5.130 ;
        RECT -132.200 4.130 -131.200 4.830 ;
    END
  END o_ranQ[95]
  PIN o_ranQ[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -142.425 5.015 -141.920 5.095 ;
        RECT -141.120 5.015 -140.215 5.105 ;
        RECT -142.425 4.835 -140.215 5.015 ;
      LAYER mcon ;
        RECT -142.235 4.925 -142.065 5.095 ;
        RECT -140.870 4.925 -140.700 5.095 ;
      LAYER met1 ;
        RECT -142.300 4.830 -140.610 5.130 ;
        RECT -142.120 4.130 -141.120 4.830 ;
    END
  END o_ranQ[97]
  PIN o_ranQ[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -147.385 10.825 -145.175 11.005 ;
        RECT -147.385 10.745 -146.880 10.825 ;
        RECT -146.080 10.735 -145.175 10.825 ;
      LAYER mcon ;
        RECT -147.195 10.745 -147.025 10.915 ;
        RECT -145.830 10.745 -145.660 10.915 ;
      LAYER met1 ;
        RECT -147.080 11.010 -146.080 11.710 ;
        RECT -147.260 10.710 -145.570 11.010 ;
    END
  END o_ranQ[98]
  PIN o_ranQ[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -152.345 5.015 -151.840 5.095 ;
        RECT -151.040 5.015 -150.135 5.105 ;
        RECT -152.345 4.835 -150.135 5.015 ;
      LAYER mcon ;
        RECT -152.155 4.925 -151.985 5.095 ;
        RECT -150.790 4.925 -150.620 5.095 ;
      LAYER met1 ;
        RECT -152.220 4.830 -150.530 5.130 ;
        RECT -152.040 4.130 -151.040 4.830 ;
    END
  END o_ranQ[99]
  PIN o_ranQ[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -137.465 10.825 -135.255 11.005 ;
        RECT -137.465 10.745 -136.960 10.825 ;
        RECT -136.160 10.735 -135.255 10.825 ;
      LAYER mcon ;
        RECT -137.275 10.745 -137.105 10.915 ;
        RECT -135.910 10.745 -135.740 10.915 ;
      LAYER met1 ;
        RECT -137.160 11.010 -136.160 11.710 ;
        RECT -137.340 10.710 -135.650 11.010 ;
    END
  END o_ranQ[96]
  PIN o_ranQ[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -157.305 10.825 -155.095 11.005 ;
        RECT -157.305 10.745 -156.800 10.825 ;
        RECT -156.000 10.735 -155.095 10.825 ;
      LAYER mcon ;
        RECT -157.115 10.745 -156.945 10.915 ;
        RECT -155.750 10.745 -155.580 10.915 ;
      LAYER met1 ;
        RECT -157.000 11.010 -156.000 11.710 ;
        RECT -157.180 10.710 -155.490 11.010 ;
    END
  END o_ranQ[100]
  PIN o_ranQ[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -162.265 5.015 -161.760 5.095 ;
        RECT -160.960 5.015 -160.055 5.105 ;
        RECT -162.265 4.835 -160.055 5.015 ;
      LAYER mcon ;
        RECT -162.075 4.925 -161.905 5.095 ;
        RECT -160.710 4.925 -160.540 5.095 ;
      LAYER met1 ;
        RECT -162.140 4.830 -160.450 5.130 ;
        RECT -161.960 4.130 -160.960 4.830 ;
    END
  END o_ranQ[101]
  PIN o_ranQ[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -167.225 10.825 -165.015 11.005 ;
        RECT -167.225 10.745 -166.720 10.825 ;
        RECT -165.920 10.735 -165.015 10.825 ;
      LAYER mcon ;
        RECT -167.035 10.745 -166.865 10.915 ;
        RECT -165.670 10.745 -165.500 10.915 ;
      LAYER met1 ;
        RECT -166.920 11.010 -165.920 11.710 ;
        RECT -167.100 10.710 -165.410 11.010 ;
    END
  END o_ranQ[102]
  PIN o_ranQ[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -172.185 5.015 -171.680 5.095 ;
        RECT -170.880 5.015 -169.975 5.105 ;
        RECT -172.185 4.835 -169.975 5.015 ;
      LAYER mcon ;
        RECT -171.995 4.925 -171.825 5.095 ;
        RECT -170.630 4.925 -170.460 5.095 ;
      LAYER met1 ;
        RECT -172.060 4.830 -170.370 5.130 ;
        RECT -171.880 4.130 -170.880 4.830 ;
    END
  END o_ranQ[103]
  PIN o_ranQ[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -177.145 10.825 -174.935 11.005 ;
        RECT -177.145 10.745 -176.640 10.825 ;
        RECT -175.840 10.735 -174.935 10.825 ;
      LAYER mcon ;
        RECT -176.955 10.745 -176.785 10.915 ;
        RECT -175.590 10.745 -175.420 10.915 ;
      LAYER met1 ;
        RECT -176.840 11.010 -175.840 11.710 ;
        RECT -177.020 10.710 -175.330 11.010 ;
    END
  END o_ranQ[104]
  PIN o_ranQ[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -182.105 5.015 -181.600 5.095 ;
        RECT -180.800 5.015 -179.895 5.105 ;
        RECT -182.105 4.835 -179.895 5.015 ;
      LAYER mcon ;
        RECT -181.915 4.925 -181.745 5.095 ;
        RECT -180.550 4.925 -180.380 5.095 ;
      LAYER met1 ;
        RECT -181.980 4.830 -180.290 5.130 ;
        RECT -181.800 4.130 -180.800 4.830 ;
    END
  END o_ranQ[105]
  PIN o_ranQ[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -187.065 10.825 -184.855 11.005 ;
        RECT -187.065 10.745 -186.560 10.825 ;
        RECT -185.760 10.735 -184.855 10.825 ;
      LAYER mcon ;
        RECT -186.875 10.745 -186.705 10.915 ;
        RECT -185.510 10.745 -185.340 10.915 ;
      LAYER met1 ;
        RECT -186.760 11.010 -185.760 11.710 ;
        RECT -186.940 10.710 -185.250 11.010 ;
    END
  END o_ranQ[106]
  PIN o_ranQ[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -192.025 5.015 -191.520 5.095 ;
        RECT -190.720 5.015 -189.815 5.105 ;
        RECT -192.025 4.835 -189.815 5.015 ;
      LAYER mcon ;
        RECT -191.835 4.925 -191.665 5.095 ;
        RECT -190.470 4.925 -190.300 5.095 ;
      LAYER met1 ;
        RECT -191.900 4.830 -190.210 5.130 ;
        RECT -191.720 4.130 -190.720 4.830 ;
    END
  END o_ranQ[107]
  PIN o_ranQ[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -196.985 10.825 -194.775 11.005 ;
        RECT -196.985 10.745 -196.480 10.825 ;
        RECT -195.680 10.735 -194.775 10.825 ;
      LAYER mcon ;
        RECT -196.795 10.745 -196.625 10.915 ;
        RECT -195.430 10.745 -195.260 10.915 ;
      LAYER met1 ;
        RECT -196.680 11.010 -195.680 11.710 ;
        RECT -196.860 10.710 -195.170 11.010 ;
    END
  END o_ranQ[108]
  PIN o_ranQ[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -201.945 5.015 -201.440 5.095 ;
        RECT -200.640 5.015 -199.735 5.105 ;
        RECT -201.945 4.835 -199.735 5.015 ;
      LAYER mcon ;
        RECT -201.755 4.925 -201.585 5.095 ;
        RECT -200.390 4.925 -200.220 5.095 ;
      LAYER met1 ;
        RECT -201.820 4.830 -200.130 5.130 ;
        RECT -201.640 4.130 -200.640 4.830 ;
    END
  END o_ranQ[109]
  PIN o_ranQ[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -206.905 10.825 -204.695 11.005 ;
        RECT -206.905 10.745 -206.400 10.825 ;
        RECT -205.600 10.735 -204.695 10.825 ;
      LAYER mcon ;
        RECT -206.715 10.745 -206.545 10.915 ;
        RECT -205.350 10.745 -205.180 10.915 ;
      LAYER met1 ;
        RECT -206.600 11.010 -205.600 11.710 ;
        RECT -206.780 10.710 -205.090 11.010 ;
    END
  END o_ranQ[110]
  PIN o_ranQ[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -211.865 5.015 -211.360 5.095 ;
        RECT -210.560 5.015 -209.655 5.105 ;
        RECT -211.865 4.835 -209.655 5.015 ;
      LAYER mcon ;
        RECT -211.675 4.925 -211.505 5.095 ;
        RECT -210.310 4.925 -210.140 5.095 ;
      LAYER met1 ;
        RECT -211.740 4.830 -210.050 5.130 ;
        RECT -211.560 4.130 -210.560 4.830 ;
    END
  END o_ranQ[111]
  PIN o_ranQ[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -221.785 5.015 -221.280 5.095 ;
        RECT -220.480 5.015 -219.575 5.105 ;
        RECT -221.785 4.835 -219.575 5.015 ;
      LAYER mcon ;
        RECT -221.595 4.925 -221.425 5.095 ;
        RECT -220.230 4.925 -220.060 5.095 ;
      LAYER met1 ;
        RECT -221.660 4.830 -219.970 5.130 ;
        RECT -221.480 4.130 -220.480 4.830 ;
    END
  END o_ranQ[113]
  PIN o_ranQ[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -226.745 10.825 -224.535 11.005 ;
        RECT -226.745 10.745 -226.240 10.825 ;
        RECT -225.440 10.735 -224.535 10.825 ;
      LAYER mcon ;
        RECT -226.555 10.745 -226.385 10.915 ;
        RECT -225.190 10.745 -225.020 10.915 ;
      LAYER met1 ;
        RECT -226.440 11.010 -225.440 11.710 ;
        RECT -226.620 10.710 -224.930 11.010 ;
    END
  END o_ranQ[114]
  PIN o_ranQ[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -231.705 5.015 -231.200 5.095 ;
        RECT -230.400 5.015 -229.495 5.105 ;
        RECT -231.705 4.835 -229.495 5.015 ;
      LAYER mcon ;
        RECT -231.515 4.925 -231.345 5.095 ;
        RECT -230.150 4.925 -229.980 5.095 ;
      LAYER met1 ;
        RECT -231.580 4.830 -229.890 5.130 ;
        RECT -231.400 4.130 -230.400 4.830 ;
    END
  END o_ranQ[115]
  PIN o_ranQ[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -216.825 10.825 -214.615 11.005 ;
        RECT -216.825 10.745 -216.320 10.825 ;
        RECT -215.520 10.735 -214.615 10.825 ;
      LAYER mcon ;
        RECT -216.635 10.745 -216.465 10.915 ;
        RECT -215.270 10.745 -215.100 10.915 ;
      LAYER met1 ;
        RECT -216.520 11.010 -215.520 11.710 ;
        RECT -216.700 10.710 -215.010 11.010 ;
    END
  END o_ranQ[112]
  PIN o_ranQ[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -236.665 10.825 -234.455 11.005 ;
        RECT -236.665 10.745 -236.160 10.825 ;
        RECT -235.360 10.735 -234.455 10.825 ;
      LAYER mcon ;
        RECT -236.475 10.745 -236.305 10.915 ;
        RECT -235.110 10.745 -234.940 10.915 ;
      LAYER met1 ;
        RECT -236.360 11.010 -235.360 11.710 ;
        RECT -236.540 10.710 -234.850 11.010 ;
    END
  END o_ranQ[116]
  PIN o_ranQ[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -241.625 5.015 -241.120 5.095 ;
        RECT -240.320 5.015 -239.415 5.105 ;
        RECT -241.625 4.835 -239.415 5.015 ;
      LAYER mcon ;
        RECT -241.435 4.925 -241.265 5.095 ;
        RECT -240.070 4.925 -239.900 5.095 ;
      LAYER met1 ;
        RECT -241.500 4.830 -239.810 5.130 ;
        RECT -241.320 4.130 -240.320 4.830 ;
    END
  END o_ranQ[117]
  PIN o_ranQ[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -246.585 10.825 -244.375 11.005 ;
        RECT -246.585 10.745 -246.080 10.825 ;
        RECT -245.280 10.735 -244.375 10.825 ;
      LAYER mcon ;
        RECT -246.395 10.745 -246.225 10.915 ;
        RECT -245.030 10.745 -244.860 10.915 ;
      LAYER met1 ;
        RECT -246.280 11.010 -245.280 11.710 ;
        RECT -246.460 10.710 -244.770 11.010 ;
    END
  END o_ranQ[118]
  PIN o_ranQ[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -251.545 5.015 -251.040 5.095 ;
        RECT -250.240 5.015 -249.335 5.105 ;
        RECT -251.545 4.835 -249.335 5.015 ;
      LAYER mcon ;
        RECT -251.355 4.925 -251.185 5.095 ;
        RECT -249.990 4.925 -249.820 5.095 ;
      LAYER met1 ;
        RECT -251.420 4.830 -249.730 5.130 ;
        RECT -251.240 4.130 -250.240 4.830 ;
    END
  END o_ranQ[119]
  PIN o_ranQ[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -256.505 10.825 -254.295 11.005 ;
        RECT -256.505 10.745 -256.000 10.825 ;
        RECT -255.200 10.735 -254.295 10.825 ;
      LAYER mcon ;
        RECT -256.315 10.745 -256.145 10.915 ;
        RECT -254.950 10.745 -254.780 10.915 ;
      LAYER met1 ;
        RECT -256.200 11.010 -255.200 11.710 ;
        RECT -256.380 10.710 -254.690 11.010 ;
    END
  END o_ranQ[120]
  PIN o_ranQ[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -261.465 5.015 -260.960 5.095 ;
        RECT -260.160 5.015 -259.255 5.105 ;
        RECT -261.465 4.835 -259.255 5.015 ;
      LAYER mcon ;
        RECT -261.275 4.925 -261.105 5.095 ;
        RECT -259.910 4.925 -259.740 5.095 ;
      LAYER met1 ;
        RECT -261.340 4.830 -259.650 5.130 ;
        RECT -261.160 4.130 -260.160 4.830 ;
    END
  END o_ranQ[121]
  PIN o_ranQ[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -266.425 10.825 -264.215 11.005 ;
        RECT -266.425 10.745 -265.920 10.825 ;
        RECT -265.120 10.735 -264.215 10.825 ;
      LAYER mcon ;
        RECT -266.235 10.745 -266.065 10.915 ;
        RECT -264.870 10.745 -264.700 10.915 ;
      LAYER met1 ;
        RECT -266.120 11.010 -265.120 11.710 ;
        RECT -266.300 10.710 -264.610 11.010 ;
    END
  END o_ranQ[122]
  PIN o_ranQ[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -271.385 5.015 -270.880 5.095 ;
        RECT -270.080 5.015 -269.175 5.105 ;
        RECT -271.385 4.835 -269.175 5.015 ;
      LAYER mcon ;
        RECT -271.195 4.925 -271.025 5.095 ;
        RECT -269.830 4.925 -269.660 5.095 ;
      LAYER met1 ;
        RECT -271.260 4.830 -269.570 5.130 ;
        RECT -271.080 4.130 -270.080 4.830 ;
    END
  END o_ranQ[123]
  PIN o_ranQ[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -276.345 10.825 -274.135 11.005 ;
        RECT -276.345 10.745 -275.840 10.825 ;
        RECT -275.040 10.735 -274.135 10.825 ;
      LAYER mcon ;
        RECT -276.155 10.745 -275.985 10.915 ;
        RECT -274.790 10.745 -274.620 10.915 ;
      LAYER met1 ;
        RECT -276.040 11.010 -275.040 11.710 ;
        RECT -276.220 10.710 -274.530 11.010 ;
    END
  END o_ranQ[124]
  PIN o_ranQ[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -281.305 5.015 -280.800 5.095 ;
        RECT -280.000 5.015 -279.095 5.105 ;
        RECT -281.305 4.835 -279.095 5.015 ;
      LAYER mcon ;
        RECT -281.115 4.925 -280.945 5.095 ;
        RECT -279.750 4.925 -279.580 5.095 ;
      LAYER met1 ;
        RECT -281.180 4.830 -279.490 5.130 ;
        RECT -281.000 4.130 -280.000 4.830 ;
    END
  END o_ranQ[125]
  PIN o_ranQ[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -286.265 10.825 -284.055 11.005 ;
        RECT -286.265 10.745 -285.760 10.825 ;
        RECT -284.960 10.735 -284.055 10.825 ;
      LAYER mcon ;
        RECT -286.075 10.745 -285.905 10.915 ;
        RECT -284.710 10.745 -284.540 10.915 ;
      LAYER met1 ;
        RECT -285.960 11.010 -284.960 11.710 ;
        RECT -286.140 10.710 -284.450 11.010 ;
    END
  END o_ranQ[126]
  PIN o_ranQ[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -291.225 5.015 -290.720 5.095 ;
        RECT -289.920 5.015 -289.015 5.105 ;
        RECT -291.225 4.835 -289.015 5.015 ;
      LAYER mcon ;
        RECT -291.035 4.925 -290.865 5.095 ;
        RECT -289.670 4.925 -289.500 5.095 ;
      LAYER met1 ;
        RECT -291.100 4.830 -289.410 5.130 ;
        RECT -290.920 4.130 -289.920 4.830 ;
    END
  END o_ranQ[127]
  PIN o_ranQ[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 16.655 -83.935 17.160 -83.855 ;
        RECT 17.960 -83.935 18.865 -83.845 ;
        RECT 16.655 -84.115 18.865 -83.935 ;
      LAYER mcon ;
        RECT 16.845 -84.025 17.015 -83.855 ;
        RECT 18.210 -84.025 18.380 -83.855 ;
      LAYER met1 ;
        RECT 16.780 -84.120 18.470 -83.820 ;
        RECT 16.960 -84.820 17.960 -84.120 ;
    END
  END o_ranQ[129]
  PIN o_ranQ[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 11.695 -78.125 13.905 -77.945 ;
        RECT 11.695 -78.205 12.200 -78.125 ;
        RECT 13.000 -78.215 13.905 -78.125 ;
      LAYER mcon ;
        RECT 11.885 -78.205 12.055 -78.035 ;
        RECT 13.250 -78.205 13.420 -78.035 ;
      LAYER met1 ;
        RECT 12.000 -77.940 13.000 -77.240 ;
        RECT 11.820 -78.240 13.510 -77.940 ;
    END
  END o_ranQ[130]
  PIN o_ranQ[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 6.735 -83.935 7.240 -83.855 ;
        RECT 8.040 -83.935 8.945 -83.845 ;
        RECT 6.735 -84.115 8.945 -83.935 ;
      LAYER mcon ;
        RECT 6.925 -84.025 7.095 -83.855 ;
        RECT 8.290 -84.025 8.460 -83.855 ;
      LAYER met1 ;
        RECT 6.860 -84.120 8.550 -83.820 ;
        RECT 7.040 -84.820 8.040 -84.120 ;
    END
  END o_ranQ[131]
  PIN o_ranQ[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 21.615 -78.125 23.825 -77.945 ;
        RECT 21.615 -78.205 22.120 -78.125 ;
        RECT 22.920 -78.215 23.825 -78.125 ;
      LAYER mcon ;
        RECT 21.805 -78.205 21.975 -78.035 ;
        RECT 23.170 -78.205 23.340 -78.035 ;
      LAYER met1 ;
        RECT 21.920 -77.940 22.920 -77.240 ;
        RECT 21.740 -78.240 23.430 -77.940 ;
    END
  END o_ranQ[128]
  PIN o_ranQ[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 1.775 -78.125 3.985 -77.945 ;
        RECT 1.775 -78.205 2.280 -78.125 ;
        RECT 3.080 -78.215 3.985 -78.125 ;
      LAYER mcon ;
        RECT 1.965 -78.205 2.135 -78.035 ;
        RECT 3.330 -78.205 3.500 -78.035 ;
      LAYER met1 ;
        RECT 2.080 -77.940 3.080 -77.240 ;
        RECT 1.900 -78.240 3.590 -77.940 ;
    END
  END o_ranQ[132]
  PIN o_ranQ[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -3.185 -83.935 -2.680 -83.855 ;
        RECT -1.880 -83.935 -0.975 -83.845 ;
        RECT -3.185 -84.115 -0.975 -83.935 ;
      LAYER mcon ;
        RECT -2.995 -84.025 -2.825 -83.855 ;
        RECT -1.630 -84.025 -1.460 -83.855 ;
      LAYER met1 ;
        RECT -3.060 -84.120 -1.370 -83.820 ;
        RECT -2.880 -84.820 -1.880 -84.120 ;
    END
  END o_ranQ[133]
  PIN o_ranQ[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -8.145 -78.125 -5.935 -77.945 ;
        RECT -8.145 -78.205 -7.640 -78.125 ;
        RECT -6.840 -78.215 -5.935 -78.125 ;
      LAYER mcon ;
        RECT -7.955 -78.205 -7.785 -78.035 ;
        RECT -6.590 -78.205 -6.420 -78.035 ;
      LAYER met1 ;
        RECT -7.840 -77.940 -6.840 -77.240 ;
        RECT -8.020 -78.240 -6.330 -77.940 ;
    END
  END o_ranQ[134]
  PIN o_ranQ[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -13.105 -83.935 -12.600 -83.855 ;
        RECT -11.800 -83.935 -10.895 -83.845 ;
        RECT -13.105 -84.115 -10.895 -83.935 ;
      LAYER mcon ;
        RECT -12.915 -84.025 -12.745 -83.855 ;
        RECT -11.550 -84.025 -11.380 -83.855 ;
      LAYER met1 ;
        RECT -12.980 -84.120 -11.290 -83.820 ;
        RECT -12.800 -84.820 -11.800 -84.120 ;
    END
  END o_ranQ[135]
  PIN o_ranQ[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -18.065 -78.125 -15.855 -77.945 ;
        RECT -18.065 -78.205 -17.560 -78.125 ;
        RECT -16.760 -78.215 -15.855 -78.125 ;
      LAYER mcon ;
        RECT -17.875 -78.205 -17.705 -78.035 ;
        RECT -16.510 -78.205 -16.340 -78.035 ;
      LAYER met1 ;
        RECT -17.760 -77.940 -16.760 -77.240 ;
        RECT -17.940 -78.240 -16.250 -77.940 ;
    END
  END o_ranQ[136]
  PIN o_ranQ[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -23.025 -83.935 -22.520 -83.855 ;
        RECT -21.720 -83.935 -20.815 -83.845 ;
        RECT -23.025 -84.115 -20.815 -83.935 ;
      LAYER mcon ;
        RECT -22.835 -84.025 -22.665 -83.855 ;
        RECT -21.470 -84.025 -21.300 -83.855 ;
      LAYER met1 ;
        RECT -22.900 -84.120 -21.210 -83.820 ;
        RECT -22.720 -84.820 -21.720 -84.120 ;
    END
  END o_ranQ[137]
  PIN o_ranQ[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -27.985 -78.125 -25.775 -77.945 ;
        RECT -27.985 -78.205 -27.480 -78.125 ;
        RECT -26.680 -78.215 -25.775 -78.125 ;
      LAYER mcon ;
        RECT -27.795 -78.205 -27.625 -78.035 ;
        RECT -26.430 -78.205 -26.260 -78.035 ;
      LAYER met1 ;
        RECT -27.680 -77.940 -26.680 -77.240 ;
        RECT -27.860 -78.240 -26.170 -77.940 ;
    END
  END o_ranQ[138]
  PIN o_ranQ[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -32.945 -83.935 -32.440 -83.855 ;
        RECT -31.640 -83.935 -30.735 -83.845 ;
        RECT -32.945 -84.115 -30.735 -83.935 ;
      LAYER mcon ;
        RECT -32.755 -84.025 -32.585 -83.855 ;
        RECT -31.390 -84.025 -31.220 -83.855 ;
      LAYER met1 ;
        RECT -32.820 -84.120 -31.130 -83.820 ;
        RECT -32.640 -84.820 -31.640 -84.120 ;
    END
  END o_ranQ[139]
  PIN o_ranQ[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -37.905 -78.125 -35.695 -77.945 ;
        RECT -37.905 -78.205 -37.400 -78.125 ;
        RECT -36.600 -78.215 -35.695 -78.125 ;
      LAYER mcon ;
        RECT -37.715 -78.205 -37.545 -78.035 ;
        RECT -36.350 -78.205 -36.180 -78.035 ;
      LAYER met1 ;
        RECT -37.600 -77.940 -36.600 -77.240 ;
        RECT -37.780 -78.240 -36.090 -77.940 ;
    END
  END o_ranQ[140]
  PIN o_ranQ[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -42.865 -83.935 -42.360 -83.855 ;
        RECT -41.560 -83.935 -40.655 -83.845 ;
        RECT -42.865 -84.115 -40.655 -83.935 ;
      LAYER mcon ;
        RECT -42.675 -84.025 -42.505 -83.855 ;
        RECT -41.310 -84.025 -41.140 -83.855 ;
      LAYER met1 ;
        RECT -42.740 -84.120 -41.050 -83.820 ;
        RECT -42.560 -84.820 -41.560 -84.120 ;
    END
  END o_ranQ[141]
  PIN o_ranQ[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -47.825 -78.125 -45.615 -77.945 ;
        RECT -47.825 -78.205 -47.320 -78.125 ;
        RECT -46.520 -78.215 -45.615 -78.125 ;
      LAYER mcon ;
        RECT -47.635 -78.205 -47.465 -78.035 ;
        RECT -46.270 -78.205 -46.100 -78.035 ;
      LAYER met1 ;
        RECT -47.520 -77.940 -46.520 -77.240 ;
        RECT -47.700 -78.240 -46.010 -77.940 ;
    END
  END o_ranQ[142]
  PIN o_ranQ[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -52.785 -83.935 -52.280 -83.855 ;
        RECT -51.480 -83.935 -50.575 -83.845 ;
        RECT -52.785 -84.115 -50.575 -83.935 ;
      LAYER mcon ;
        RECT -52.595 -84.025 -52.425 -83.855 ;
        RECT -51.230 -84.025 -51.060 -83.855 ;
      LAYER met1 ;
        RECT -52.660 -84.120 -50.970 -83.820 ;
        RECT -52.480 -84.820 -51.480 -84.120 ;
    END
  END o_ranQ[143]
  PIN o_ranQ[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -62.705 -83.935 -62.200 -83.855 ;
        RECT -61.400 -83.935 -60.495 -83.845 ;
        RECT -62.705 -84.115 -60.495 -83.935 ;
      LAYER mcon ;
        RECT -62.515 -84.025 -62.345 -83.855 ;
        RECT -61.150 -84.025 -60.980 -83.855 ;
      LAYER met1 ;
        RECT -62.580 -84.120 -60.890 -83.820 ;
        RECT -62.400 -84.820 -61.400 -84.120 ;
    END
  END o_ranQ[145]
  PIN o_ranQ[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -67.665 -78.125 -65.455 -77.945 ;
        RECT -67.665 -78.205 -67.160 -78.125 ;
        RECT -66.360 -78.215 -65.455 -78.125 ;
      LAYER mcon ;
        RECT -67.475 -78.205 -67.305 -78.035 ;
        RECT -66.110 -78.205 -65.940 -78.035 ;
      LAYER met1 ;
        RECT -67.360 -77.940 -66.360 -77.240 ;
        RECT -67.540 -78.240 -65.850 -77.940 ;
    END
  END o_ranQ[146]
  PIN o_ranQ[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -72.625 -83.935 -72.120 -83.855 ;
        RECT -71.320 -83.935 -70.415 -83.845 ;
        RECT -72.625 -84.115 -70.415 -83.935 ;
      LAYER mcon ;
        RECT -72.435 -84.025 -72.265 -83.855 ;
        RECT -71.070 -84.025 -70.900 -83.855 ;
      LAYER met1 ;
        RECT -72.500 -84.120 -70.810 -83.820 ;
        RECT -72.320 -84.820 -71.320 -84.120 ;
    END
  END o_ranQ[147]
  PIN o_ranQ[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -57.745 -78.125 -55.535 -77.945 ;
        RECT -57.745 -78.205 -57.240 -78.125 ;
        RECT -56.440 -78.215 -55.535 -78.125 ;
      LAYER mcon ;
        RECT -57.555 -78.205 -57.385 -78.035 ;
        RECT -56.190 -78.205 -56.020 -78.035 ;
      LAYER met1 ;
        RECT -57.440 -77.940 -56.440 -77.240 ;
        RECT -57.620 -78.240 -55.930 -77.940 ;
    END
  END o_ranQ[144]
  PIN o_ranQ[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -77.585 -78.125 -75.375 -77.945 ;
        RECT -77.585 -78.205 -77.080 -78.125 ;
        RECT -76.280 -78.215 -75.375 -78.125 ;
      LAYER mcon ;
        RECT -77.395 -78.205 -77.225 -78.035 ;
        RECT -76.030 -78.205 -75.860 -78.035 ;
      LAYER met1 ;
        RECT -77.280 -77.940 -76.280 -77.240 ;
        RECT -77.460 -78.240 -75.770 -77.940 ;
    END
  END o_ranQ[148]
  PIN o_ranQ[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -82.545 -83.935 -82.040 -83.855 ;
        RECT -81.240 -83.935 -80.335 -83.845 ;
        RECT -82.545 -84.115 -80.335 -83.935 ;
      LAYER mcon ;
        RECT -82.355 -84.025 -82.185 -83.855 ;
        RECT -80.990 -84.025 -80.820 -83.855 ;
      LAYER met1 ;
        RECT -82.420 -84.120 -80.730 -83.820 ;
        RECT -82.240 -84.820 -81.240 -84.120 ;
    END
  END o_ranQ[149]
  PIN o_ranQ[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -87.505 -78.125 -85.295 -77.945 ;
        RECT -87.505 -78.205 -87.000 -78.125 ;
        RECT -86.200 -78.215 -85.295 -78.125 ;
      LAYER mcon ;
        RECT -87.315 -78.205 -87.145 -78.035 ;
        RECT -85.950 -78.205 -85.780 -78.035 ;
      LAYER met1 ;
        RECT -87.200 -77.940 -86.200 -77.240 ;
        RECT -87.380 -78.240 -85.690 -77.940 ;
    END
  END o_ranQ[150]
  PIN o_ranQ[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -92.465 -83.935 -91.960 -83.855 ;
        RECT -91.160 -83.935 -90.255 -83.845 ;
        RECT -92.465 -84.115 -90.255 -83.935 ;
      LAYER mcon ;
        RECT -92.275 -84.025 -92.105 -83.855 ;
        RECT -90.910 -84.025 -90.740 -83.855 ;
      LAYER met1 ;
        RECT -92.340 -84.120 -90.650 -83.820 ;
        RECT -92.160 -84.820 -91.160 -84.120 ;
    END
  END o_ranQ[151]
  PIN o_ranQ[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -97.425 -78.125 -95.215 -77.945 ;
        RECT -97.425 -78.205 -96.920 -78.125 ;
        RECT -96.120 -78.215 -95.215 -78.125 ;
      LAYER mcon ;
        RECT -97.235 -78.205 -97.065 -78.035 ;
        RECT -95.870 -78.205 -95.700 -78.035 ;
      LAYER met1 ;
        RECT -97.120 -77.940 -96.120 -77.240 ;
        RECT -97.300 -78.240 -95.610 -77.940 ;
    END
  END o_ranQ[152]
  PIN o_ranQ[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -102.385 -83.935 -101.880 -83.855 ;
        RECT -101.080 -83.935 -100.175 -83.845 ;
        RECT -102.385 -84.115 -100.175 -83.935 ;
      LAYER mcon ;
        RECT -102.195 -84.025 -102.025 -83.855 ;
        RECT -100.830 -84.025 -100.660 -83.855 ;
      LAYER met1 ;
        RECT -102.260 -84.120 -100.570 -83.820 ;
        RECT -102.080 -84.820 -101.080 -84.120 ;
    END
  END o_ranQ[153]
  PIN o_ranQ[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -107.345 -78.125 -105.135 -77.945 ;
        RECT -107.345 -78.205 -106.840 -78.125 ;
        RECT -106.040 -78.215 -105.135 -78.125 ;
      LAYER mcon ;
        RECT -107.155 -78.205 -106.985 -78.035 ;
        RECT -105.790 -78.205 -105.620 -78.035 ;
      LAYER met1 ;
        RECT -107.040 -77.940 -106.040 -77.240 ;
        RECT -107.220 -78.240 -105.530 -77.940 ;
    END
  END o_ranQ[154]
  PIN o_ranQ[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -112.305 -83.935 -111.800 -83.855 ;
        RECT -111.000 -83.935 -110.095 -83.845 ;
        RECT -112.305 -84.115 -110.095 -83.935 ;
      LAYER mcon ;
        RECT -112.115 -84.025 -111.945 -83.855 ;
        RECT -110.750 -84.025 -110.580 -83.855 ;
      LAYER met1 ;
        RECT -112.180 -84.120 -110.490 -83.820 ;
        RECT -112.000 -84.820 -111.000 -84.120 ;
    END
  END o_ranQ[155]
  PIN o_ranQ[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -117.265 -78.125 -115.055 -77.945 ;
        RECT -117.265 -78.205 -116.760 -78.125 ;
        RECT -115.960 -78.215 -115.055 -78.125 ;
      LAYER mcon ;
        RECT -117.075 -78.205 -116.905 -78.035 ;
        RECT -115.710 -78.205 -115.540 -78.035 ;
      LAYER met1 ;
        RECT -116.960 -77.940 -115.960 -77.240 ;
        RECT -117.140 -78.240 -115.450 -77.940 ;
    END
  END o_ranQ[156]
  PIN o_ranQ[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -122.225 -83.935 -121.720 -83.855 ;
        RECT -120.920 -83.935 -120.015 -83.845 ;
        RECT -122.225 -84.115 -120.015 -83.935 ;
      LAYER mcon ;
        RECT -122.035 -84.025 -121.865 -83.855 ;
        RECT -120.670 -84.025 -120.500 -83.855 ;
      LAYER met1 ;
        RECT -122.100 -84.120 -120.410 -83.820 ;
        RECT -121.920 -84.820 -120.920 -84.120 ;
    END
  END o_ranQ[157]
  PIN o_ranQ[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -127.185 -78.125 -124.975 -77.945 ;
        RECT -127.185 -78.205 -126.680 -78.125 ;
        RECT -125.880 -78.215 -124.975 -78.125 ;
      LAYER mcon ;
        RECT -126.995 -78.205 -126.825 -78.035 ;
        RECT -125.630 -78.205 -125.460 -78.035 ;
      LAYER met1 ;
        RECT -126.880 -77.940 -125.880 -77.240 ;
        RECT -127.060 -78.240 -125.370 -77.940 ;
    END
  END o_ranQ[158]
  PIN o_ranQ[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -132.145 -83.935 -131.640 -83.855 ;
        RECT -130.840 -83.935 -129.935 -83.845 ;
        RECT -132.145 -84.115 -129.935 -83.935 ;
      LAYER mcon ;
        RECT -131.955 -84.025 -131.785 -83.855 ;
        RECT -130.590 -84.025 -130.420 -83.855 ;
      LAYER met1 ;
        RECT -132.020 -84.120 -130.330 -83.820 ;
        RECT -131.840 -84.820 -130.840 -84.120 ;
    END
  END o_ranQ[159]
  PIN o_ranQ[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -142.065 -83.935 -141.560 -83.855 ;
        RECT -140.760 -83.935 -139.855 -83.845 ;
        RECT -142.065 -84.115 -139.855 -83.935 ;
      LAYER mcon ;
        RECT -141.875 -84.025 -141.705 -83.855 ;
        RECT -140.510 -84.025 -140.340 -83.855 ;
      LAYER met1 ;
        RECT -141.940 -84.120 -140.250 -83.820 ;
        RECT -141.760 -84.820 -140.760 -84.120 ;
    END
  END o_ranQ[161]
  PIN o_ranQ[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -147.025 -78.125 -144.815 -77.945 ;
        RECT -147.025 -78.205 -146.520 -78.125 ;
        RECT -145.720 -78.215 -144.815 -78.125 ;
      LAYER mcon ;
        RECT -146.835 -78.205 -146.665 -78.035 ;
        RECT -145.470 -78.205 -145.300 -78.035 ;
      LAYER met1 ;
        RECT -146.720 -77.940 -145.720 -77.240 ;
        RECT -146.900 -78.240 -145.210 -77.940 ;
    END
  END o_ranQ[162]
  PIN o_ranQ[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -151.985 -83.935 -151.480 -83.855 ;
        RECT -150.680 -83.935 -149.775 -83.845 ;
        RECT -151.985 -84.115 -149.775 -83.935 ;
      LAYER mcon ;
        RECT -151.795 -84.025 -151.625 -83.855 ;
        RECT -150.430 -84.025 -150.260 -83.855 ;
      LAYER met1 ;
        RECT -151.860 -84.120 -150.170 -83.820 ;
        RECT -151.680 -84.820 -150.680 -84.120 ;
    END
  END o_ranQ[163]
  PIN o_ranQ[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -137.105 -78.125 -134.895 -77.945 ;
        RECT -137.105 -78.205 -136.600 -78.125 ;
        RECT -135.800 -78.215 -134.895 -78.125 ;
      LAYER mcon ;
        RECT -136.915 -78.205 -136.745 -78.035 ;
        RECT -135.550 -78.205 -135.380 -78.035 ;
      LAYER met1 ;
        RECT -136.800 -77.940 -135.800 -77.240 ;
        RECT -136.980 -78.240 -135.290 -77.940 ;
    END
  END o_ranQ[160]
  PIN o_ranQ[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -156.945 -78.125 -154.735 -77.945 ;
        RECT -156.945 -78.205 -156.440 -78.125 ;
        RECT -155.640 -78.215 -154.735 -78.125 ;
      LAYER mcon ;
        RECT -156.755 -78.205 -156.585 -78.035 ;
        RECT -155.390 -78.205 -155.220 -78.035 ;
      LAYER met1 ;
        RECT -156.640 -77.940 -155.640 -77.240 ;
        RECT -156.820 -78.240 -155.130 -77.940 ;
    END
  END o_ranQ[164]
  PIN o_ranQ[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -161.905 -83.935 -161.400 -83.855 ;
        RECT -160.600 -83.935 -159.695 -83.845 ;
        RECT -161.905 -84.115 -159.695 -83.935 ;
      LAYER mcon ;
        RECT -161.715 -84.025 -161.545 -83.855 ;
        RECT -160.350 -84.025 -160.180 -83.855 ;
      LAYER met1 ;
        RECT -161.780 -84.120 -160.090 -83.820 ;
        RECT -161.600 -84.820 -160.600 -84.120 ;
    END
  END o_ranQ[165]
  PIN o_ranQ[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -166.865 -78.125 -164.655 -77.945 ;
        RECT -166.865 -78.205 -166.360 -78.125 ;
        RECT -165.560 -78.215 -164.655 -78.125 ;
      LAYER mcon ;
        RECT -166.675 -78.205 -166.505 -78.035 ;
        RECT -165.310 -78.205 -165.140 -78.035 ;
      LAYER met1 ;
        RECT -166.560 -77.940 -165.560 -77.240 ;
        RECT -166.740 -78.240 -165.050 -77.940 ;
    END
  END o_ranQ[166]
  PIN o_ranQ[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -171.825 -83.935 -171.320 -83.855 ;
        RECT -170.520 -83.935 -169.615 -83.845 ;
        RECT -171.825 -84.115 -169.615 -83.935 ;
      LAYER mcon ;
        RECT -171.635 -84.025 -171.465 -83.855 ;
        RECT -170.270 -84.025 -170.100 -83.855 ;
      LAYER met1 ;
        RECT -171.700 -84.120 -170.010 -83.820 ;
        RECT -171.520 -84.820 -170.520 -84.120 ;
    END
  END o_ranQ[167]
  PIN o_ranQ[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -176.785 -78.125 -174.575 -77.945 ;
        RECT -176.785 -78.205 -176.280 -78.125 ;
        RECT -175.480 -78.215 -174.575 -78.125 ;
      LAYER mcon ;
        RECT -176.595 -78.205 -176.425 -78.035 ;
        RECT -175.230 -78.205 -175.060 -78.035 ;
      LAYER met1 ;
        RECT -176.480 -77.940 -175.480 -77.240 ;
        RECT -176.660 -78.240 -174.970 -77.940 ;
    END
  END o_ranQ[168]
  PIN o_ranQ[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -181.745 -83.935 -181.240 -83.855 ;
        RECT -180.440 -83.935 -179.535 -83.845 ;
        RECT -181.745 -84.115 -179.535 -83.935 ;
      LAYER mcon ;
        RECT -181.555 -84.025 -181.385 -83.855 ;
        RECT -180.190 -84.025 -180.020 -83.855 ;
      LAYER met1 ;
        RECT -181.620 -84.120 -179.930 -83.820 ;
        RECT -181.440 -84.820 -180.440 -84.120 ;
    END
  END o_ranQ[169]
  PIN o_ranQ[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -186.705 -78.125 -184.495 -77.945 ;
        RECT -186.705 -78.205 -186.200 -78.125 ;
        RECT -185.400 -78.215 -184.495 -78.125 ;
      LAYER mcon ;
        RECT -186.515 -78.205 -186.345 -78.035 ;
        RECT -185.150 -78.205 -184.980 -78.035 ;
      LAYER met1 ;
        RECT -186.400 -77.940 -185.400 -77.240 ;
        RECT -186.580 -78.240 -184.890 -77.940 ;
    END
  END o_ranQ[170]
  PIN o_ranQ[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -191.665 -83.935 -191.160 -83.855 ;
        RECT -190.360 -83.935 -189.455 -83.845 ;
        RECT -191.665 -84.115 -189.455 -83.935 ;
      LAYER mcon ;
        RECT -191.475 -84.025 -191.305 -83.855 ;
        RECT -190.110 -84.025 -189.940 -83.855 ;
      LAYER met1 ;
        RECT -191.540 -84.120 -189.850 -83.820 ;
        RECT -191.360 -84.820 -190.360 -84.120 ;
    END
  END o_ranQ[171]
  PIN o_ranQ[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -196.625 -78.125 -194.415 -77.945 ;
        RECT -196.625 -78.205 -196.120 -78.125 ;
        RECT -195.320 -78.215 -194.415 -78.125 ;
      LAYER mcon ;
        RECT -196.435 -78.205 -196.265 -78.035 ;
        RECT -195.070 -78.205 -194.900 -78.035 ;
      LAYER met1 ;
        RECT -196.320 -77.940 -195.320 -77.240 ;
        RECT -196.500 -78.240 -194.810 -77.940 ;
    END
  END o_ranQ[172]
  PIN o_ranQ[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -201.585 -83.935 -201.080 -83.855 ;
        RECT -200.280 -83.935 -199.375 -83.845 ;
        RECT -201.585 -84.115 -199.375 -83.935 ;
      LAYER mcon ;
        RECT -201.395 -84.025 -201.225 -83.855 ;
        RECT -200.030 -84.025 -199.860 -83.855 ;
      LAYER met1 ;
        RECT -201.460 -84.120 -199.770 -83.820 ;
        RECT -201.280 -84.820 -200.280 -84.120 ;
    END
  END o_ranQ[173]
  PIN o_ranQ[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -206.545 -78.125 -204.335 -77.945 ;
        RECT -206.545 -78.205 -206.040 -78.125 ;
        RECT -205.240 -78.215 -204.335 -78.125 ;
      LAYER mcon ;
        RECT -206.355 -78.205 -206.185 -78.035 ;
        RECT -204.990 -78.205 -204.820 -78.035 ;
      LAYER met1 ;
        RECT -206.240 -77.940 -205.240 -77.240 ;
        RECT -206.420 -78.240 -204.730 -77.940 ;
    END
  END o_ranQ[174]
  PIN o_ranQ[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -211.505 -83.935 -211.000 -83.855 ;
        RECT -210.200 -83.935 -209.295 -83.845 ;
        RECT -211.505 -84.115 -209.295 -83.935 ;
      LAYER mcon ;
        RECT -211.315 -84.025 -211.145 -83.855 ;
        RECT -209.950 -84.025 -209.780 -83.855 ;
      LAYER met1 ;
        RECT -211.380 -84.120 -209.690 -83.820 ;
        RECT -211.200 -84.820 -210.200 -84.120 ;
    END
  END o_ranQ[175]
  PIN o_ranQ[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -221.425 -83.935 -220.920 -83.855 ;
        RECT -220.120 -83.935 -219.215 -83.845 ;
        RECT -221.425 -84.115 -219.215 -83.935 ;
      LAYER mcon ;
        RECT -221.235 -84.025 -221.065 -83.855 ;
        RECT -219.870 -84.025 -219.700 -83.855 ;
      LAYER met1 ;
        RECT -221.300 -84.120 -219.610 -83.820 ;
        RECT -221.120 -84.820 -220.120 -84.120 ;
    END
  END o_ranQ[177]
  PIN o_ranQ[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -226.385 -78.125 -224.175 -77.945 ;
        RECT -226.385 -78.205 -225.880 -78.125 ;
        RECT -225.080 -78.215 -224.175 -78.125 ;
      LAYER mcon ;
        RECT -226.195 -78.205 -226.025 -78.035 ;
        RECT -224.830 -78.205 -224.660 -78.035 ;
      LAYER met1 ;
        RECT -226.080 -77.940 -225.080 -77.240 ;
        RECT -226.260 -78.240 -224.570 -77.940 ;
    END
  END o_ranQ[178]
  PIN o_ranQ[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -231.345 -83.935 -230.840 -83.855 ;
        RECT -230.040 -83.935 -229.135 -83.845 ;
        RECT -231.345 -84.115 -229.135 -83.935 ;
      LAYER mcon ;
        RECT -231.155 -84.025 -230.985 -83.855 ;
        RECT -229.790 -84.025 -229.620 -83.855 ;
      LAYER met1 ;
        RECT -231.220 -84.120 -229.530 -83.820 ;
        RECT -231.040 -84.820 -230.040 -84.120 ;
    END
  END o_ranQ[179]
  PIN o_ranQ[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -216.465 -78.125 -214.255 -77.945 ;
        RECT -216.465 -78.205 -215.960 -78.125 ;
        RECT -215.160 -78.215 -214.255 -78.125 ;
      LAYER mcon ;
        RECT -216.275 -78.205 -216.105 -78.035 ;
        RECT -214.910 -78.205 -214.740 -78.035 ;
      LAYER met1 ;
        RECT -216.160 -77.940 -215.160 -77.240 ;
        RECT -216.340 -78.240 -214.650 -77.940 ;
    END
  END o_ranQ[176]
  PIN o_ranQ[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -236.305 -78.125 -234.095 -77.945 ;
        RECT -236.305 -78.205 -235.800 -78.125 ;
        RECT -235.000 -78.215 -234.095 -78.125 ;
      LAYER mcon ;
        RECT -236.115 -78.205 -235.945 -78.035 ;
        RECT -234.750 -78.205 -234.580 -78.035 ;
      LAYER met1 ;
        RECT -236.000 -77.940 -235.000 -77.240 ;
        RECT -236.180 -78.240 -234.490 -77.940 ;
    END
  END o_ranQ[180]
  PIN o_ranQ[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -241.265 -83.935 -240.760 -83.855 ;
        RECT -239.960 -83.935 -239.055 -83.845 ;
        RECT -241.265 -84.115 -239.055 -83.935 ;
      LAYER mcon ;
        RECT -241.075 -84.025 -240.905 -83.855 ;
        RECT -239.710 -84.025 -239.540 -83.855 ;
      LAYER met1 ;
        RECT -241.140 -84.120 -239.450 -83.820 ;
        RECT -240.960 -84.820 -239.960 -84.120 ;
    END
  END o_ranQ[181]
  PIN o_ranQ[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -246.225 -78.125 -244.015 -77.945 ;
        RECT -246.225 -78.205 -245.720 -78.125 ;
        RECT -244.920 -78.215 -244.015 -78.125 ;
      LAYER mcon ;
        RECT -246.035 -78.205 -245.865 -78.035 ;
        RECT -244.670 -78.205 -244.500 -78.035 ;
      LAYER met1 ;
        RECT -245.920 -77.940 -244.920 -77.240 ;
        RECT -246.100 -78.240 -244.410 -77.940 ;
    END
  END o_ranQ[182]
  PIN o_ranQ[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -251.185 -83.935 -250.680 -83.855 ;
        RECT -249.880 -83.935 -248.975 -83.845 ;
        RECT -251.185 -84.115 -248.975 -83.935 ;
      LAYER mcon ;
        RECT -250.995 -84.025 -250.825 -83.855 ;
        RECT -249.630 -84.025 -249.460 -83.855 ;
      LAYER met1 ;
        RECT -251.060 -84.120 -249.370 -83.820 ;
        RECT -250.880 -84.820 -249.880 -84.120 ;
    END
  END o_ranQ[183]
  PIN o_ranQ[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -256.145 -78.125 -253.935 -77.945 ;
        RECT -256.145 -78.205 -255.640 -78.125 ;
        RECT -254.840 -78.215 -253.935 -78.125 ;
      LAYER mcon ;
        RECT -255.955 -78.205 -255.785 -78.035 ;
        RECT -254.590 -78.205 -254.420 -78.035 ;
      LAYER met1 ;
        RECT -255.840 -77.940 -254.840 -77.240 ;
        RECT -256.020 -78.240 -254.330 -77.940 ;
    END
  END o_ranQ[184]
  PIN o_ranQ[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -261.105 -83.935 -260.600 -83.855 ;
        RECT -259.800 -83.935 -258.895 -83.845 ;
        RECT -261.105 -84.115 -258.895 -83.935 ;
      LAYER mcon ;
        RECT -260.915 -84.025 -260.745 -83.855 ;
        RECT -259.550 -84.025 -259.380 -83.855 ;
      LAYER met1 ;
        RECT -260.980 -84.120 -259.290 -83.820 ;
        RECT -260.800 -84.820 -259.800 -84.120 ;
    END
  END o_ranQ[185]
  PIN o_ranQ[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -266.065 -78.125 -263.855 -77.945 ;
        RECT -266.065 -78.205 -265.560 -78.125 ;
        RECT -264.760 -78.215 -263.855 -78.125 ;
      LAYER mcon ;
        RECT -265.875 -78.205 -265.705 -78.035 ;
        RECT -264.510 -78.205 -264.340 -78.035 ;
      LAYER met1 ;
        RECT -265.760 -77.940 -264.760 -77.240 ;
        RECT -265.940 -78.240 -264.250 -77.940 ;
    END
  END o_ranQ[186]
  PIN o_ranQ[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -271.025 -83.935 -270.520 -83.855 ;
        RECT -269.720 -83.935 -268.815 -83.845 ;
        RECT -271.025 -84.115 -268.815 -83.935 ;
      LAYER mcon ;
        RECT -270.835 -84.025 -270.665 -83.855 ;
        RECT -269.470 -84.025 -269.300 -83.855 ;
      LAYER met1 ;
        RECT -270.900 -84.120 -269.210 -83.820 ;
        RECT -270.720 -84.820 -269.720 -84.120 ;
    END
  END o_ranQ[187]
  PIN o_ranQ[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -275.985 -78.125 -273.775 -77.945 ;
        RECT -275.985 -78.205 -275.480 -78.125 ;
        RECT -274.680 -78.215 -273.775 -78.125 ;
      LAYER mcon ;
        RECT -275.795 -78.205 -275.625 -78.035 ;
        RECT -274.430 -78.205 -274.260 -78.035 ;
      LAYER met1 ;
        RECT -275.680 -77.940 -274.680 -77.240 ;
        RECT -275.860 -78.240 -274.170 -77.940 ;
    END
  END o_ranQ[188]
  PIN o_ranQ[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -280.945 -83.935 -280.440 -83.855 ;
        RECT -279.640 -83.935 -278.735 -83.845 ;
        RECT -280.945 -84.115 -278.735 -83.935 ;
      LAYER mcon ;
        RECT -280.755 -84.025 -280.585 -83.855 ;
        RECT -279.390 -84.025 -279.220 -83.855 ;
      LAYER met1 ;
        RECT -280.820 -84.120 -279.130 -83.820 ;
        RECT -280.640 -84.820 -279.640 -84.120 ;
    END
  END o_ranQ[189]
  PIN o_ranQ[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -285.905 -78.125 -283.695 -77.945 ;
        RECT -285.905 -78.205 -285.400 -78.125 ;
        RECT -284.600 -78.215 -283.695 -78.125 ;
      LAYER mcon ;
        RECT -285.715 -78.205 -285.545 -78.035 ;
        RECT -284.350 -78.205 -284.180 -78.035 ;
      LAYER met1 ;
        RECT -285.600 -77.940 -284.600 -77.240 ;
        RECT -285.780 -78.240 -284.090 -77.940 ;
    END
  END o_ranQ[190]
  PIN o_ranQ[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -290.865 -83.935 -290.360 -83.855 ;
        RECT -289.560 -83.935 -288.655 -83.845 ;
        RECT -290.865 -84.115 -288.655 -83.935 ;
      LAYER mcon ;
        RECT -290.675 -84.025 -290.505 -83.855 ;
        RECT -289.310 -84.025 -289.140 -83.855 ;
      LAYER met1 ;
        RECT -290.740 -84.120 -289.050 -83.820 ;
        RECT -290.560 -84.820 -289.560 -84.120 ;
    END
  END o_ranQ[191]
  PIN o_ranQ[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 14.895 -178.515 15.400 -178.435 ;
        RECT 16.200 -178.515 17.105 -178.425 ;
        RECT 14.895 -178.695 17.105 -178.515 ;
      LAYER mcon ;
        RECT 15.085 -178.605 15.255 -178.435 ;
        RECT 16.450 -178.605 16.620 -178.435 ;
      LAYER met1 ;
        RECT 15.020 -178.700 16.710 -178.400 ;
        RECT 15.200 -179.400 16.200 -178.700 ;
    END
  END o_ranQ[193]
  PIN o_ranQ[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 9.935 -172.705 12.145 -172.525 ;
        RECT 9.935 -172.785 10.440 -172.705 ;
        RECT 11.240 -172.795 12.145 -172.705 ;
      LAYER mcon ;
        RECT 10.125 -172.785 10.295 -172.615 ;
        RECT 11.490 -172.785 11.660 -172.615 ;
      LAYER met1 ;
        RECT 10.240 -172.520 11.240 -171.820 ;
        RECT 10.060 -172.820 11.750 -172.520 ;
    END
  END o_ranQ[194]
  PIN o_ranQ[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 4.975 -178.515 5.480 -178.435 ;
        RECT 6.280 -178.515 7.185 -178.425 ;
        RECT 4.975 -178.695 7.185 -178.515 ;
      LAYER mcon ;
        RECT 5.165 -178.605 5.335 -178.435 ;
        RECT 6.530 -178.605 6.700 -178.435 ;
      LAYER met1 ;
        RECT 5.100 -178.700 6.790 -178.400 ;
        RECT 5.280 -179.400 6.280 -178.700 ;
    END
  END o_ranQ[195]
  PIN o_ranQ[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 19.855 -172.705 22.065 -172.525 ;
        RECT 19.855 -172.785 20.360 -172.705 ;
        RECT 21.160 -172.795 22.065 -172.705 ;
      LAYER mcon ;
        RECT 20.045 -172.785 20.215 -172.615 ;
        RECT 21.410 -172.785 21.580 -172.615 ;
      LAYER met1 ;
        RECT 20.160 -172.520 21.160 -171.820 ;
        RECT 19.980 -172.820 21.670 -172.520 ;
    END
  END o_ranQ[192]
  PIN o_ranQ[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 0.015 -172.705 2.225 -172.525 ;
        RECT 0.015 -172.785 0.520 -172.705 ;
        RECT 1.320 -172.795 2.225 -172.705 ;
      LAYER mcon ;
        RECT 0.205 -172.785 0.375 -172.615 ;
        RECT 1.570 -172.785 1.740 -172.615 ;
      LAYER met1 ;
        RECT 0.320 -172.520 1.320 -171.820 ;
        RECT 0.140 -172.820 1.830 -172.520 ;
    END
  END o_ranQ[196]
  PIN o_ranQ[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -4.945 -178.515 -4.440 -178.435 ;
        RECT -3.640 -178.515 -2.735 -178.425 ;
        RECT -4.945 -178.695 -2.735 -178.515 ;
      LAYER mcon ;
        RECT -4.755 -178.605 -4.585 -178.435 ;
        RECT -3.390 -178.605 -3.220 -178.435 ;
      LAYER met1 ;
        RECT -4.820 -178.700 -3.130 -178.400 ;
        RECT -4.640 -179.400 -3.640 -178.700 ;
    END
  END o_ranQ[197]
  PIN o_ranQ[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -9.905 -172.705 -7.695 -172.525 ;
        RECT -9.905 -172.785 -9.400 -172.705 ;
        RECT -8.600 -172.795 -7.695 -172.705 ;
      LAYER mcon ;
        RECT -9.715 -172.785 -9.545 -172.615 ;
        RECT -8.350 -172.785 -8.180 -172.615 ;
      LAYER met1 ;
        RECT -9.600 -172.520 -8.600 -171.820 ;
        RECT -9.780 -172.820 -8.090 -172.520 ;
    END
  END o_ranQ[198]
  PIN o_ranQ[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -14.865 -178.515 -14.360 -178.435 ;
        RECT -13.560 -178.515 -12.655 -178.425 ;
        RECT -14.865 -178.695 -12.655 -178.515 ;
      LAYER mcon ;
        RECT -14.675 -178.605 -14.505 -178.435 ;
        RECT -13.310 -178.605 -13.140 -178.435 ;
      LAYER met1 ;
        RECT -14.740 -178.700 -13.050 -178.400 ;
        RECT -14.560 -179.400 -13.560 -178.700 ;
    END
  END o_ranQ[199]
  PIN o_ranQ[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -19.825 -172.705 -17.615 -172.525 ;
        RECT -19.825 -172.785 -19.320 -172.705 ;
        RECT -18.520 -172.795 -17.615 -172.705 ;
      LAYER mcon ;
        RECT -19.635 -172.785 -19.465 -172.615 ;
        RECT -18.270 -172.785 -18.100 -172.615 ;
      LAYER met1 ;
        RECT -19.520 -172.520 -18.520 -171.820 ;
        RECT -19.700 -172.820 -18.010 -172.520 ;
    END
  END o_ranQ[200]
  PIN o_ranQ[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -24.785 -178.515 -24.280 -178.435 ;
        RECT -23.480 -178.515 -22.575 -178.425 ;
        RECT -24.785 -178.695 -22.575 -178.515 ;
      LAYER mcon ;
        RECT -24.595 -178.605 -24.425 -178.435 ;
        RECT -23.230 -178.605 -23.060 -178.435 ;
      LAYER met1 ;
        RECT -24.660 -178.700 -22.970 -178.400 ;
        RECT -24.480 -179.400 -23.480 -178.700 ;
    END
  END o_ranQ[201]
  PIN o_ranQ[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -29.745 -172.705 -27.535 -172.525 ;
        RECT -29.745 -172.785 -29.240 -172.705 ;
        RECT -28.440 -172.795 -27.535 -172.705 ;
      LAYER mcon ;
        RECT -29.555 -172.785 -29.385 -172.615 ;
        RECT -28.190 -172.785 -28.020 -172.615 ;
      LAYER met1 ;
        RECT -29.440 -172.520 -28.440 -171.820 ;
        RECT -29.620 -172.820 -27.930 -172.520 ;
    END
  END o_ranQ[202]
  PIN o_ranQ[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -34.705 -178.515 -34.200 -178.435 ;
        RECT -33.400 -178.515 -32.495 -178.425 ;
        RECT -34.705 -178.695 -32.495 -178.515 ;
      LAYER mcon ;
        RECT -34.515 -178.605 -34.345 -178.435 ;
        RECT -33.150 -178.605 -32.980 -178.435 ;
      LAYER met1 ;
        RECT -34.580 -178.700 -32.890 -178.400 ;
        RECT -34.400 -179.400 -33.400 -178.700 ;
    END
  END o_ranQ[203]
  PIN o_ranQ[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -39.665 -172.705 -37.455 -172.525 ;
        RECT -39.665 -172.785 -39.160 -172.705 ;
        RECT -38.360 -172.795 -37.455 -172.705 ;
      LAYER mcon ;
        RECT -39.475 -172.785 -39.305 -172.615 ;
        RECT -38.110 -172.785 -37.940 -172.615 ;
      LAYER met1 ;
        RECT -39.360 -172.520 -38.360 -171.820 ;
        RECT -39.540 -172.820 -37.850 -172.520 ;
    END
  END o_ranQ[204]
  PIN o_ranQ[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -44.625 -178.515 -44.120 -178.435 ;
        RECT -43.320 -178.515 -42.415 -178.425 ;
        RECT -44.625 -178.695 -42.415 -178.515 ;
      LAYER mcon ;
        RECT -44.435 -178.605 -44.265 -178.435 ;
        RECT -43.070 -178.605 -42.900 -178.435 ;
      LAYER met1 ;
        RECT -44.500 -178.700 -42.810 -178.400 ;
        RECT -44.320 -179.400 -43.320 -178.700 ;
    END
  END o_ranQ[205]
  PIN o_ranQ[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -49.585 -172.705 -47.375 -172.525 ;
        RECT -49.585 -172.785 -49.080 -172.705 ;
        RECT -48.280 -172.795 -47.375 -172.705 ;
      LAYER mcon ;
        RECT -49.395 -172.785 -49.225 -172.615 ;
        RECT -48.030 -172.785 -47.860 -172.615 ;
      LAYER met1 ;
        RECT -49.280 -172.520 -48.280 -171.820 ;
        RECT -49.460 -172.820 -47.770 -172.520 ;
    END
  END o_ranQ[206]
  PIN o_ranQ[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -54.545 -178.515 -54.040 -178.435 ;
        RECT -53.240 -178.515 -52.335 -178.425 ;
        RECT -54.545 -178.695 -52.335 -178.515 ;
      LAYER mcon ;
        RECT -54.355 -178.605 -54.185 -178.435 ;
        RECT -52.990 -178.605 -52.820 -178.435 ;
      LAYER met1 ;
        RECT -54.420 -178.700 -52.730 -178.400 ;
        RECT -54.240 -179.400 -53.240 -178.700 ;
    END
  END o_ranQ[207]
  PIN o_ranQ[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -64.465 -178.515 -63.960 -178.435 ;
        RECT -63.160 -178.515 -62.255 -178.425 ;
        RECT -64.465 -178.695 -62.255 -178.515 ;
      LAYER mcon ;
        RECT -64.275 -178.605 -64.105 -178.435 ;
        RECT -62.910 -178.605 -62.740 -178.435 ;
      LAYER met1 ;
        RECT -64.340 -178.700 -62.650 -178.400 ;
        RECT -64.160 -179.400 -63.160 -178.700 ;
    END
  END o_ranQ[209]
  PIN o_ranQ[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -69.425 -172.705 -67.215 -172.525 ;
        RECT -69.425 -172.785 -68.920 -172.705 ;
        RECT -68.120 -172.795 -67.215 -172.705 ;
      LAYER mcon ;
        RECT -69.235 -172.785 -69.065 -172.615 ;
        RECT -67.870 -172.785 -67.700 -172.615 ;
      LAYER met1 ;
        RECT -69.120 -172.520 -68.120 -171.820 ;
        RECT -69.300 -172.820 -67.610 -172.520 ;
    END
  END o_ranQ[210]
  PIN o_ranQ[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -74.385 -178.515 -73.880 -178.435 ;
        RECT -73.080 -178.515 -72.175 -178.425 ;
        RECT -74.385 -178.695 -72.175 -178.515 ;
      LAYER mcon ;
        RECT -74.195 -178.605 -74.025 -178.435 ;
        RECT -72.830 -178.605 -72.660 -178.435 ;
      LAYER met1 ;
        RECT -74.260 -178.700 -72.570 -178.400 ;
        RECT -74.080 -179.400 -73.080 -178.700 ;
    END
  END o_ranQ[211]
  PIN o_ranQ[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -59.505 -172.705 -57.295 -172.525 ;
        RECT -59.505 -172.785 -59.000 -172.705 ;
        RECT -58.200 -172.795 -57.295 -172.705 ;
      LAYER mcon ;
        RECT -59.315 -172.785 -59.145 -172.615 ;
        RECT -57.950 -172.785 -57.780 -172.615 ;
      LAYER met1 ;
        RECT -59.200 -172.520 -58.200 -171.820 ;
        RECT -59.380 -172.820 -57.690 -172.520 ;
    END
  END o_ranQ[208]
  PIN o_ranQ[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -79.345 -172.705 -77.135 -172.525 ;
        RECT -79.345 -172.785 -78.840 -172.705 ;
        RECT -78.040 -172.795 -77.135 -172.705 ;
      LAYER mcon ;
        RECT -79.155 -172.785 -78.985 -172.615 ;
        RECT -77.790 -172.785 -77.620 -172.615 ;
      LAYER met1 ;
        RECT -79.040 -172.520 -78.040 -171.820 ;
        RECT -79.220 -172.820 -77.530 -172.520 ;
    END
  END o_ranQ[212]
  PIN o_ranQ[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -84.305 -178.515 -83.800 -178.435 ;
        RECT -83.000 -178.515 -82.095 -178.425 ;
        RECT -84.305 -178.695 -82.095 -178.515 ;
      LAYER mcon ;
        RECT -84.115 -178.605 -83.945 -178.435 ;
        RECT -82.750 -178.605 -82.580 -178.435 ;
      LAYER met1 ;
        RECT -84.180 -178.700 -82.490 -178.400 ;
        RECT -84.000 -179.400 -83.000 -178.700 ;
    END
  END o_ranQ[213]
  PIN o_ranQ[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -89.265 -172.705 -87.055 -172.525 ;
        RECT -89.265 -172.785 -88.760 -172.705 ;
        RECT -87.960 -172.795 -87.055 -172.705 ;
      LAYER mcon ;
        RECT -89.075 -172.785 -88.905 -172.615 ;
        RECT -87.710 -172.785 -87.540 -172.615 ;
      LAYER met1 ;
        RECT -88.960 -172.520 -87.960 -171.820 ;
        RECT -89.140 -172.820 -87.450 -172.520 ;
    END
  END o_ranQ[214]
  PIN o_ranQ[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -94.225 -178.515 -93.720 -178.435 ;
        RECT -92.920 -178.515 -92.015 -178.425 ;
        RECT -94.225 -178.695 -92.015 -178.515 ;
      LAYER mcon ;
        RECT -94.035 -178.605 -93.865 -178.435 ;
        RECT -92.670 -178.605 -92.500 -178.435 ;
      LAYER met1 ;
        RECT -94.100 -178.700 -92.410 -178.400 ;
        RECT -93.920 -179.400 -92.920 -178.700 ;
    END
  END o_ranQ[215]
  PIN o_ranQ[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -99.185 -172.705 -96.975 -172.525 ;
        RECT -99.185 -172.785 -98.680 -172.705 ;
        RECT -97.880 -172.795 -96.975 -172.705 ;
      LAYER mcon ;
        RECT -98.995 -172.785 -98.825 -172.615 ;
        RECT -97.630 -172.785 -97.460 -172.615 ;
      LAYER met1 ;
        RECT -98.880 -172.520 -97.880 -171.820 ;
        RECT -99.060 -172.820 -97.370 -172.520 ;
    END
  END o_ranQ[216]
  PIN o_ranQ[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -104.145 -178.515 -103.640 -178.435 ;
        RECT -102.840 -178.515 -101.935 -178.425 ;
        RECT -104.145 -178.695 -101.935 -178.515 ;
      LAYER mcon ;
        RECT -103.955 -178.605 -103.785 -178.435 ;
        RECT -102.590 -178.605 -102.420 -178.435 ;
      LAYER met1 ;
        RECT -104.020 -178.700 -102.330 -178.400 ;
        RECT -103.840 -179.400 -102.840 -178.700 ;
    END
  END o_ranQ[217]
  PIN o_ranQ[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -109.105 -172.705 -106.895 -172.525 ;
        RECT -109.105 -172.785 -108.600 -172.705 ;
        RECT -107.800 -172.795 -106.895 -172.705 ;
      LAYER mcon ;
        RECT -108.915 -172.785 -108.745 -172.615 ;
        RECT -107.550 -172.785 -107.380 -172.615 ;
      LAYER met1 ;
        RECT -108.800 -172.520 -107.800 -171.820 ;
        RECT -108.980 -172.820 -107.290 -172.520 ;
    END
  END o_ranQ[218]
  PIN o_ranQ[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -114.065 -178.515 -113.560 -178.435 ;
        RECT -112.760 -178.515 -111.855 -178.425 ;
        RECT -114.065 -178.695 -111.855 -178.515 ;
      LAYER mcon ;
        RECT -113.875 -178.605 -113.705 -178.435 ;
        RECT -112.510 -178.605 -112.340 -178.435 ;
      LAYER met1 ;
        RECT -113.940 -178.700 -112.250 -178.400 ;
        RECT -113.760 -179.400 -112.760 -178.700 ;
    END
  END o_ranQ[219]
  PIN o_ranQ[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -119.025 -172.705 -116.815 -172.525 ;
        RECT -119.025 -172.785 -118.520 -172.705 ;
        RECT -117.720 -172.795 -116.815 -172.705 ;
      LAYER mcon ;
        RECT -118.835 -172.785 -118.665 -172.615 ;
        RECT -117.470 -172.785 -117.300 -172.615 ;
      LAYER met1 ;
        RECT -118.720 -172.520 -117.720 -171.820 ;
        RECT -118.900 -172.820 -117.210 -172.520 ;
    END
  END o_ranQ[220]
  PIN o_ranQ[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -123.985 -178.515 -123.480 -178.435 ;
        RECT -122.680 -178.515 -121.775 -178.425 ;
        RECT -123.985 -178.695 -121.775 -178.515 ;
      LAYER mcon ;
        RECT -123.795 -178.605 -123.625 -178.435 ;
        RECT -122.430 -178.605 -122.260 -178.435 ;
      LAYER met1 ;
        RECT -123.860 -178.700 -122.170 -178.400 ;
        RECT -123.680 -179.400 -122.680 -178.700 ;
    END
  END o_ranQ[221]
  PIN o_ranQ[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -128.945 -172.705 -126.735 -172.525 ;
        RECT -128.945 -172.785 -128.440 -172.705 ;
        RECT -127.640 -172.795 -126.735 -172.705 ;
      LAYER mcon ;
        RECT -128.755 -172.785 -128.585 -172.615 ;
        RECT -127.390 -172.785 -127.220 -172.615 ;
      LAYER met1 ;
        RECT -128.640 -172.520 -127.640 -171.820 ;
        RECT -128.820 -172.820 -127.130 -172.520 ;
    END
  END o_ranQ[222]
  PIN o_ranQ[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -133.905 -178.515 -133.400 -178.435 ;
        RECT -132.600 -178.515 -131.695 -178.425 ;
        RECT -133.905 -178.695 -131.695 -178.515 ;
      LAYER mcon ;
        RECT -133.715 -178.605 -133.545 -178.435 ;
        RECT -132.350 -178.605 -132.180 -178.435 ;
      LAYER met1 ;
        RECT -133.780 -178.700 -132.090 -178.400 ;
        RECT -133.600 -179.400 -132.600 -178.700 ;
    END
  END o_ranQ[223]
  PIN o_ranQ[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -143.825 -178.515 -143.320 -178.435 ;
        RECT -142.520 -178.515 -141.615 -178.425 ;
        RECT -143.825 -178.695 -141.615 -178.515 ;
      LAYER mcon ;
        RECT -143.635 -178.605 -143.465 -178.435 ;
        RECT -142.270 -178.605 -142.100 -178.435 ;
      LAYER met1 ;
        RECT -143.700 -178.700 -142.010 -178.400 ;
        RECT -143.520 -179.400 -142.520 -178.700 ;
    END
  END o_ranQ[225]
  PIN o_ranQ[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -148.785 -172.705 -146.575 -172.525 ;
        RECT -148.785 -172.785 -148.280 -172.705 ;
        RECT -147.480 -172.795 -146.575 -172.705 ;
      LAYER mcon ;
        RECT -148.595 -172.785 -148.425 -172.615 ;
        RECT -147.230 -172.785 -147.060 -172.615 ;
      LAYER met1 ;
        RECT -148.480 -172.520 -147.480 -171.820 ;
        RECT -148.660 -172.820 -146.970 -172.520 ;
    END
  END o_ranQ[226]
  PIN o_ranQ[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -153.745 -178.515 -153.240 -178.435 ;
        RECT -152.440 -178.515 -151.535 -178.425 ;
        RECT -153.745 -178.695 -151.535 -178.515 ;
      LAYER mcon ;
        RECT -153.555 -178.605 -153.385 -178.435 ;
        RECT -152.190 -178.605 -152.020 -178.435 ;
      LAYER met1 ;
        RECT -153.620 -178.700 -151.930 -178.400 ;
        RECT -153.440 -179.400 -152.440 -178.700 ;
    END
  END o_ranQ[227]
  PIN o_ranQ[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -138.865 -172.705 -136.655 -172.525 ;
        RECT -138.865 -172.785 -138.360 -172.705 ;
        RECT -137.560 -172.795 -136.655 -172.705 ;
      LAYER mcon ;
        RECT -138.675 -172.785 -138.505 -172.615 ;
        RECT -137.310 -172.785 -137.140 -172.615 ;
      LAYER met1 ;
        RECT -138.560 -172.520 -137.560 -171.820 ;
        RECT -138.740 -172.820 -137.050 -172.520 ;
    END
  END o_ranQ[224]
  PIN o_ranQ[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -158.705 -172.705 -156.495 -172.525 ;
        RECT -158.705 -172.785 -158.200 -172.705 ;
        RECT -157.400 -172.795 -156.495 -172.705 ;
      LAYER mcon ;
        RECT -158.515 -172.785 -158.345 -172.615 ;
        RECT -157.150 -172.785 -156.980 -172.615 ;
      LAYER met1 ;
        RECT -158.400 -172.520 -157.400 -171.820 ;
        RECT -158.580 -172.820 -156.890 -172.520 ;
    END
  END o_ranQ[228]
  PIN o_ranQ[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -163.665 -178.515 -163.160 -178.435 ;
        RECT -162.360 -178.515 -161.455 -178.425 ;
        RECT -163.665 -178.695 -161.455 -178.515 ;
      LAYER mcon ;
        RECT -163.475 -178.605 -163.305 -178.435 ;
        RECT -162.110 -178.605 -161.940 -178.435 ;
      LAYER met1 ;
        RECT -163.540 -178.700 -161.850 -178.400 ;
        RECT -163.360 -179.400 -162.360 -178.700 ;
    END
  END o_ranQ[229]
  PIN o_ranQ[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -168.625 -172.705 -166.415 -172.525 ;
        RECT -168.625 -172.785 -168.120 -172.705 ;
        RECT -167.320 -172.795 -166.415 -172.705 ;
      LAYER mcon ;
        RECT -168.435 -172.785 -168.265 -172.615 ;
        RECT -167.070 -172.785 -166.900 -172.615 ;
      LAYER met1 ;
        RECT -168.320 -172.520 -167.320 -171.820 ;
        RECT -168.500 -172.820 -166.810 -172.520 ;
    END
  END o_ranQ[230]
  PIN o_ranQ[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -173.585 -178.515 -173.080 -178.435 ;
        RECT -172.280 -178.515 -171.375 -178.425 ;
        RECT -173.585 -178.695 -171.375 -178.515 ;
      LAYER mcon ;
        RECT -173.395 -178.605 -173.225 -178.435 ;
        RECT -172.030 -178.605 -171.860 -178.435 ;
      LAYER met1 ;
        RECT -173.460 -178.700 -171.770 -178.400 ;
        RECT -173.280 -179.400 -172.280 -178.700 ;
    END
  END o_ranQ[231]
  PIN o_ranQ[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -178.545 -172.705 -176.335 -172.525 ;
        RECT -178.545 -172.785 -178.040 -172.705 ;
        RECT -177.240 -172.795 -176.335 -172.705 ;
      LAYER mcon ;
        RECT -178.355 -172.785 -178.185 -172.615 ;
        RECT -176.990 -172.785 -176.820 -172.615 ;
      LAYER met1 ;
        RECT -178.240 -172.520 -177.240 -171.820 ;
        RECT -178.420 -172.820 -176.730 -172.520 ;
    END
  END o_ranQ[232]
  PIN o_ranQ[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -183.505 -178.515 -183.000 -178.435 ;
        RECT -182.200 -178.515 -181.295 -178.425 ;
        RECT -183.505 -178.695 -181.295 -178.515 ;
      LAYER mcon ;
        RECT -183.315 -178.605 -183.145 -178.435 ;
        RECT -181.950 -178.605 -181.780 -178.435 ;
      LAYER met1 ;
        RECT -183.380 -178.700 -181.690 -178.400 ;
        RECT -183.200 -179.400 -182.200 -178.700 ;
    END
  END o_ranQ[233]
  PIN o_ranQ[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -188.465 -172.705 -186.255 -172.525 ;
        RECT -188.465 -172.785 -187.960 -172.705 ;
        RECT -187.160 -172.795 -186.255 -172.705 ;
      LAYER mcon ;
        RECT -188.275 -172.785 -188.105 -172.615 ;
        RECT -186.910 -172.785 -186.740 -172.615 ;
      LAYER met1 ;
        RECT -188.160 -172.520 -187.160 -171.820 ;
        RECT -188.340 -172.820 -186.650 -172.520 ;
    END
  END o_ranQ[234]
  PIN o_ranQ[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -193.425 -178.515 -192.920 -178.435 ;
        RECT -192.120 -178.515 -191.215 -178.425 ;
        RECT -193.425 -178.695 -191.215 -178.515 ;
      LAYER mcon ;
        RECT -193.235 -178.605 -193.065 -178.435 ;
        RECT -191.870 -178.605 -191.700 -178.435 ;
      LAYER met1 ;
        RECT -193.300 -178.700 -191.610 -178.400 ;
        RECT -193.120 -179.400 -192.120 -178.700 ;
    END
  END o_ranQ[235]
  PIN o_ranQ[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -198.385 -172.705 -196.175 -172.525 ;
        RECT -198.385 -172.785 -197.880 -172.705 ;
        RECT -197.080 -172.795 -196.175 -172.705 ;
      LAYER mcon ;
        RECT -198.195 -172.785 -198.025 -172.615 ;
        RECT -196.830 -172.785 -196.660 -172.615 ;
      LAYER met1 ;
        RECT -198.080 -172.520 -197.080 -171.820 ;
        RECT -198.260 -172.820 -196.570 -172.520 ;
    END
  END o_ranQ[236]
  PIN o_ranQ[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -203.345 -178.515 -202.840 -178.435 ;
        RECT -202.040 -178.515 -201.135 -178.425 ;
        RECT -203.345 -178.695 -201.135 -178.515 ;
      LAYER mcon ;
        RECT -203.155 -178.605 -202.985 -178.435 ;
        RECT -201.790 -178.605 -201.620 -178.435 ;
      LAYER met1 ;
        RECT -203.220 -178.700 -201.530 -178.400 ;
        RECT -203.040 -179.400 -202.040 -178.700 ;
    END
  END o_ranQ[237]
  PIN o_ranQ[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -208.305 -172.705 -206.095 -172.525 ;
        RECT -208.305 -172.785 -207.800 -172.705 ;
        RECT -207.000 -172.795 -206.095 -172.705 ;
      LAYER mcon ;
        RECT -208.115 -172.785 -207.945 -172.615 ;
        RECT -206.750 -172.785 -206.580 -172.615 ;
      LAYER met1 ;
        RECT -208.000 -172.520 -207.000 -171.820 ;
        RECT -208.180 -172.820 -206.490 -172.520 ;
    END
  END o_ranQ[238]
  PIN o_ranQ[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -213.265 -178.515 -212.760 -178.435 ;
        RECT -211.960 -178.515 -211.055 -178.425 ;
        RECT -213.265 -178.695 -211.055 -178.515 ;
      LAYER mcon ;
        RECT -213.075 -178.605 -212.905 -178.435 ;
        RECT -211.710 -178.605 -211.540 -178.435 ;
      LAYER met1 ;
        RECT -213.140 -178.700 -211.450 -178.400 ;
        RECT -212.960 -179.400 -211.960 -178.700 ;
    END
  END o_ranQ[239]
  PIN o_ranQ[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -223.185 -178.515 -222.680 -178.435 ;
        RECT -221.880 -178.515 -220.975 -178.425 ;
        RECT -223.185 -178.695 -220.975 -178.515 ;
      LAYER mcon ;
        RECT -222.995 -178.605 -222.825 -178.435 ;
        RECT -221.630 -178.605 -221.460 -178.435 ;
      LAYER met1 ;
        RECT -223.060 -178.700 -221.370 -178.400 ;
        RECT -222.880 -179.400 -221.880 -178.700 ;
    END
  END o_ranQ[241]
  PIN o_ranQ[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -228.145 -172.705 -225.935 -172.525 ;
        RECT -228.145 -172.785 -227.640 -172.705 ;
        RECT -226.840 -172.795 -225.935 -172.705 ;
      LAYER mcon ;
        RECT -227.955 -172.785 -227.785 -172.615 ;
        RECT -226.590 -172.785 -226.420 -172.615 ;
      LAYER met1 ;
        RECT -227.840 -172.520 -226.840 -171.820 ;
        RECT -228.020 -172.820 -226.330 -172.520 ;
    END
  END o_ranQ[242]
  PIN o_ranQ[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -233.105 -178.515 -232.600 -178.435 ;
        RECT -231.800 -178.515 -230.895 -178.425 ;
        RECT -233.105 -178.695 -230.895 -178.515 ;
      LAYER mcon ;
        RECT -232.915 -178.605 -232.745 -178.435 ;
        RECT -231.550 -178.605 -231.380 -178.435 ;
      LAYER met1 ;
        RECT -232.980 -178.700 -231.290 -178.400 ;
        RECT -232.800 -179.400 -231.800 -178.700 ;
    END
  END o_ranQ[243]
  PIN o_ranQ[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -218.225 -172.705 -216.015 -172.525 ;
        RECT -218.225 -172.785 -217.720 -172.705 ;
        RECT -216.920 -172.795 -216.015 -172.705 ;
      LAYER mcon ;
        RECT -218.035 -172.785 -217.865 -172.615 ;
        RECT -216.670 -172.785 -216.500 -172.615 ;
      LAYER met1 ;
        RECT -217.920 -172.520 -216.920 -171.820 ;
        RECT -218.100 -172.820 -216.410 -172.520 ;
    END
  END o_ranQ[240]
  PIN o_ranQ[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -238.065 -172.705 -235.855 -172.525 ;
        RECT -238.065 -172.785 -237.560 -172.705 ;
        RECT -236.760 -172.795 -235.855 -172.705 ;
      LAYER mcon ;
        RECT -237.875 -172.785 -237.705 -172.615 ;
        RECT -236.510 -172.785 -236.340 -172.615 ;
      LAYER met1 ;
        RECT -237.760 -172.520 -236.760 -171.820 ;
        RECT -237.940 -172.820 -236.250 -172.520 ;
    END
  END o_ranQ[244]
  PIN o_ranQ[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -243.025 -178.515 -242.520 -178.435 ;
        RECT -241.720 -178.515 -240.815 -178.425 ;
        RECT -243.025 -178.695 -240.815 -178.515 ;
      LAYER mcon ;
        RECT -242.835 -178.605 -242.665 -178.435 ;
        RECT -241.470 -178.605 -241.300 -178.435 ;
      LAYER met1 ;
        RECT -242.900 -178.700 -241.210 -178.400 ;
        RECT -242.720 -179.400 -241.720 -178.700 ;
    END
  END o_ranQ[245]
  PIN o_ranQ[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -247.985 -172.705 -245.775 -172.525 ;
        RECT -247.985 -172.785 -247.480 -172.705 ;
        RECT -246.680 -172.795 -245.775 -172.705 ;
      LAYER mcon ;
        RECT -247.795 -172.785 -247.625 -172.615 ;
        RECT -246.430 -172.785 -246.260 -172.615 ;
      LAYER met1 ;
        RECT -247.680 -172.520 -246.680 -171.820 ;
        RECT -247.860 -172.820 -246.170 -172.520 ;
    END
  END o_ranQ[246]
  PIN o_ranQ[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -252.945 -178.515 -252.440 -178.435 ;
        RECT -251.640 -178.515 -250.735 -178.425 ;
        RECT -252.945 -178.695 -250.735 -178.515 ;
      LAYER mcon ;
        RECT -252.755 -178.605 -252.585 -178.435 ;
        RECT -251.390 -178.605 -251.220 -178.435 ;
      LAYER met1 ;
        RECT -252.820 -178.700 -251.130 -178.400 ;
        RECT -252.640 -179.400 -251.640 -178.700 ;
    END
  END o_ranQ[247]
  PIN o_ranQ[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -257.905 -172.705 -255.695 -172.525 ;
        RECT -257.905 -172.785 -257.400 -172.705 ;
        RECT -256.600 -172.795 -255.695 -172.705 ;
      LAYER mcon ;
        RECT -257.715 -172.785 -257.545 -172.615 ;
        RECT -256.350 -172.785 -256.180 -172.615 ;
      LAYER met1 ;
        RECT -257.600 -172.520 -256.600 -171.820 ;
        RECT -257.780 -172.820 -256.090 -172.520 ;
    END
  END o_ranQ[248]
  PIN o_ranQ[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -262.865 -178.515 -262.360 -178.435 ;
        RECT -261.560 -178.515 -260.655 -178.425 ;
        RECT -262.865 -178.695 -260.655 -178.515 ;
      LAYER mcon ;
        RECT -262.675 -178.605 -262.505 -178.435 ;
        RECT -261.310 -178.605 -261.140 -178.435 ;
      LAYER met1 ;
        RECT -262.740 -178.700 -261.050 -178.400 ;
        RECT -262.560 -179.400 -261.560 -178.700 ;
    END
  END o_ranQ[249]
  PIN o_ranQ[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -267.825 -172.705 -265.615 -172.525 ;
        RECT -267.825 -172.785 -267.320 -172.705 ;
        RECT -266.520 -172.795 -265.615 -172.705 ;
      LAYER mcon ;
        RECT -267.635 -172.785 -267.465 -172.615 ;
        RECT -266.270 -172.785 -266.100 -172.615 ;
      LAYER met1 ;
        RECT -267.520 -172.520 -266.520 -171.820 ;
        RECT -267.700 -172.820 -266.010 -172.520 ;
    END
  END o_ranQ[250]
  PIN o_ranQ[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -272.785 -178.515 -272.280 -178.435 ;
        RECT -271.480 -178.515 -270.575 -178.425 ;
        RECT -272.785 -178.695 -270.575 -178.515 ;
      LAYER mcon ;
        RECT -272.595 -178.605 -272.425 -178.435 ;
        RECT -271.230 -178.605 -271.060 -178.435 ;
      LAYER met1 ;
        RECT -272.660 -178.700 -270.970 -178.400 ;
        RECT -272.480 -179.400 -271.480 -178.700 ;
    END
  END o_ranQ[251]
  PIN o_ranQ[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -277.745 -172.705 -275.535 -172.525 ;
        RECT -277.745 -172.785 -277.240 -172.705 ;
        RECT -276.440 -172.795 -275.535 -172.705 ;
      LAYER mcon ;
        RECT -277.555 -172.785 -277.385 -172.615 ;
        RECT -276.190 -172.785 -276.020 -172.615 ;
      LAYER met1 ;
        RECT -277.440 -172.520 -276.440 -171.820 ;
        RECT -277.620 -172.820 -275.930 -172.520 ;
    END
  END o_ranQ[252]
  PIN o_ranQ[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -282.705 -178.515 -282.200 -178.435 ;
        RECT -281.400 -178.515 -280.495 -178.425 ;
        RECT -282.705 -178.695 -280.495 -178.515 ;
      LAYER mcon ;
        RECT -282.515 -178.605 -282.345 -178.435 ;
        RECT -281.150 -178.605 -280.980 -178.435 ;
      LAYER met1 ;
        RECT -282.580 -178.700 -280.890 -178.400 ;
        RECT -282.400 -179.400 -281.400 -178.700 ;
    END
  END o_ranQ[253]
  PIN o_ranQ[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -287.665 -172.705 -285.455 -172.525 ;
        RECT -287.665 -172.785 -287.160 -172.705 ;
        RECT -286.360 -172.795 -285.455 -172.705 ;
      LAYER mcon ;
        RECT -287.475 -172.785 -287.305 -172.615 ;
        RECT -286.110 -172.785 -285.940 -172.615 ;
      LAYER met1 ;
        RECT -287.360 -172.520 -286.360 -171.820 ;
        RECT -287.540 -172.820 -285.850 -172.520 ;
    END
  END o_ranQ[254]
  PIN o_ranQ[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT -292.625 -178.515 -292.120 -178.435 ;
        RECT -291.320 -178.515 -290.415 -178.425 ;
        RECT -292.625 -178.695 -290.415 -178.515 ;
      LAYER mcon ;
        RECT -292.435 -178.605 -292.265 -178.435 ;
        RECT -291.070 -178.605 -290.900 -178.435 ;
      LAYER met1 ;
        RECT -292.500 -178.700 -290.810 -178.400 ;
        RECT -292.320 -179.400 -291.320 -178.700 ;
    END
  END o_ranQ[255]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -283.195 93.570 -279.425 95.330 ;
        RECT -273.275 93.570 -269.505 95.330 ;
        RECT -263.355 93.570 -259.585 95.330 ;
        RECT -253.435 93.570 -249.665 95.330 ;
        RECT -243.515 93.570 -239.745 95.330 ;
        RECT -233.595 93.570 -229.825 95.330 ;
        RECT -223.675 93.570 -219.905 95.330 ;
        RECT -213.755 93.570 -209.985 95.330 ;
        RECT -203.835 93.570 -200.065 95.330 ;
        RECT -193.915 93.570 -190.145 95.330 ;
        RECT -183.995 93.570 -180.225 95.330 ;
        RECT -174.075 93.570 -170.305 95.330 ;
        RECT -164.155 93.570 -160.385 95.330 ;
        RECT -154.235 93.570 -150.465 95.330 ;
        RECT -144.315 93.570 -140.545 95.330 ;
        RECT -134.395 93.570 -130.625 95.330 ;
        RECT -124.475 93.570 -120.705 95.330 ;
        RECT -114.555 93.570 -110.785 95.330 ;
        RECT -104.635 93.570 -100.865 95.330 ;
        RECT -94.715 93.570 -90.945 95.330 ;
        RECT -84.795 93.570 -81.025 95.330 ;
        RECT -74.875 93.570 -71.105 95.330 ;
        RECT -64.955 93.570 -61.185 95.330 ;
        RECT -55.035 93.570 -51.265 95.330 ;
        RECT -45.115 93.570 -41.345 95.330 ;
        RECT -35.195 93.570 -31.425 95.330 ;
        RECT -25.275 93.570 -21.505 95.330 ;
        RECT -15.355 93.570 -11.585 95.330 ;
        RECT -5.435 93.570 -1.665 95.330 ;
        RECT 4.485 93.570 8.255 95.330 ;
        RECT 14.405 93.570 18.175 95.330 ;
        RECT 24.325 95.095 25.930 95.330 ;
        RECT 24.325 95.090 26.440 95.095 ;
        RECT 24.325 93.570 26.630 95.090 ;
        RECT -281.730 93.520 -280.890 93.570 ;
        RECT -288.070 91.915 -284.470 93.520 ;
        RECT -283.110 90.420 -279.510 92.025 ;
        RECT -278.150 91.915 -274.550 93.520 ;
        RECT -271.810 93.510 -270.970 93.570 ;
        RECT -261.890 93.520 -261.050 93.570 ;
        RECT -273.190 90.420 -269.590 92.025 ;
        RECT -268.230 91.915 -264.630 93.520 ;
        RECT -263.270 90.420 -259.670 92.025 ;
        RECT -258.310 91.915 -254.710 93.520 ;
        RECT -251.970 93.510 -251.130 93.570 ;
        RECT -242.050 93.520 -241.210 93.570 ;
        RECT -253.350 90.420 -249.750 92.025 ;
        RECT -248.390 91.915 -244.790 93.520 ;
        RECT -243.430 90.420 -239.830 92.025 ;
        RECT -238.470 91.915 -234.870 93.520 ;
        RECT -232.130 93.510 -231.290 93.570 ;
        RECT -222.210 93.520 -221.370 93.570 ;
        RECT -233.510 90.420 -229.910 92.025 ;
        RECT -228.550 91.915 -224.950 93.520 ;
        RECT -223.590 90.420 -219.990 92.025 ;
        RECT -218.630 91.915 -215.030 93.520 ;
        RECT -212.290 93.510 -211.450 93.570 ;
        RECT -202.370 93.520 -201.530 93.570 ;
        RECT -213.670 90.420 -210.070 92.025 ;
        RECT -208.710 91.915 -205.110 93.520 ;
        RECT -203.750 90.420 -200.150 92.025 ;
        RECT -198.790 91.915 -195.190 93.520 ;
        RECT -192.450 93.510 -191.610 93.570 ;
        RECT -182.530 93.520 -181.690 93.570 ;
        RECT -193.830 90.420 -190.230 92.025 ;
        RECT -188.870 91.915 -185.270 93.520 ;
        RECT -183.910 90.420 -180.310 92.025 ;
        RECT -178.950 91.915 -175.350 93.520 ;
        RECT -172.610 93.510 -171.770 93.570 ;
        RECT -162.690 93.520 -161.850 93.570 ;
        RECT -173.990 90.420 -170.390 92.025 ;
        RECT -169.030 91.915 -165.430 93.520 ;
        RECT -164.070 90.420 -160.470 92.025 ;
        RECT -159.110 91.915 -155.510 93.520 ;
        RECT -152.770 93.510 -151.930 93.570 ;
        RECT -142.850 93.520 -142.010 93.570 ;
        RECT -154.150 90.420 -150.550 92.025 ;
        RECT -149.190 91.915 -145.590 93.520 ;
        RECT -144.230 90.420 -140.630 92.025 ;
        RECT -139.270 91.915 -135.670 93.520 ;
        RECT -132.930 93.510 -132.090 93.570 ;
        RECT -123.010 93.520 -122.170 93.570 ;
        RECT -134.310 90.420 -130.710 92.025 ;
        RECT -129.350 91.915 -125.750 93.520 ;
        RECT -124.390 90.420 -120.790 92.025 ;
        RECT -119.430 91.915 -115.830 93.520 ;
        RECT -113.090 93.510 -112.250 93.570 ;
        RECT -103.170 93.520 -102.330 93.570 ;
        RECT -114.470 90.420 -110.870 92.025 ;
        RECT -109.510 91.915 -105.910 93.520 ;
        RECT -104.550 90.420 -100.950 92.025 ;
        RECT -99.590 91.915 -95.990 93.520 ;
        RECT -93.250 93.510 -92.410 93.570 ;
        RECT -83.330 93.520 -82.490 93.570 ;
        RECT -94.630 90.420 -91.030 92.025 ;
        RECT -89.670 91.915 -86.070 93.520 ;
        RECT -84.710 90.420 -81.110 92.025 ;
        RECT -79.750 91.915 -76.150 93.520 ;
        RECT -73.410 93.510 -72.570 93.570 ;
        RECT -63.490 93.520 -62.650 93.570 ;
        RECT -74.790 90.420 -71.190 92.025 ;
        RECT -69.830 91.915 -66.230 93.520 ;
        RECT -64.870 90.420 -61.270 92.025 ;
        RECT -59.910 91.915 -56.310 93.520 ;
        RECT -53.570 93.510 -52.730 93.570 ;
        RECT -43.650 93.520 -42.810 93.570 ;
        RECT -54.950 90.420 -51.350 92.025 ;
        RECT -49.990 91.915 -46.390 93.520 ;
        RECT -45.030 90.420 -41.430 92.025 ;
        RECT -40.070 91.915 -36.470 93.520 ;
        RECT -33.730 93.510 -32.890 93.570 ;
        RECT -23.810 93.520 -22.970 93.570 ;
        RECT -35.110 90.420 -31.510 92.025 ;
        RECT -30.150 91.915 -26.550 93.520 ;
        RECT -25.190 90.420 -21.590 92.025 ;
        RECT -20.230 91.915 -16.630 93.520 ;
        RECT -13.890 93.510 -13.050 93.570 ;
        RECT -3.970 93.520 -3.130 93.570 ;
        RECT -15.270 90.420 -11.670 92.025 ;
        RECT -10.310 91.915 -6.710 93.520 ;
        RECT -5.350 90.420 -1.750 92.025 ;
        RECT -0.390 91.915 3.210 93.520 ;
        RECT 5.950 93.510 6.790 93.570 ;
        RECT 15.870 93.520 16.710 93.570 ;
        RECT 25.790 93.520 26.630 93.570 ;
        RECT 4.570 90.420 8.170 92.025 ;
        RECT 9.530 91.915 13.130 93.520 ;
        RECT 14.490 90.420 18.090 92.025 ;
        RECT 19.450 91.915 23.050 93.520 ;
        RECT 24.410 90.420 26.630 92.025 ;
        RECT -288.155 88.610 -284.385 90.370 ;
        RECT -278.235 88.610 -274.465 90.370 ;
        RECT -268.315 88.610 -264.545 90.370 ;
        RECT -258.395 88.610 -254.625 90.370 ;
        RECT -248.475 88.610 -244.705 90.370 ;
        RECT -238.555 88.610 -234.785 90.370 ;
        RECT -228.635 88.610 -224.865 90.370 ;
        RECT -218.715 88.610 -214.945 90.370 ;
        RECT -208.795 88.610 -205.025 90.370 ;
        RECT -198.875 88.610 -195.105 90.370 ;
        RECT -188.955 88.610 -185.185 90.370 ;
        RECT -179.035 88.610 -175.265 90.370 ;
        RECT -169.115 88.610 -165.345 90.370 ;
        RECT -159.195 88.610 -155.425 90.370 ;
        RECT -149.275 88.610 -145.505 90.370 ;
        RECT -139.355 88.610 -135.585 90.370 ;
        RECT -129.435 88.610 -125.665 90.370 ;
        RECT -119.515 88.610 -115.745 90.370 ;
        RECT -109.595 88.610 -105.825 90.370 ;
        RECT -99.675 88.610 -95.905 90.370 ;
        RECT -89.755 88.610 -85.985 90.370 ;
        RECT -79.835 88.610 -76.065 90.370 ;
        RECT -69.915 88.610 -66.145 90.370 ;
        RECT -59.995 88.610 -56.225 90.370 ;
        RECT -50.075 88.610 -46.305 90.370 ;
        RECT -40.155 88.610 -36.385 90.370 ;
        RECT -30.235 88.610 -26.465 90.370 ;
        RECT -20.315 88.610 -16.545 90.370 ;
        RECT -10.395 88.610 -6.625 90.370 ;
        RECT -0.475 88.610 3.295 90.370 ;
        RECT 9.445 88.610 13.215 90.370 ;
        RECT 19.365 88.610 23.135 90.370 ;
        RECT -285.215 9.520 -281.445 11.280 ;
        RECT -275.295 9.520 -271.525 11.280 ;
        RECT -265.375 9.520 -261.605 11.280 ;
        RECT -255.455 9.520 -251.685 11.280 ;
        RECT -245.535 9.520 -241.765 11.280 ;
        RECT -235.615 9.520 -231.845 11.280 ;
        RECT -225.695 9.520 -221.925 11.280 ;
        RECT -215.775 9.520 -212.005 11.280 ;
        RECT -205.855 9.520 -202.085 11.280 ;
        RECT -195.935 9.520 -192.165 11.280 ;
        RECT -186.015 9.520 -182.245 11.280 ;
        RECT -176.095 9.520 -172.325 11.280 ;
        RECT -166.175 9.520 -162.405 11.280 ;
        RECT -156.255 9.520 -152.485 11.280 ;
        RECT -146.335 9.520 -142.565 11.280 ;
        RECT -136.415 9.520 -132.645 11.280 ;
        RECT -126.495 9.520 -122.725 11.280 ;
        RECT -116.575 9.520 -112.805 11.280 ;
        RECT -106.655 9.520 -102.885 11.280 ;
        RECT -96.735 9.520 -92.965 11.280 ;
        RECT -86.815 9.520 -83.045 11.280 ;
        RECT -76.895 9.520 -73.125 11.280 ;
        RECT -66.975 9.520 -63.205 11.280 ;
        RECT -57.055 9.520 -53.285 11.280 ;
        RECT -47.135 9.520 -43.365 11.280 ;
        RECT -37.215 9.520 -33.445 11.280 ;
        RECT -27.295 9.520 -23.525 11.280 ;
        RECT -17.375 9.520 -13.605 11.280 ;
        RECT -7.455 9.520 -3.685 11.280 ;
        RECT 2.465 9.520 6.235 11.280 ;
        RECT 12.385 9.520 16.155 11.280 ;
        RECT 22.305 11.045 23.910 11.280 ;
        RECT 22.305 11.040 24.420 11.045 ;
        RECT 22.305 9.520 24.610 11.040 ;
        RECT -283.750 9.470 -282.910 9.520 ;
        RECT -290.090 7.865 -286.490 9.470 ;
        RECT -285.130 6.370 -281.530 7.975 ;
        RECT -280.170 7.865 -276.570 9.470 ;
        RECT -273.830 9.460 -272.990 9.520 ;
        RECT -263.910 9.470 -263.070 9.520 ;
        RECT -275.210 6.370 -271.610 7.975 ;
        RECT -270.250 7.865 -266.650 9.470 ;
        RECT -265.290 6.370 -261.690 7.975 ;
        RECT -260.330 7.865 -256.730 9.470 ;
        RECT -253.990 9.460 -253.150 9.520 ;
        RECT -244.070 9.470 -243.230 9.520 ;
        RECT -255.370 6.370 -251.770 7.975 ;
        RECT -250.410 7.865 -246.810 9.470 ;
        RECT -245.450 6.370 -241.850 7.975 ;
        RECT -240.490 7.865 -236.890 9.470 ;
        RECT -234.150 9.460 -233.310 9.520 ;
        RECT -224.230 9.470 -223.390 9.520 ;
        RECT -235.530 6.370 -231.930 7.975 ;
        RECT -230.570 7.865 -226.970 9.470 ;
        RECT -225.610 6.370 -222.010 7.975 ;
        RECT -220.650 7.865 -217.050 9.470 ;
        RECT -214.310 9.460 -213.470 9.520 ;
        RECT -204.390 9.470 -203.550 9.520 ;
        RECT -215.690 6.370 -212.090 7.975 ;
        RECT -210.730 7.865 -207.130 9.470 ;
        RECT -205.770 6.370 -202.170 7.975 ;
        RECT -200.810 7.865 -197.210 9.470 ;
        RECT -194.470 9.460 -193.630 9.520 ;
        RECT -184.550 9.470 -183.710 9.520 ;
        RECT -195.850 6.370 -192.250 7.975 ;
        RECT -190.890 7.865 -187.290 9.470 ;
        RECT -185.930 6.370 -182.330 7.975 ;
        RECT -180.970 7.865 -177.370 9.470 ;
        RECT -174.630 9.460 -173.790 9.520 ;
        RECT -164.710 9.470 -163.870 9.520 ;
        RECT -176.010 6.370 -172.410 7.975 ;
        RECT -171.050 7.865 -167.450 9.470 ;
        RECT -166.090 6.370 -162.490 7.975 ;
        RECT -161.130 7.865 -157.530 9.470 ;
        RECT -154.790 9.460 -153.950 9.520 ;
        RECT -144.870 9.470 -144.030 9.520 ;
        RECT -156.170 6.370 -152.570 7.975 ;
        RECT -151.210 7.865 -147.610 9.470 ;
        RECT -146.250 6.370 -142.650 7.975 ;
        RECT -141.290 7.865 -137.690 9.470 ;
        RECT -134.950 9.460 -134.110 9.520 ;
        RECT -125.030 9.470 -124.190 9.520 ;
        RECT -136.330 6.370 -132.730 7.975 ;
        RECT -131.370 7.865 -127.770 9.470 ;
        RECT -126.410 6.370 -122.810 7.975 ;
        RECT -121.450 7.865 -117.850 9.470 ;
        RECT -115.110 9.460 -114.270 9.520 ;
        RECT -105.190 9.470 -104.350 9.520 ;
        RECT -116.490 6.370 -112.890 7.975 ;
        RECT -111.530 7.865 -107.930 9.470 ;
        RECT -106.570 6.370 -102.970 7.975 ;
        RECT -101.610 7.865 -98.010 9.470 ;
        RECT -95.270 9.460 -94.430 9.520 ;
        RECT -85.350 9.470 -84.510 9.520 ;
        RECT -96.650 6.370 -93.050 7.975 ;
        RECT -91.690 7.865 -88.090 9.470 ;
        RECT -86.730 6.370 -83.130 7.975 ;
        RECT -81.770 7.865 -78.170 9.470 ;
        RECT -75.430 9.460 -74.590 9.520 ;
        RECT -65.510 9.470 -64.670 9.520 ;
        RECT -76.810 6.370 -73.210 7.975 ;
        RECT -71.850 7.865 -68.250 9.470 ;
        RECT -66.890 6.370 -63.290 7.975 ;
        RECT -61.930 7.865 -58.330 9.470 ;
        RECT -55.590 9.460 -54.750 9.520 ;
        RECT -45.670 9.470 -44.830 9.520 ;
        RECT -56.970 6.370 -53.370 7.975 ;
        RECT -52.010 7.865 -48.410 9.470 ;
        RECT -47.050 6.370 -43.450 7.975 ;
        RECT -42.090 7.865 -38.490 9.470 ;
        RECT -35.750 9.460 -34.910 9.520 ;
        RECT -25.830 9.470 -24.990 9.520 ;
        RECT -37.130 6.370 -33.530 7.975 ;
        RECT -32.170 7.865 -28.570 9.470 ;
        RECT -27.210 6.370 -23.610 7.975 ;
        RECT -22.250 7.865 -18.650 9.470 ;
        RECT -15.910 9.460 -15.070 9.520 ;
        RECT -5.990 9.470 -5.150 9.520 ;
        RECT -17.290 6.370 -13.690 7.975 ;
        RECT -12.330 7.865 -8.730 9.470 ;
        RECT -7.370 6.370 -3.770 7.975 ;
        RECT -2.410 7.865 1.190 9.470 ;
        RECT 3.930 9.460 4.770 9.520 ;
        RECT 13.850 9.470 14.690 9.520 ;
        RECT 23.770 9.470 24.610 9.520 ;
        RECT 2.550 6.370 6.150 7.975 ;
        RECT 7.510 7.865 11.110 9.470 ;
        RECT 12.470 6.370 16.070 7.975 ;
        RECT 17.430 7.865 21.030 9.470 ;
        RECT 22.390 6.370 24.610 7.975 ;
        RECT -290.175 4.560 -286.405 6.320 ;
        RECT -280.255 4.560 -276.485 6.320 ;
        RECT -270.335 4.560 -266.565 6.320 ;
        RECT -260.415 4.560 -256.645 6.320 ;
        RECT -250.495 4.560 -246.725 6.320 ;
        RECT -240.575 4.560 -236.805 6.320 ;
        RECT -230.655 4.560 -226.885 6.320 ;
        RECT -220.735 4.560 -216.965 6.320 ;
        RECT -210.815 4.560 -207.045 6.320 ;
        RECT -200.895 4.560 -197.125 6.320 ;
        RECT -190.975 4.560 -187.205 6.320 ;
        RECT -181.055 4.560 -177.285 6.320 ;
        RECT -171.135 4.560 -167.365 6.320 ;
        RECT -161.215 4.560 -157.445 6.320 ;
        RECT -151.295 4.560 -147.525 6.320 ;
        RECT -141.375 4.560 -137.605 6.320 ;
        RECT -131.455 4.560 -127.685 6.320 ;
        RECT -121.535 4.560 -117.765 6.320 ;
        RECT -111.615 4.560 -107.845 6.320 ;
        RECT -101.695 4.560 -97.925 6.320 ;
        RECT -91.775 4.560 -88.005 6.320 ;
        RECT -81.855 4.560 -78.085 6.320 ;
        RECT -71.935 4.560 -68.165 6.320 ;
        RECT -62.015 4.560 -58.245 6.320 ;
        RECT -52.095 4.560 -48.325 6.320 ;
        RECT -42.175 4.560 -38.405 6.320 ;
        RECT -32.255 4.560 -28.485 6.320 ;
        RECT -22.335 4.560 -18.565 6.320 ;
        RECT -12.415 4.560 -8.645 6.320 ;
        RECT -2.495 4.560 1.275 6.320 ;
        RECT 7.425 4.560 11.195 6.320 ;
        RECT 17.345 4.560 21.115 6.320 ;
        RECT -284.855 -79.430 -281.085 -77.670 ;
        RECT -274.935 -79.430 -271.165 -77.670 ;
        RECT -265.015 -79.430 -261.245 -77.670 ;
        RECT -255.095 -79.430 -251.325 -77.670 ;
        RECT -245.175 -79.430 -241.405 -77.670 ;
        RECT -235.255 -79.430 -231.485 -77.670 ;
        RECT -225.335 -79.430 -221.565 -77.670 ;
        RECT -215.415 -79.430 -211.645 -77.670 ;
        RECT -205.495 -79.430 -201.725 -77.670 ;
        RECT -195.575 -79.430 -191.805 -77.670 ;
        RECT -185.655 -79.430 -181.885 -77.670 ;
        RECT -175.735 -79.430 -171.965 -77.670 ;
        RECT -165.815 -79.430 -162.045 -77.670 ;
        RECT -155.895 -79.430 -152.125 -77.670 ;
        RECT -145.975 -79.430 -142.205 -77.670 ;
        RECT -136.055 -79.430 -132.285 -77.670 ;
        RECT -126.135 -79.430 -122.365 -77.670 ;
        RECT -116.215 -79.430 -112.445 -77.670 ;
        RECT -106.295 -79.430 -102.525 -77.670 ;
        RECT -96.375 -79.430 -92.605 -77.670 ;
        RECT -86.455 -79.430 -82.685 -77.670 ;
        RECT -76.535 -79.430 -72.765 -77.670 ;
        RECT -66.615 -79.430 -62.845 -77.670 ;
        RECT -56.695 -79.430 -52.925 -77.670 ;
        RECT -46.775 -79.430 -43.005 -77.670 ;
        RECT -36.855 -79.430 -33.085 -77.670 ;
        RECT -26.935 -79.430 -23.165 -77.670 ;
        RECT -17.015 -79.430 -13.245 -77.670 ;
        RECT -7.095 -79.430 -3.325 -77.670 ;
        RECT 2.825 -79.430 6.595 -77.670 ;
        RECT 12.745 -79.430 16.515 -77.670 ;
        RECT 22.665 -77.905 24.270 -77.670 ;
        RECT 22.665 -77.910 24.780 -77.905 ;
        RECT 22.665 -79.430 24.970 -77.910 ;
        RECT -283.390 -79.480 -282.550 -79.430 ;
        RECT -289.730 -81.085 -286.130 -79.480 ;
        RECT -284.770 -82.580 -281.170 -80.975 ;
        RECT -279.810 -81.085 -276.210 -79.480 ;
        RECT -273.470 -79.490 -272.630 -79.430 ;
        RECT -263.550 -79.480 -262.710 -79.430 ;
        RECT -274.850 -82.580 -271.250 -80.975 ;
        RECT -269.890 -81.085 -266.290 -79.480 ;
        RECT -264.930 -82.580 -261.330 -80.975 ;
        RECT -259.970 -81.085 -256.370 -79.480 ;
        RECT -253.630 -79.490 -252.790 -79.430 ;
        RECT -243.710 -79.480 -242.870 -79.430 ;
        RECT -255.010 -82.580 -251.410 -80.975 ;
        RECT -250.050 -81.085 -246.450 -79.480 ;
        RECT -245.090 -82.580 -241.490 -80.975 ;
        RECT -240.130 -81.085 -236.530 -79.480 ;
        RECT -233.790 -79.490 -232.950 -79.430 ;
        RECT -223.870 -79.480 -223.030 -79.430 ;
        RECT -235.170 -82.580 -231.570 -80.975 ;
        RECT -230.210 -81.085 -226.610 -79.480 ;
        RECT -225.250 -82.580 -221.650 -80.975 ;
        RECT -220.290 -81.085 -216.690 -79.480 ;
        RECT -213.950 -79.490 -213.110 -79.430 ;
        RECT -204.030 -79.480 -203.190 -79.430 ;
        RECT -215.330 -82.580 -211.730 -80.975 ;
        RECT -210.370 -81.085 -206.770 -79.480 ;
        RECT -205.410 -82.580 -201.810 -80.975 ;
        RECT -200.450 -81.085 -196.850 -79.480 ;
        RECT -194.110 -79.490 -193.270 -79.430 ;
        RECT -184.190 -79.480 -183.350 -79.430 ;
        RECT -195.490 -82.580 -191.890 -80.975 ;
        RECT -190.530 -81.085 -186.930 -79.480 ;
        RECT -185.570 -82.580 -181.970 -80.975 ;
        RECT -180.610 -81.085 -177.010 -79.480 ;
        RECT -174.270 -79.490 -173.430 -79.430 ;
        RECT -164.350 -79.480 -163.510 -79.430 ;
        RECT -175.650 -82.580 -172.050 -80.975 ;
        RECT -170.690 -81.085 -167.090 -79.480 ;
        RECT -165.730 -82.580 -162.130 -80.975 ;
        RECT -160.770 -81.085 -157.170 -79.480 ;
        RECT -154.430 -79.490 -153.590 -79.430 ;
        RECT -144.510 -79.480 -143.670 -79.430 ;
        RECT -155.810 -82.580 -152.210 -80.975 ;
        RECT -150.850 -81.085 -147.250 -79.480 ;
        RECT -145.890 -82.580 -142.290 -80.975 ;
        RECT -140.930 -81.085 -137.330 -79.480 ;
        RECT -134.590 -79.490 -133.750 -79.430 ;
        RECT -124.670 -79.480 -123.830 -79.430 ;
        RECT -135.970 -82.580 -132.370 -80.975 ;
        RECT -131.010 -81.085 -127.410 -79.480 ;
        RECT -126.050 -82.580 -122.450 -80.975 ;
        RECT -121.090 -81.085 -117.490 -79.480 ;
        RECT -114.750 -79.490 -113.910 -79.430 ;
        RECT -104.830 -79.480 -103.990 -79.430 ;
        RECT -116.130 -82.580 -112.530 -80.975 ;
        RECT -111.170 -81.085 -107.570 -79.480 ;
        RECT -106.210 -82.580 -102.610 -80.975 ;
        RECT -101.250 -81.085 -97.650 -79.480 ;
        RECT -94.910 -79.490 -94.070 -79.430 ;
        RECT -84.990 -79.480 -84.150 -79.430 ;
        RECT -96.290 -82.580 -92.690 -80.975 ;
        RECT -91.330 -81.085 -87.730 -79.480 ;
        RECT -86.370 -82.580 -82.770 -80.975 ;
        RECT -81.410 -81.085 -77.810 -79.480 ;
        RECT -75.070 -79.490 -74.230 -79.430 ;
        RECT -65.150 -79.480 -64.310 -79.430 ;
        RECT -76.450 -82.580 -72.850 -80.975 ;
        RECT -71.490 -81.085 -67.890 -79.480 ;
        RECT -66.530 -82.580 -62.930 -80.975 ;
        RECT -61.570 -81.085 -57.970 -79.480 ;
        RECT -55.230 -79.490 -54.390 -79.430 ;
        RECT -45.310 -79.480 -44.470 -79.430 ;
        RECT -56.610 -82.580 -53.010 -80.975 ;
        RECT -51.650 -81.085 -48.050 -79.480 ;
        RECT -46.690 -82.580 -43.090 -80.975 ;
        RECT -41.730 -81.085 -38.130 -79.480 ;
        RECT -35.390 -79.490 -34.550 -79.430 ;
        RECT -25.470 -79.480 -24.630 -79.430 ;
        RECT -36.770 -82.580 -33.170 -80.975 ;
        RECT -31.810 -81.085 -28.210 -79.480 ;
        RECT -26.850 -82.580 -23.250 -80.975 ;
        RECT -21.890 -81.085 -18.290 -79.480 ;
        RECT -15.550 -79.490 -14.710 -79.430 ;
        RECT -5.630 -79.480 -4.790 -79.430 ;
        RECT -16.930 -82.580 -13.330 -80.975 ;
        RECT -11.970 -81.085 -8.370 -79.480 ;
        RECT -7.010 -82.580 -3.410 -80.975 ;
        RECT -2.050 -81.085 1.550 -79.480 ;
        RECT 4.290 -79.490 5.130 -79.430 ;
        RECT 14.210 -79.480 15.050 -79.430 ;
        RECT 24.130 -79.480 24.970 -79.430 ;
        RECT 2.910 -82.580 6.510 -80.975 ;
        RECT 7.870 -81.085 11.470 -79.480 ;
        RECT 12.830 -82.580 16.430 -80.975 ;
        RECT 17.790 -81.085 21.390 -79.480 ;
        RECT 22.750 -82.580 24.970 -80.975 ;
        RECT -289.815 -84.390 -286.045 -82.630 ;
        RECT -279.895 -84.390 -276.125 -82.630 ;
        RECT -269.975 -84.390 -266.205 -82.630 ;
        RECT -260.055 -84.390 -256.285 -82.630 ;
        RECT -250.135 -84.390 -246.365 -82.630 ;
        RECT -240.215 -84.390 -236.445 -82.630 ;
        RECT -230.295 -84.390 -226.525 -82.630 ;
        RECT -220.375 -84.390 -216.605 -82.630 ;
        RECT -210.455 -84.390 -206.685 -82.630 ;
        RECT -200.535 -84.390 -196.765 -82.630 ;
        RECT -190.615 -84.390 -186.845 -82.630 ;
        RECT -180.695 -84.390 -176.925 -82.630 ;
        RECT -170.775 -84.390 -167.005 -82.630 ;
        RECT -160.855 -84.390 -157.085 -82.630 ;
        RECT -150.935 -84.390 -147.165 -82.630 ;
        RECT -141.015 -84.390 -137.245 -82.630 ;
        RECT -131.095 -84.390 -127.325 -82.630 ;
        RECT -121.175 -84.390 -117.405 -82.630 ;
        RECT -111.255 -84.390 -107.485 -82.630 ;
        RECT -101.335 -84.390 -97.565 -82.630 ;
        RECT -91.415 -84.390 -87.645 -82.630 ;
        RECT -81.495 -84.390 -77.725 -82.630 ;
        RECT -71.575 -84.390 -67.805 -82.630 ;
        RECT -61.655 -84.390 -57.885 -82.630 ;
        RECT -51.735 -84.390 -47.965 -82.630 ;
        RECT -41.815 -84.390 -38.045 -82.630 ;
        RECT -31.895 -84.390 -28.125 -82.630 ;
        RECT -21.975 -84.390 -18.205 -82.630 ;
        RECT -12.055 -84.390 -8.285 -82.630 ;
        RECT -2.135 -84.390 1.635 -82.630 ;
        RECT 7.785 -84.390 11.555 -82.630 ;
        RECT 17.705 -84.390 21.475 -82.630 ;
        RECT -286.615 -174.010 -282.845 -172.250 ;
        RECT -276.695 -174.010 -272.925 -172.250 ;
        RECT -266.775 -174.010 -263.005 -172.250 ;
        RECT -256.855 -174.010 -253.085 -172.250 ;
        RECT -246.935 -174.010 -243.165 -172.250 ;
        RECT -237.015 -174.010 -233.245 -172.250 ;
        RECT -227.095 -174.010 -223.325 -172.250 ;
        RECT -217.175 -174.010 -213.405 -172.250 ;
        RECT -207.255 -174.010 -203.485 -172.250 ;
        RECT -197.335 -174.010 -193.565 -172.250 ;
        RECT -187.415 -174.010 -183.645 -172.250 ;
        RECT -177.495 -174.010 -173.725 -172.250 ;
        RECT -167.575 -174.010 -163.805 -172.250 ;
        RECT -157.655 -174.010 -153.885 -172.250 ;
        RECT -147.735 -174.010 -143.965 -172.250 ;
        RECT -137.815 -174.010 -134.045 -172.250 ;
        RECT -127.895 -174.010 -124.125 -172.250 ;
        RECT -117.975 -174.010 -114.205 -172.250 ;
        RECT -108.055 -174.010 -104.285 -172.250 ;
        RECT -98.135 -174.010 -94.365 -172.250 ;
        RECT -88.215 -174.010 -84.445 -172.250 ;
        RECT -78.295 -174.010 -74.525 -172.250 ;
        RECT -68.375 -174.010 -64.605 -172.250 ;
        RECT -58.455 -174.010 -54.685 -172.250 ;
        RECT -48.535 -174.010 -44.765 -172.250 ;
        RECT -38.615 -174.010 -34.845 -172.250 ;
        RECT -28.695 -174.010 -24.925 -172.250 ;
        RECT -18.775 -174.010 -15.005 -172.250 ;
        RECT -8.855 -174.010 -5.085 -172.250 ;
        RECT 1.065 -174.010 4.835 -172.250 ;
        RECT 10.985 -174.010 14.755 -172.250 ;
        RECT 20.905 -172.485 22.510 -172.250 ;
        RECT 20.905 -172.490 23.020 -172.485 ;
        RECT 20.905 -174.010 23.210 -172.490 ;
        RECT -285.150 -174.060 -284.310 -174.010 ;
        RECT -291.490 -175.665 -287.890 -174.060 ;
        RECT -286.530 -177.160 -282.930 -175.555 ;
        RECT -281.570 -175.665 -277.970 -174.060 ;
        RECT -275.230 -174.070 -274.390 -174.010 ;
        RECT -265.310 -174.060 -264.470 -174.010 ;
        RECT -276.610 -177.160 -273.010 -175.555 ;
        RECT -271.650 -175.665 -268.050 -174.060 ;
        RECT -266.690 -177.160 -263.090 -175.555 ;
        RECT -261.730 -175.665 -258.130 -174.060 ;
        RECT -255.390 -174.070 -254.550 -174.010 ;
        RECT -245.470 -174.060 -244.630 -174.010 ;
        RECT -256.770 -177.160 -253.170 -175.555 ;
        RECT -251.810 -175.665 -248.210 -174.060 ;
        RECT -246.850 -177.160 -243.250 -175.555 ;
        RECT -241.890 -175.665 -238.290 -174.060 ;
        RECT -235.550 -174.070 -234.710 -174.010 ;
        RECT -225.630 -174.060 -224.790 -174.010 ;
        RECT -236.930 -177.160 -233.330 -175.555 ;
        RECT -231.970 -175.665 -228.370 -174.060 ;
        RECT -227.010 -177.160 -223.410 -175.555 ;
        RECT -222.050 -175.665 -218.450 -174.060 ;
        RECT -215.710 -174.070 -214.870 -174.010 ;
        RECT -205.790 -174.060 -204.950 -174.010 ;
        RECT -217.090 -177.160 -213.490 -175.555 ;
        RECT -212.130 -175.665 -208.530 -174.060 ;
        RECT -207.170 -177.160 -203.570 -175.555 ;
        RECT -202.210 -175.665 -198.610 -174.060 ;
        RECT -195.870 -174.070 -195.030 -174.010 ;
        RECT -185.950 -174.060 -185.110 -174.010 ;
        RECT -197.250 -177.160 -193.650 -175.555 ;
        RECT -192.290 -175.665 -188.690 -174.060 ;
        RECT -187.330 -177.160 -183.730 -175.555 ;
        RECT -182.370 -175.665 -178.770 -174.060 ;
        RECT -176.030 -174.070 -175.190 -174.010 ;
        RECT -166.110 -174.060 -165.270 -174.010 ;
        RECT -177.410 -177.160 -173.810 -175.555 ;
        RECT -172.450 -175.665 -168.850 -174.060 ;
        RECT -167.490 -177.160 -163.890 -175.555 ;
        RECT -162.530 -175.665 -158.930 -174.060 ;
        RECT -156.190 -174.070 -155.350 -174.010 ;
        RECT -146.270 -174.060 -145.430 -174.010 ;
        RECT -157.570 -177.160 -153.970 -175.555 ;
        RECT -152.610 -175.665 -149.010 -174.060 ;
        RECT -147.650 -177.160 -144.050 -175.555 ;
        RECT -142.690 -175.665 -139.090 -174.060 ;
        RECT -136.350 -174.070 -135.510 -174.010 ;
        RECT -126.430 -174.060 -125.590 -174.010 ;
        RECT -137.730 -177.160 -134.130 -175.555 ;
        RECT -132.770 -175.665 -129.170 -174.060 ;
        RECT -127.810 -177.160 -124.210 -175.555 ;
        RECT -122.850 -175.665 -119.250 -174.060 ;
        RECT -116.510 -174.070 -115.670 -174.010 ;
        RECT -106.590 -174.060 -105.750 -174.010 ;
        RECT -117.890 -177.160 -114.290 -175.555 ;
        RECT -112.930 -175.665 -109.330 -174.060 ;
        RECT -107.970 -177.160 -104.370 -175.555 ;
        RECT -103.010 -175.665 -99.410 -174.060 ;
        RECT -96.670 -174.070 -95.830 -174.010 ;
        RECT -86.750 -174.060 -85.910 -174.010 ;
        RECT -98.050 -177.160 -94.450 -175.555 ;
        RECT -93.090 -175.665 -89.490 -174.060 ;
        RECT -88.130 -177.160 -84.530 -175.555 ;
        RECT -83.170 -175.665 -79.570 -174.060 ;
        RECT -76.830 -174.070 -75.990 -174.010 ;
        RECT -66.910 -174.060 -66.070 -174.010 ;
        RECT -78.210 -177.160 -74.610 -175.555 ;
        RECT -73.250 -175.665 -69.650 -174.060 ;
        RECT -68.290 -177.160 -64.690 -175.555 ;
        RECT -63.330 -175.665 -59.730 -174.060 ;
        RECT -56.990 -174.070 -56.150 -174.010 ;
        RECT -47.070 -174.060 -46.230 -174.010 ;
        RECT -58.370 -177.160 -54.770 -175.555 ;
        RECT -53.410 -175.665 -49.810 -174.060 ;
        RECT -48.450 -177.160 -44.850 -175.555 ;
        RECT -43.490 -175.665 -39.890 -174.060 ;
        RECT -37.150 -174.070 -36.310 -174.010 ;
        RECT -27.230 -174.060 -26.390 -174.010 ;
        RECT -38.530 -177.160 -34.930 -175.555 ;
        RECT -33.570 -175.665 -29.970 -174.060 ;
        RECT -28.610 -177.160 -25.010 -175.555 ;
        RECT -23.650 -175.665 -20.050 -174.060 ;
        RECT -17.310 -174.070 -16.470 -174.010 ;
        RECT -7.390 -174.060 -6.550 -174.010 ;
        RECT -18.690 -177.160 -15.090 -175.555 ;
        RECT -13.730 -175.665 -10.130 -174.060 ;
        RECT -8.770 -177.160 -5.170 -175.555 ;
        RECT -3.810 -175.665 -0.210 -174.060 ;
        RECT 2.530 -174.070 3.370 -174.010 ;
        RECT 12.450 -174.060 13.290 -174.010 ;
        RECT 22.370 -174.060 23.210 -174.010 ;
        RECT 1.150 -177.160 4.750 -175.555 ;
        RECT 6.110 -175.665 9.710 -174.060 ;
        RECT 11.070 -177.160 14.670 -175.555 ;
        RECT 16.030 -175.665 19.630 -174.060 ;
        RECT 20.990 -177.160 23.210 -175.555 ;
        RECT -291.575 -178.970 -287.805 -177.210 ;
        RECT -281.655 -178.970 -277.885 -177.210 ;
        RECT -271.735 -178.970 -267.965 -177.210 ;
        RECT -261.815 -178.970 -258.045 -177.210 ;
        RECT -251.895 -178.970 -248.125 -177.210 ;
        RECT -241.975 -178.970 -238.205 -177.210 ;
        RECT -232.055 -178.970 -228.285 -177.210 ;
        RECT -222.135 -178.970 -218.365 -177.210 ;
        RECT -212.215 -178.970 -208.445 -177.210 ;
        RECT -202.295 -178.970 -198.525 -177.210 ;
        RECT -192.375 -178.970 -188.605 -177.210 ;
        RECT -182.455 -178.970 -178.685 -177.210 ;
        RECT -172.535 -178.970 -168.765 -177.210 ;
        RECT -162.615 -178.970 -158.845 -177.210 ;
        RECT -152.695 -178.970 -148.925 -177.210 ;
        RECT -142.775 -178.970 -139.005 -177.210 ;
        RECT -132.855 -178.970 -129.085 -177.210 ;
        RECT -122.935 -178.970 -119.165 -177.210 ;
        RECT -113.015 -178.970 -109.245 -177.210 ;
        RECT -103.095 -178.970 -99.325 -177.210 ;
        RECT -93.175 -178.970 -89.405 -177.210 ;
        RECT -83.255 -178.970 -79.485 -177.210 ;
        RECT -73.335 -178.970 -69.565 -177.210 ;
        RECT -63.415 -178.970 -59.645 -177.210 ;
        RECT -53.495 -178.970 -49.725 -177.210 ;
        RECT -43.575 -178.970 -39.805 -177.210 ;
        RECT -33.655 -178.970 -29.885 -177.210 ;
        RECT -23.735 -178.970 -19.965 -177.210 ;
        RECT -13.815 -178.970 -10.045 -177.210 ;
        RECT -3.895 -178.970 -0.125 -177.210 ;
        RECT 6.025 -178.970 9.795 -177.210 ;
        RECT 15.945 -178.970 19.715 -177.210 ;
      LAYER li1 ;
        RECT -281.865 94.990 -281.695 95.140 ;
        RECT -280.925 94.990 -280.755 95.140 ;
        RECT -281.865 94.820 -280.755 94.990 ;
        RECT -281.865 94.615 -281.695 94.820 ;
        RECT -282.625 94.285 -281.695 94.615 ;
        RECT -281.865 93.760 -281.695 94.285 ;
        RECT -281.455 93.655 -281.165 94.820 ;
        RECT -280.925 94.615 -280.755 94.820 ;
        RECT -271.945 94.990 -271.775 95.140 ;
        RECT -271.005 94.990 -270.835 95.140 ;
        RECT -271.945 94.820 -270.835 94.990 ;
        RECT -271.945 94.615 -271.775 94.820 ;
        RECT -280.925 94.285 -279.995 94.615 ;
        RECT -272.705 94.285 -271.775 94.615 ;
        RECT -280.925 93.760 -280.755 94.285 ;
        RECT -271.945 93.760 -271.775 94.285 ;
        RECT -271.535 93.655 -271.245 94.820 ;
        RECT -271.005 94.615 -270.835 94.820 ;
        RECT -262.025 94.990 -261.855 95.140 ;
        RECT -261.085 94.990 -260.915 95.140 ;
        RECT -262.025 94.820 -260.915 94.990 ;
        RECT -262.025 94.615 -261.855 94.820 ;
        RECT -271.005 94.285 -270.075 94.615 ;
        RECT -262.785 94.285 -261.855 94.615 ;
        RECT -271.005 93.760 -270.835 94.285 ;
        RECT -262.025 93.760 -261.855 94.285 ;
        RECT -261.615 93.655 -261.325 94.820 ;
        RECT -261.085 94.615 -260.915 94.820 ;
        RECT -252.105 94.990 -251.935 95.140 ;
        RECT -251.165 94.990 -250.995 95.140 ;
        RECT -252.105 94.820 -250.995 94.990 ;
        RECT -252.105 94.615 -251.935 94.820 ;
        RECT -261.085 94.285 -260.155 94.615 ;
        RECT -252.865 94.285 -251.935 94.615 ;
        RECT -261.085 93.760 -260.915 94.285 ;
        RECT -252.105 93.760 -251.935 94.285 ;
        RECT -251.695 93.655 -251.405 94.820 ;
        RECT -251.165 94.615 -250.995 94.820 ;
        RECT -242.185 94.990 -242.015 95.140 ;
        RECT -241.245 94.990 -241.075 95.140 ;
        RECT -242.185 94.820 -241.075 94.990 ;
        RECT -242.185 94.615 -242.015 94.820 ;
        RECT -251.165 94.285 -250.235 94.615 ;
        RECT -242.945 94.285 -242.015 94.615 ;
        RECT -251.165 93.760 -250.995 94.285 ;
        RECT -242.185 93.760 -242.015 94.285 ;
        RECT -241.775 93.655 -241.485 94.820 ;
        RECT -241.245 94.615 -241.075 94.820 ;
        RECT -232.265 94.990 -232.095 95.140 ;
        RECT -231.325 94.990 -231.155 95.140 ;
        RECT -232.265 94.820 -231.155 94.990 ;
        RECT -232.265 94.615 -232.095 94.820 ;
        RECT -241.245 94.285 -240.315 94.615 ;
        RECT -233.025 94.285 -232.095 94.615 ;
        RECT -241.245 93.760 -241.075 94.285 ;
        RECT -232.265 93.760 -232.095 94.285 ;
        RECT -231.855 93.655 -231.565 94.820 ;
        RECT -231.325 94.615 -231.155 94.820 ;
        RECT -222.345 94.990 -222.175 95.140 ;
        RECT -221.405 94.990 -221.235 95.140 ;
        RECT -222.345 94.820 -221.235 94.990 ;
        RECT -222.345 94.615 -222.175 94.820 ;
        RECT -231.325 94.285 -230.395 94.615 ;
        RECT -223.105 94.285 -222.175 94.615 ;
        RECT -231.325 93.760 -231.155 94.285 ;
        RECT -222.345 93.760 -222.175 94.285 ;
        RECT -221.935 93.655 -221.645 94.820 ;
        RECT -221.405 94.615 -221.235 94.820 ;
        RECT -212.425 94.990 -212.255 95.140 ;
        RECT -211.485 94.990 -211.315 95.140 ;
        RECT -212.425 94.820 -211.315 94.990 ;
        RECT -212.425 94.615 -212.255 94.820 ;
        RECT -221.405 94.285 -220.475 94.615 ;
        RECT -213.185 94.285 -212.255 94.615 ;
        RECT -221.405 93.760 -221.235 94.285 ;
        RECT -212.425 93.760 -212.255 94.285 ;
        RECT -212.015 93.655 -211.725 94.820 ;
        RECT -211.485 94.615 -211.315 94.820 ;
        RECT -202.505 94.990 -202.335 95.140 ;
        RECT -201.565 94.990 -201.395 95.140 ;
        RECT -202.505 94.820 -201.395 94.990 ;
        RECT -202.505 94.615 -202.335 94.820 ;
        RECT -211.485 94.285 -210.555 94.615 ;
        RECT -203.265 94.285 -202.335 94.615 ;
        RECT -211.485 93.760 -211.315 94.285 ;
        RECT -202.505 93.760 -202.335 94.285 ;
        RECT -202.095 93.655 -201.805 94.820 ;
        RECT -201.565 94.615 -201.395 94.820 ;
        RECT -192.585 94.990 -192.415 95.140 ;
        RECT -191.645 94.990 -191.475 95.140 ;
        RECT -192.585 94.820 -191.475 94.990 ;
        RECT -192.585 94.615 -192.415 94.820 ;
        RECT -201.565 94.285 -200.635 94.615 ;
        RECT -193.345 94.285 -192.415 94.615 ;
        RECT -201.565 93.760 -201.395 94.285 ;
        RECT -192.585 93.760 -192.415 94.285 ;
        RECT -192.175 93.655 -191.885 94.820 ;
        RECT -191.645 94.615 -191.475 94.820 ;
        RECT -182.665 94.990 -182.495 95.140 ;
        RECT -181.725 94.990 -181.555 95.140 ;
        RECT -182.665 94.820 -181.555 94.990 ;
        RECT -182.665 94.615 -182.495 94.820 ;
        RECT -191.645 94.285 -190.715 94.615 ;
        RECT -183.425 94.285 -182.495 94.615 ;
        RECT -191.645 93.760 -191.475 94.285 ;
        RECT -182.665 93.760 -182.495 94.285 ;
        RECT -182.255 93.655 -181.965 94.820 ;
        RECT -181.725 94.615 -181.555 94.820 ;
        RECT -172.745 94.990 -172.575 95.140 ;
        RECT -171.805 94.990 -171.635 95.140 ;
        RECT -172.745 94.820 -171.635 94.990 ;
        RECT -172.745 94.615 -172.575 94.820 ;
        RECT -181.725 94.285 -180.795 94.615 ;
        RECT -173.505 94.285 -172.575 94.615 ;
        RECT -181.725 93.760 -181.555 94.285 ;
        RECT -172.745 93.760 -172.575 94.285 ;
        RECT -172.335 93.655 -172.045 94.820 ;
        RECT -171.805 94.615 -171.635 94.820 ;
        RECT -162.825 94.990 -162.655 95.140 ;
        RECT -161.885 94.990 -161.715 95.140 ;
        RECT -162.825 94.820 -161.715 94.990 ;
        RECT -162.825 94.615 -162.655 94.820 ;
        RECT -171.805 94.285 -170.875 94.615 ;
        RECT -163.585 94.285 -162.655 94.615 ;
        RECT -171.805 93.760 -171.635 94.285 ;
        RECT -162.825 93.760 -162.655 94.285 ;
        RECT -162.415 93.655 -162.125 94.820 ;
        RECT -161.885 94.615 -161.715 94.820 ;
        RECT -152.905 94.990 -152.735 95.140 ;
        RECT -151.965 94.990 -151.795 95.140 ;
        RECT -152.905 94.820 -151.795 94.990 ;
        RECT -152.905 94.615 -152.735 94.820 ;
        RECT -161.885 94.285 -160.955 94.615 ;
        RECT -153.665 94.285 -152.735 94.615 ;
        RECT -161.885 93.760 -161.715 94.285 ;
        RECT -152.905 93.760 -152.735 94.285 ;
        RECT -152.495 93.655 -152.205 94.820 ;
        RECT -151.965 94.615 -151.795 94.820 ;
        RECT -142.985 94.990 -142.815 95.140 ;
        RECT -142.045 94.990 -141.875 95.140 ;
        RECT -142.985 94.820 -141.875 94.990 ;
        RECT -142.985 94.615 -142.815 94.820 ;
        RECT -151.965 94.285 -151.035 94.615 ;
        RECT -143.745 94.285 -142.815 94.615 ;
        RECT -151.965 93.760 -151.795 94.285 ;
        RECT -142.985 93.760 -142.815 94.285 ;
        RECT -142.575 93.655 -142.285 94.820 ;
        RECT -142.045 94.615 -141.875 94.820 ;
        RECT -133.065 94.990 -132.895 95.140 ;
        RECT -132.125 94.990 -131.955 95.140 ;
        RECT -133.065 94.820 -131.955 94.990 ;
        RECT -133.065 94.615 -132.895 94.820 ;
        RECT -142.045 94.285 -141.115 94.615 ;
        RECT -133.825 94.285 -132.895 94.615 ;
        RECT -142.045 93.760 -141.875 94.285 ;
        RECT -133.065 93.760 -132.895 94.285 ;
        RECT -132.655 93.655 -132.365 94.820 ;
        RECT -132.125 94.615 -131.955 94.820 ;
        RECT -123.145 94.990 -122.975 95.140 ;
        RECT -122.205 94.990 -122.035 95.140 ;
        RECT -123.145 94.820 -122.035 94.990 ;
        RECT -123.145 94.615 -122.975 94.820 ;
        RECT -132.125 94.285 -131.195 94.615 ;
        RECT -123.905 94.285 -122.975 94.615 ;
        RECT -132.125 93.760 -131.955 94.285 ;
        RECT -123.145 93.760 -122.975 94.285 ;
        RECT -122.735 93.655 -122.445 94.820 ;
        RECT -122.205 94.615 -122.035 94.820 ;
        RECT -113.225 94.990 -113.055 95.140 ;
        RECT -112.285 94.990 -112.115 95.140 ;
        RECT -113.225 94.820 -112.115 94.990 ;
        RECT -113.225 94.615 -113.055 94.820 ;
        RECT -122.205 94.285 -121.275 94.615 ;
        RECT -113.985 94.285 -113.055 94.615 ;
        RECT -122.205 93.760 -122.035 94.285 ;
        RECT -113.225 93.760 -113.055 94.285 ;
        RECT -112.815 93.655 -112.525 94.820 ;
        RECT -112.285 94.615 -112.115 94.820 ;
        RECT -103.305 94.990 -103.135 95.140 ;
        RECT -102.365 94.990 -102.195 95.140 ;
        RECT -103.305 94.820 -102.195 94.990 ;
        RECT -103.305 94.615 -103.135 94.820 ;
        RECT -112.285 94.285 -111.355 94.615 ;
        RECT -104.065 94.285 -103.135 94.615 ;
        RECT -112.285 93.760 -112.115 94.285 ;
        RECT -103.305 93.760 -103.135 94.285 ;
        RECT -102.895 93.655 -102.605 94.820 ;
        RECT -102.365 94.615 -102.195 94.820 ;
        RECT -93.385 94.990 -93.215 95.140 ;
        RECT -92.445 94.990 -92.275 95.140 ;
        RECT -93.385 94.820 -92.275 94.990 ;
        RECT -93.385 94.615 -93.215 94.820 ;
        RECT -102.365 94.285 -101.435 94.615 ;
        RECT -94.145 94.285 -93.215 94.615 ;
        RECT -102.365 93.760 -102.195 94.285 ;
        RECT -93.385 93.760 -93.215 94.285 ;
        RECT -92.975 93.655 -92.685 94.820 ;
        RECT -92.445 94.615 -92.275 94.820 ;
        RECT -83.465 94.990 -83.295 95.140 ;
        RECT -82.525 94.990 -82.355 95.140 ;
        RECT -83.465 94.820 -82.355 94.990 ;
        RECT -83.465 94.615 -83.295 94.820 ;
        RECT -92.445 94.285 -91.515 94.615 ;
        RECT -84.225 94.285 -83.295 94.615 ;
        RECT -92.445 93.760 -92.275 94.285 ;
        RECT -83.465 93.760 -83.295 94.285 ;
        RECT -83.055 93.655 -82.765 94.820 ;
        RECT -82.525 94.615 -82.355 94.820 ;
        RECT -73.545 94.990 -73.375 95.140 ;
        RECT -72.605 94.990 -72.435 95.140 ;
        RECT -73.545 94.820 -72.435 94.990 ;
        RECT -73.545 94.615 -73.375 94.820 ;
        RECT -82.525 94.285 -81.595 94.615 ;
        RECT -74.305 94.285 -73.375 94.615 ;
        RECT -82.525 93.760 -82.355 94.285 ;
        RECT -73.545 93.760 -73.375 94.285 ;
        RECT -73.135 93.655 -72.845 94.820 ;
        RECT -72.605 94.615 -72.435 94.820 ;
        RECT -63.625 94.990 -63.455 95.140 ;
        RECT -62.685 94.990 -62.515 95.140 ;
        RECT -63.625 94.820 -62.515 94.990 ;
        RECT -63.625 94.615 -63.455 94.820 ;
        RECT -72.605 94.285 -71.675 94.615 ;
        RECT -64.385 94.285 -63.455 94.615 ;
        RECT -72.605 93.760 -72.435 94.285 ;
        RECT -63.625 93.760 -63.455 94.285 ;
        RECT -63.215 93.655 -62.925 94.820 ;
        RECT -62.685 94.615 -62.515 94.820 ;
        RECT -53.705 94.990 -53.535 95.140 ;
        RECT -52.765 94.990 -52.595 95.140 ;
        RECT -53.705 94.820 -52.595 94.990 ;
        RECT -53.705 94.615 -53.535 94.820 ;
        RECT -62.685 94.285 -61.755 94.615 ;
        RECT -54.465 94.285 -53.535 94.615 ;
        RECT -62.685 93.760 -62.515 94.285 ;
        RECT -53.705 93.760 -53.535 94.285 ;
        RECT -53.295 93.655 -53.005 94.820 ;
        RECT -52.765 94.615 -52.595 94.820 ;
        RECT -43.785 94.990 -43.615 95.140 ;
        RECT -42.845 94.990 -42.675 95.140 ;
        RECT -43.785 94.820 -42.675 94.990 ;
        RECT -43.785 94.615 -43.615 94.820 ;
        RECT -52.765 94.285 -51.835 94.615 ;
        RECT -44.545 94.285 -43.615 94.615 ;
        RECT -52.765 93.760 -52.595 94.285 ;
        RECT -43.785 93.760 -43.615 94.285 ;
        RECT -43.375 93.655 -43.085 94.820 ;
        RECT -42.845 94.615 -42.675 94.820 ;
        RECT -33.865 94.990 -33.695 95.140 ;
        RECT -32.925 94.990 -32.755 95.140 ;
        RECT -33.865 94.820 -32.755 94.990 ;
        RECT -33.865 94.615 -33.695 94.820 ;
        RECT -42.845 94.285 -41.915 94.615 ;
        RECT -34.625 94.285 -33.695 94.615 ;
        RECT -42.845 93.760 -42.675 94.285 ;
        RECT -33.865 93.760 -33.695 94.285 ;
        RECT -33.455 93.655 -33.165 94.820 ;
        RECT -32.925 94.615 -32.755 94.820 ;
        RECT -23.945 94.990 -23.775 95.140 ;
        RECT -23.005 94.990 -22.835 95.140 ;
        RECT -23.945 94.820 -22.835 94.990 ;
        RECT -23.945 94.615 -23.775 94.820 ;
        RECT -32.925 94.285 -31.995 94.615 ;
        RECT -24.705 94.285 -23.775 94.615 ;
        RECT -32.925 93.760 -32.755 94.285 ;
        RECT -23.945 93.760 -23.775 94.285 ;
        RECT -23.535 93.655 -23.245 94.820 ;
        RECT -23.005 94.615 -22.835 94.820 ;
        RECT -14.025 94.990 -13.855 95.140 ;
        RECT -13.085 94.990 -12.915 95.140 ;
        RECT -14.025 94.820 -12.915 94.990 ;
        RECT -14.025 94.615 -13.855 94.820 ;
        RECT -23.005 94.285 -22.075 94.615 ;
        RECT -14.785 94.285 -13.855 94.615 ;
        RECT -23.005 93.760 -22.835 94.285 ;
        RECT -14.025 93.760 -13.855 94.285 ;
        RECT -13.615 93.655 -13.325 94.820 ;
        RECT -13.085 94.615 -12.915 94.820 ;
        RECT -4.105 94.990 -3.935 95.140 ;
        RECT -3.165 94.990 -2.995 95.140 ;
        RECT -4.105 94.820 -2.995 94.990 ;
        RECT -4.105 94.615 -3.935 94.820 ;
        RECT -13.085 94.285 -12.155 94.615 ;
        RECT -4.865 94.285 -3.935 94.615 ;
        RECT -13.085 93.760 -12.915 94.285 ;
        RECT -4.105 93.760 -3.935 94.285 ;
        RECT -3.695 93.655 -3.405 94.820 ;
        RECT -3.165 94.615 -2.995 94.820 ;
        RECT 5.815 94.990 5.985 95.140 ;
        RECT 6.755 94.990 6.925 95.140 ;
        RECT 5.815 94.820 6.925 94.990 ;
        RECT 5.815 94.615 5.985 94.820 ;
        RECT -3.165 94.285 -2.235 94.615 ;
        RECT 5.055 94.285 5.985 94.615 ;
        RECT -3.165 93.760 -2.995 94.285 ;
        RECT 5.815 93.760 5.985 94.285 ;
        RECT 6.225 93.655 6.515 94.820 ;
        RECT 6.755 94.615 6.925 94.820 ;
        RECT 15.735 94.990 15.905 95.140 ;
        RECT 16.675 94.990 16.845 95.140 ;
        RECT 15.735 94.820 16.845 94.990 ;
        RECT 15.735 94.615 15.905 94.820 ;
        RECT 6.755 94.285 7.685 94.615 ;
        RECT 14.975 94.285 15.905 94.615 ;
        RECT 6.755 93.760 6.925 94.285 ;
        RECT 15.735 93.760 15.905 94.285 ;
        RECT 16.145 93.655 16.435 94.820 ;
        RECT 16.675 94.615 16.845 94.820 ;
        RECT 25.655 94.990 25.825 95.140 ;
        RECT 25.655 94.820 26.440 94.990 ;
        RECT 25.655 94.615 25.825 94.820 ;
        RECT 16.675 94.285 17.605 94.615 ;
        RECT 24.895 94.285 25.825 94.615 ;
        RECT 16.675 93.760 16.845 94.285 ;
        RECT 25.655 93.760 25.825 94.285 ;
        RECT 26.065 93.655 26.355 94.820 ;
        RECT -287.880 93.245 -284.660 93.415 ;
        RECT -277.960 93.245 -274.740 93.415 ;
        RECT -268.040 93.245 -264.820 93.415 ;
        RECT -258.120 93.245 -254.900 93.415 ;
        RECT -248.200 93.245 -244.980 93.415 ;
        RECT -238.280 93.245 -235.060 93.415 ;
        RECT -228.360 93.245 -225.140 93.415 ;
        RECT -218.440 93.245 -215.220 93.415 ;
        RECT -208.520 93.245 -205.300 93.415 ;
        RECT -198.600 93.245 -195.380 93.415 ;
        RECT -188.680 93.245 -185.460 93.415 ;
        RECT -178.760 93.245 -175.540 93.415 ;
        RECT -168.840 93.245 -165.620 93.415 ;
        RECT -158.920 93.245 -155.700 93.415 ;
        RECT -149.000 93.245 -145.780 93.415 ;
        RECT -139.080 93.245 -135.860 93.415 ;
        RECT -129.160 93.245 -125.940 93.415 ;
        RECT -119.240 93.245 -116.020 93.415 ;
        RECT -109.320 93.245 -106.100 93.415 ;
        RECT -99.400 93.245 -96.180 93.415 ;
        RECT -89.480 93.245 -86.260 93.415 ;
        RECT -79.560 93.245 -76.340 93.415 ;
        RECT -69.640 93.245 -66.420 93.415 ;
        RECT -59.720 93.245 -56.500 93.415 ;
        RECT -49.800 93.245 -46.580 93.415 ;
        RECT -39.880 93.245 -36.660 93.415 ;
        RECT -29.960 93.245 -26.740 93.415 ;
        RECT -20.040 93.245 -16.820 93.415 ;
        RECT -10.120 93.245 -6.900 93.415 ;
        RECT -0.200 93.245 3.020 93.415 ;
        RECT 9.720 93.245 12.940 93.415 ;
        RECT 19.640 93.245 22.860 93.415 ;
        RECT -287.795 92.105 -287.535 93.245 ;
        RECT -286.865 92.105 -286.585 93.245 ;
        RECT -286.415 92.080 -286.125 93.245 ;
        RECT -285.955 92.105 -285.675 93.245 ;
        RECT -285.005 92.105 -284.745 93.245 ;
        RECT -277.875 92.105 -277.615 93.245 ;
        RECT -276.945 92.105 -276.665 93.245 ;
        RECT -276.495 92.080 -276.205 93.245 ;
        RECT -276.035 92.105 -275.755 93.245 ;
        RECT -275.085 92.105 -274.825 93.245 ;
        RECT -267.955 92.105 -267.695 93.245 ;
        RECT -267.025 92.105 -266.745 93.245 ;
        RECT -266.575 92.080 -266.285 93.245 ;
        RECT -266.115 92.105 -265.835 93.245 ;
        RECT -265.165 92.105 -264.905 93.245 ;
        RECT -258.035 92.105 -257.775 93.245 ;
        RECT -257.105 92.105 -256.825 93.245 ;
        RECT -256.655 92.080 -256.365 93.245 ;
        RECT -256.195 92.105 -255.915 93.245 ;
        RECT -255.245 92.105 -254.985 93.245 ;
        RECT -248.115 92.105 -247.855 93.245 ;
        RECT -247.185 92.105 -246.905 93.245 ;
        RECT -246.735 92.080 -246.445 93.245 ;
        RECT -246.275 92.105 -245.995 93.245 ;
        RECT -245.325 92.105 -245.065 93.245 ;
        RECT -238.195 92.105 -237.935 93.245 ;
        RECT -237.265 92.105 -236.985 93.245 ;
        RECT -236.815 92.080 -236.525 93.245 ;
        RECT -236.355 92.105 -236.075 93.245 ;
        RECT -235.405 92.105 -235.145 93.245 ;
        RECT -228.275 92.105 -228.015 93.245 ;
        RECT -227.345 92.105 -227.065 93.245 ;
        RECT -226.895 92.080 -226.605 93.245 ;
        RECT -226.435 92.105 -226.155 93.245 ;
        RECT -225.485 92.105 -225.225 93.245 ;
        RECT -218.355 92.105 -218.095 93.245 ;
        RECT -217.425 92.105 -217.145 93.245 ;
        RECT -216.975 92.080 -216.685 93.245 ;
        RECT -216.515 92.105 -216.235 93.245 ;
        RECT -215.565 92.105 -215.305 93.245 ;
        RECT -208.435 92.105 -208.175 93.245 ;
        RECT -207.505 92.105 -207.225 93.245 ;
        RECT -207.055 92.080 -206.765 93.245 ;
        RECT -206.595 92.105 -206.315 93.245 ;
        RECT -205.645 92.105 -205.385 93.245 ;
        RECT -198.515 92.105 -198.255 93.245 ;
        RECT -197.585 92.105 -197.305 93.245 ;
        RECT -197.135 92.080 -196.845 93.245 ;
        RECT -196.675 92.105 -196.395 93.245 ;
        RECT -195.725 92.105 -195.465 93.245 ;
        RECT -188.595 92.105 -188.335 93.245 ;
        RECT -187.665 92.105 -187.385 93.245 ;
        RECT -187.215 92.080 -186.925 93.245 ;
        RECT -186.755 92.105 -186.475 93.245 ;
        RECT -185.805 92.105 -185.545 93.245 ;
        RECT -178.675 92.105 -178.415 93.245 ;
        RECT -177.745 92.105 -177.465 93.245 ;
        RECT -177.295 92.080 -177.005 93.245 ;
        RECT -176.835 92.105 -176.555 93.245 ;
        RECT -175.885 92.105 -175.625 93.245 ;
        RECT -168.755 92.105 -168.495 93.245 ;
        RECT -167.825 92.105 -167.545 93.245 ;
        RECT -167.375 92.080 -167.085 93.245 ;
        RECT -166.915 92.105 -166.635 93.245 ;
        RECT -165.965 92.105 -165.705 93.245 ;
        RECT -158.835 92.105 -158.575 93.245 ;
        RECT -157.905 92.105 -157.625 93.245 ;
        RECT -157.455 92.080 -157.165 93.245 ;
        RECT -156.995 92.105 -156.715 93.245 ;
        RECT -156.045 92.105 -155.785 93.245 ;
        RECT -148.915 92.105 -148.655 93.245 ;
        RECT -147.985 92.105 -147.705 93.245 ;
        RECT -147.535 92.080 -147.245 93.245 ;
        RECT -147.075 92.105 -146.795 93.245 ;
        RECT -146.125 92.105 -145.865 93.245 ;
        RECT -138.995 92.105 -138.735 93.245 ;
        RECT -138.065 92.105 -137.785 93.245 ;
        RECT -137.615 92.080 -137.325 93.245 ;
        RECT -137.155 92.105 -136.875 93.245 ;
        RECT -136.205 92.105 -135.945 93.245 ;
        RECT -129.075 92.105 -128.815 93.245 ;
        RECT -128.145 92.105 -127.865 93.245 ;
        RECT -127.695 92.080 -127.405 93.245 ;
        RECT -127.235 92.105 -126.955 93.245 ;
        RECT -126.285 92.105 -126.025 93.245 ;
        RECT -119.155 92.105 -118.895 93.245 ;
        RECT -118.225 92.105 -117.945 93.245 ;
        RECT -117.775 92.080 -117.485 93.245 ;
        RECT -117.315 92.105 -117.035 93.245 ;
        RECT -116.365 92.105 -116.105 93.245 ;
        RECT -109.235 92.105 -108.975 93.245 ;
        RECT -108.305 92.105 -108.025 93.245 ;
        RECT -107.855 92.080 -107.565 93.245 ;
        RECT -107.395 92.105 -107.115 93.245 ;
        RECT -106.445 92.105 -106.185 93.245 ;
        RECT -99.315 92.105 -99.055 93.245 ;
        RECT -98.385 92.105 -98.105 93.245 ;
        RECT -97.935 92.080 -97.645 93.245 ;
        RECT -97.475 92.105 -97.195 93.245 ;
        RECT -96.525 92.105 -96.265 93.245 ;
        RECT -89.395 92.105 -89.135 93.245 ;
        RECT -88.465 92.105 -88.185 93.245 ;
        RECT -88.015 92.080 -87.725 93.245 ;
        RECT -87.555 92.105 -87.275 93.245 ;
        RECT -86.605 92.105 -86.345 93.245 ;
        RECT -79.475 92.105 -79.215 93.245 ;
        RECT -78.545 92.105 -78.265 93.245 ;
        RECT -78.095 92.080 -77.805 93.245 ;
        RECT -77.635 92.105 -77.355 93.245 ;
        RECT -76.685 92.105 -76.425 93.245 ;
        RECT -69.555 92.105 -69.295 93.245 ;
        RECT -68.625 92.105 -68.345 93.245 ;
        RECT -68.175 92.080 -67.885 93.245 ;
        RECT -67.715 92.105 -67.435 93.245 ;
        RECT -66.765 92.105 -66.505 93.245 ;
        RECT -59.635 92.105 -59.375 93.245 ;
        RECT -58.705 92.105 -58.425 93.245 ;
        RECT -58.255 92.080 -57.965 93.245 ;
        RECT -57.795 92.105 -57.515 93.245 ;
        RECT -56.845 92.105 -56.585 93.245 ;
        RECT -49.715 92.105 -49.455 93.245 ;
        RECT -48.785 92.105 -48.505 93.245 ;
        RECT -48.335 92.080 -48.045 93.245 ;
        RECT -47.875 92.105 -47.595 93.245 ;
        RECT -46.925 92.105 -46.665 93.245 ;
        RECT -39.795 92.105 -39.535 93.245 ;
        RECT -38.865 92.105 -38.585 93.245 ;
        RECT -38.415 92.080 -38.125 93.245 ;
        RECT -37.955 92.105 -37.675 93.245 ;
        RECT -37.005 92.105 -36.745 93.245 ;
        RECT -29.875 92.105 -29.615 93.245 ;
        RECT -28.945 92.105 -28.665 93.245 ;
        RECT -28.495 92.080 -28.205 93.245 ;
        RECT -28.035 92.105 -27.755 93.245 ;
        RECT -27.085 92.105 -26.825 93.245 ;
        RECT -19.955 92.105 -19.695 93.245 ;
        RECT -19.025 92.105 -18.745 93.245 ;
        RECT -18.575 92.080 -18.285 93.245 ;
        RECT -18.115 92.105 -17.835 93.245 ;
        RECT -17.165 92.105 -16.905 93.245 ;
        RECT -10.035 92.105 -9.775 93.245 ;
        RECT -9.105 92.105 -8.825 93.245 ;
        RECT -8.655 92.080 -8.365 93.245 ;
        RECT -8.195 92.105 -7.915 93.245 ;
        RECT -7.245 92.105 -6.985 93.245 ;
        RECT -0.115 92.105 0.145 93.245 ;
        RECT 0.815 92.105 1.095 93.245 ;
        RECT 1.265 92.080 1.555 93.245 ;
        RECT 1.725 92.105 2.005 93.245 ;
        RECT 2.675 92.105 2.935 93.245 ;
        RECT 9.805 92.105 10.065 93.245 ;
        RECT 10.735 92.105 11.015 93.245 ;
        RECT 11.185 92.080 11.475 93.245 ;
        RECT 11.645 92.105 11.925 93.245 ;
        RECT 12.595 92.105 12.855 93.245 ;
        RECT 19.725 92.105 19.985 93.245 ;
        RECT 20.655 92.105 20.935 93.245 ;
        RECT 21.105 92.080 21.395 93.245 ;
        RECT 21.565 92.105 21.845 93.245 ;
        RECT 22.515 92.105 22.775 93.245 ;
        RECT -282.835 90.695 -282.575 91.835 ;
        RECT -281.905 90.695 -281.625 91.835 ;
        RECT -281.455 90.695 -281.165 91.860 ;
        RECT -280.995 90.695 -280.715 91.835 ;
        RECT -280.045 90.695 -279.785 91.835 ;
        RECT -272.915 90.695 -272.655 91.835 ;
        RECT -271.985 90.695 -271.705 91.835 ;
        RECT -271.535 90.695 -271.245 91.860 ;
        RECT -271.075 90.695 -270.795 91.835 ;
        RECT -270.125 90.695 -269.865 91.835 ;
        RECT -262.995 90.695 -262.735 91.835 ;
        RECT -262.065 90.695 -261.785 91.835 ;
        RECT -261.615 90.695 -261.325 91.860 ;
        RECT -261.155 90.695 -260.875 91.835 ;
        RECT -260.205 90.695 -259.945 91.835 ;
        RECT -253.075 90.695 -252.815 91.835 ;
        RECT -252.145 90.695 -251.865 91.835 ;
        RECT -251.695 90.695 -251.405 91.860 ;
        RECT -251.235 90.695 -250.955 91.835 ;
        RECT -250.285 90.695 -250.025 91.835 ;
        RECT -243.155 90.695 -242.895 91.835 ;
        RECT -242.225 90.695 -241.945 91.835 ;
        RECT -241.775 90.695 -241.485 91.860 ;
        RECT -241.315 90.695 -241.035 91.835 ;
        RECT -240.365 90.695 -240.105 91.835 ;
        RECT -233.235 90.695 -232.975 91.835 ;
        RECT -232.305 90.695 -232.025 91.835 ;
        RECT -231.855 90.695 -231.565 91.860 ;
        RECT -231.395 90.695 -231.115 91.835 ;
        RECT -230.445 90.695 -230.185 91.835 ;
        RECT -223.315 90.695 -223.055 91.835 ;
        RECT -222.385 90.695 -222.105 91.835 ;
        RECT -221.935 90.695 -221.645 91.860 ;
        RECT -221.475 90.695 -221.195 91.835 ;
        RECT -220.525 90.695 -220.265 91.835 ;
        RECT -213.395 90.695 -213.135 91.835 ;
        RECT -212.465 90.695 -212.185 91.835 ;
        RECT -212.015 90.695 -211.725 91.860 ;
        RECT -211.555 90.695 -211.275 91.835 ;
        RECT -210.605 90.695 -210.345 91.835 ;
        RECT -203.475 90.695 -203.215 91.835 ;
        RECT -202.545 90.695 -202.265 91.835 ;
        RECT -202.095 90.695 -201.805 91.860 ;
        RECT -201.635 90.695 -201.355 91.835 ;
        RECT -200.685 90.695 -200.425 91.835 ;
        RECT -193.555 90.695 -193.295 91.835 ;
        RECT -192.625 90.695 -192.345 91.835 ;
        RECT -192.175 90.695 -191.885 91.860 ;
        RECT -191.715 90.695 -191.435 91.835 ;
        RECT -190.765 90.695 -190.505 91.835 ;
        RECT -183.635 90.695 -183.375 91.835 ;
        RECT -182.705 90.695 -182.425 91.835 ;
        RECT -182.255 90.695 -181.965 91.860 ;
        RECT -181.795 90.695 -181.515 91.835 ;
        RECT -180.845 90.695 -180.585 91.835 ;
        RECT -173.715 90.695 -173.455 91.835 ;
        RECT -172.785 90.695 -172.505 91.835 ;
        RECT -172.335 90.695 -172.045 91.860 ;
        RECT -171.875 90.695 -171.595 91.835 ;
        RECT -170.925 90.695 -170.665 91.835 ;
        RECT -163.795 90.695 -163.535 91.835 ;
        RECT -162.865 90.695 -162.585 91.835 ;
        RECT -162.415 90.695 -162.125 91.860 ;
        RECT -161.955 90.695 -161.675 91.835 ;
        RECT -161.005 90.695 -160.745 91.835 ;
        RECT -153.875 90.695 -153.615 91.835 ;
        RECT -152.945 90.695 -152.665 91.835 ;
        RECT -152.495 90.695 -152.205 91.860 ;
        RECT -152.035 90.695 -151.755 91.835 ;
        RECT -151.085 90.695 -150.825 91.835 ;
        RECT -143.955 90.695 -143.695 91.835 ;
        RECT -143.025 90.695 -142.745 91.835 ;
        RECT -142.575 90.695 -142.285 91.860 ;
        RECT -142.115 90.695 -141.835 91.835 ;
        RECT -141.165 90.695 -140.905 91.835 ;
        RECT -134.035 90.695 -133.775 91.835 ;
        RECT -133.105 90.695 -132.825 91.835 ;
        RECT -132.655 90.695 -132.365 91.860 ;
        RECT -132.195 90.695 -131.915 91.835 ;
        RECT -131.245 90.695 -130.985 91.835 ;
        RECT -124.115 90.695 -123.855 91.835 ;
        RECT -123.185 90.695 -122.905 91.835 ;
        RECT -122.735 90.695 -122.445 91.860 ;
        RECT -122.275 90.695 -121.995 91.835 ;
        RECT -121.325 90.695 -121.065 91.835 ;
        RECT -114.195 90.695 -113.935 91.835 ;
        RECT -113.265 90.695 -112.985 91.835 ;
        RECT -112.815 90.695 -112.525 91.860 ;
        RECT -112.355 90.695 -112.075 91.835 ;
        RECT -111.405 90.695 -111.145 91.835 ;
        RECT -104.275 90.695 -104.015 91.835 ;
        RECT -103.345 90.695 -103.065 91.835 ;
        RECT -102.895 90.695 -102.605 91.860 ;
        RECT -102.435 90.695 -102.155 91.835 ;
        RECT -101.485 90.695 -101.225 91.835 ;
        RECT -94.355 90.695 -94.095 91.835 ;
        RECT -93.425 90.695 -93.145 91.835 ;
        RECT -92.975 90.695 -92.685 91.860 ;
        RECT -92.515 90.695 -92.235 91.835 ;
        RECT -91.565 90.695 -91.305 91.835 ;
        RECT -84.435 90.695 -84.175 91.835 ;
        RECT -83.505 90.695 -83.225 91.835 ;
        RECT -83.055 90.695 -82.765 91.860 ;
        RECT -82.595 90.695 -82.315 91.835 ;
        RECT -81.645 90.695 -81.385 91.835 ;
        RECT -74.515 90.695 -74.255 91.835 ;
        RECT -73.585 90.695 -73.305 91.835 ;
        RECT -73.135 90.695 -72.845 91.860 ;
        RECT -72.675 90.695 -72.395 91.835 ;
        RECT -71.725 90.695 -71.465 91.835 ;
        RECT -64.595 90.695 -64.335 91.835 ;
        RECT -63.665 90.695 -63.385 91.835 ;
        RECT -63.215 90.695 -62.925 91.860 ;
        RECT -62.755 90.695 -62.475 91.835 ;
        RECT -61.805 90.695 -61.545 91.835 ;
        RECT -54.675 90.695 -54.415 91.835 ;
        RECT -53.745 90.695 -53.465 91.835 ;
        RECT -53.295 90.695 -53.005 91.860 ;
        RECT -52.835 90.695 -52.555 91.835 ;
        RECT -51.885 90.695 -51.625 91.835 ;
        RECT -44.755 90.695 -44.495 91.835 ;
        RECT -43.825 90.695 -43.545 91.835 ;
        RECT -43.375 90.695 -43.085 91.860 ;
        RECT -42.915 90.695 -42.635 91.835 ;
        RECT -41.965 90.695 -41.705 91.835 ;
        RECT -34.835 90.695 -34.575 91.835 ;
        RECT -33.905 90.695 -33.625 91.835 ;
        RECT -33.455 90.695 -33.165 91.860 ;
        RECT -32.995 90.695 -32.715 91.835 ;
        RECT -32.045 90.695 -31.785 91.835 ;
        RECT -24.915 90.695 -24.655 91.835 ;
        RECT -23.985 90.695 -23.705 91.835 ;
        RECT -23.535 90.695 -23.245 91.860 ;
        RECT -23.075 90.695 -22.795 91.835 ;
        RECT -22.125 90.695 -21.865 91.835 ;
        RECT -14.995 90.695 -14.735 91.835 ;
        RECT -14.065 90.695 -13.785 91.835 ;
        RECT -13.615 90.695 -13.325 91.860 ;
        RECT -13.155 90.695 -12.875 91.835 ;
        RECT -12.205 90.695 -11.945 91.835 ;
        RECT -5.075 90.695 -4.815 91.835 ;
        RECT -4.145 90.695 -3.865 91.835 ;
        RECT -3.695 90.695 -3.405 91.860 ;
        RECT -3.235 90.695 -2.955 91.835 ;
        RECT -2.285 90.695 -2.025 91.835 ;
        RECT 4.845 90.695 5.105 91.835 ;
        RECT 5.775 90.695 6.055 91.835 ;
        RECT 6.225 90.695 6.515 91.860 ;
        RECT 6.685 90.695 6.965 91.835 ;
        RECT 7.635 90.695 7.895 91.835 ;
        RECT 14.765 90.695 15.025 91.835 ;
        RECT 15.695 90.695 15.975 91.835 ;
        RECT 16.145 90.695 16.435 91.860 ;
        RECT 16.605 90.695 16.885 91.835 ;
        RECT 17.555 90.695 17.815 91.835 ;
        RECT 24.685 90.695 24.945 91.835 ;
        RECT 25.615 90.695 25.895 91.835 ;
        RECT 26.065 90.695 26.355 91.860 ;
        RECT -282.920 90.525 -279.700 90.695 ;
        RECT -273.000 90.525 -269.780 90.695 ;
        RECT -263.080 90.525 -259.860 90.695 ;
        RECT -253.160 90.525 -249.940 90.695 ;
        RECT -243.240 90.525 -240.020 90.695 ;
        RECT -233.320 90.525 -230.100 90.695 ;
        RECT -223.400 90.525 -220.180 90.695 ;
        RECT -213.480 90.525 -210.260 90.695 ;
        RECT -203.560 90.525 -200.340 90.695 ;
        RECT -193.640 90.525 -190.420 90.695 ;
        RECT -183.720 90.525 -180.500 90.695 ;
        RECT -173.800 90.525 -170.580 90.695 ;
        RECT -163.880 90.525 -160.660 90.695 ;
        RECT -153.960 90.525 -150.740 90.695 ;
        RECT -144.040 90.525 -140.820 90.695 ;
        RECT -134.120 90.525 -130.900 90.695 ;
        RECT -124.200 90.525 -120.980 90.695 ;
        RECT -114.280 90.525 -111.060 90.695 ;
        RECT -104.360 90.525 -101.140 90.695 ;
        RECT -94.440 90.525 -91.220 90.695 ;
        RECT -84.520 90.525 -81.300 90.695 ;
        RECT -74.600 90.525 -71.380 90.695 ;
        RECT -64.680 90.525 -61.460 90.695 ;
        RECT -54.760 90.525 -51.540 90.695 ;
        RECT -44.840 90.525 -41.620 90.695 ;
        RECT -34.920 90.525 -31.700 90.695 ;
        RECT -25.000 90.525 -21.780 90.695 ;
        RECT -15.080 90.525 -11.860 90.695 ;
        RECT -5.160 90.525 -1.940 90.695 ;
        RECT 4.760 90.525 7.980 90.695 ;
        RECT 14.680 90.525 17.900 90.695 ;
        RECT 24.600 90.525 26.440 90.695 ;
        RECT -286.825 90.110 -286.655 90.180 ;
        RECT -285.885 90.110 -285.715 90.180 ;
        RECT -286.825 89.940 -285.715 90.110 ;
        RECT -286.825 89.655 -286.655 89.940 ;
        RECT -287.585 89.325 -286.655 89.655 ;
        RECT -286.825 88.800 -286.655 89.325 ;
        RECT -286.415 88.775 -286.125 89.940 ;
        RECT -285.885 89.655 -285.715 89.940 ;
        RECT -276.905 90.110 -276.735 90.180 ;
        RECT -275.965 90.110 -275.795 90.180 ;
        RECT -276.905 89.940 -275.795 90.110 ;
        RECT -276.905 89.655 -276.735 89.940 ;
        RECT -285.885 89.325 -284.955 89.655 ;
        RECT -277.665 89.325 -276.735 89.655 ;
        RECT -285.885 88.800 -285.715 89.325 ;
        RECT -276.905 88.800 -276.735 89.325 ;
        RECT -276.495 88.775 -276.205 89.940 ;
        RECT -275.965 89.655 -275.795 89.940 ;
        RECT -266.985 90.110 -266.815 90.180 ;
        RECT -266.045 90.110 -265.875 90.180 ;
        RECT -266.985 89.940 -265.875 90.110 ;
        RECT -266.985 89.655 -266.815 89.940 ;
        RECT -275.965 89.325 -275.035 89.655 ;
        RECT -267.745 89.325 -266.815 89.655 ;
        RECT -275.965 88.800 -275.795 89.325 ;
        RECT -266.985 88.800 -266.815 89.325 ;
        RECT -266.575 88.775 -266.285 89.940 ;
        RECT -266.045 89.655 -265.875 89.940 ;
        RECT -257.065 90.110 -256.895 90.180 ;
        RECT -256.125 90.110 -255.955 90.180 ;
        RECT -257.065 89.940 -255.955 90.110 ;
        RECT -257.065 89.655 -256.895 89.940 ;
        RECT -266.045 89.325 -265.115 89.655 ;
        RECT -257.825 89.325 -256.895 89.655 ;
        RECT -266.045 88.800 -265.875 89.325 ;
        RECT -257.065 88.800 -256.895 89.325 ;
        RECT -256.655 88.775 -256.365 89.940 ;
        RECT -256.125 89.655 -255.955 89.940 ;
        RECT -247.145 90.110 -246.975 90.180 ;
        RECT -246.205 90.110 -246.035 90.180 ;
        RECT -247.145 89.940 -246.035 90.110 ;
        RECT -247.145 89.655 -246.975 89.940 ;
        RECT -256.125 89.325 -255.195 89.655 ;
        RECT -247.905 89.325 -246.975 89.655 ;
        RECT -256.125 88.800 -255.955 89.325 ;
        RECT -247.145 88.800 -246.975 89.325 ;
        RECT -246.735 88.775 -246.445 89.940 ;
        RECT -246.205 89.655 -246.035 89.940 ;
        RECT -237.225 90.110 -237.055 90.180 ;
        RECT -236.285 90.110 -236.115 90.180 ;
        RECT -237.225 89.940 -236.115 90.110 ;
        RECT -237.225 89.655 -237.055 89.940 ;
        RECT -246.205 89.325 -245.275 89.655 ;
        RECT -237.985 89.325 -237.055 89.655 ;
        RECT -246.205 88.800 -246.035 89.325 ;
        RECT -237.225 88.800 -237.055 89.325 ;
        RECT -236.815 88.775 -236.525 89.940 ;
        RECT -236.285 89.655 -236.115 89.940 ;
        RECT -227.305 90.110 -227.135 90.180 ;
        RECT -226.365 90.110 -226.195 90.180 ;
        RECT -227.305 89.940 -226.195 90.110 ;
        RECT -227.305 89.655 -227.135 89.940 ;
        RECT -236.285 89.325 -235.355 89.655 ;
        RECT -228.065 89.325 -227.135 89.655 ;
        RECT -236.285 88.800 -236.115 89.325 ;
        RECT -227.305 88.800 -227.135 89.325 ;
        RECT -226.895 88.775 -226.605 89.940 ;
        RECT -226.365 89.655 -226.195 89.940 ;
        RECT -217.385 90.110 -217.215 90.180 ;
        RECT -216.445 90.110 -216.275 90.180 ;
        RECT -217.385 89.940 -216.275 90.110 ;
        RECT -217.385 89.655 -217.215 89.940 ;
        RECT -226.365 89.325 -225.435 89.655 ;
        RECT -218.145 89.325 -217.215 89.655 ;
        RECT -226.365 88.800 -226.195 89.325 ;
        RECT -217.385 88.800 -217.215 89.325 ;
        RECT -216.975 88.775 -216.685 89.940 ;
        RECT -216.445 89.655 -216.275 89.940 ;
        RECT -207.465 90.110 -207.295 90.180 ;
        RECT -206.525 90.110 -206.355 90.180 ;
        RECT -207.465 89.940 -206.355 90.110 ;
        RECT -207.465 89.655 -207.295 89.940 ;
        RECT -216.445 89.325 -215.515 89.655 ;
        RECT -208.225 89.325 -207.295 89.655 ;
        RECT -216.445 88.800 -216.275 89.325 ;
        RECT -207.465 88.800 -207.295 89.325 ;
        RECT -207.055 88.775 -206.765 89.940 ;
        RECT -206.525 89.655 -206.355 89.940 ;
        RECT -197.545 90.110 -197.375 90.180 ;
        RECT -196.605 90.110 -196.435 90.180 ;
        RECT -197.545 89.940 -196.435 90.110 ;
        RECT -197.545 89.655 -197.375 89.940 ;
        RECT -206.525 89.325 -205.595 89.655 ;
        RECT -198.305 89.325 -197.375 89.655 ;
        RECT -206.525 88.800 -206.355 89.325 ;
        RECT -197.545 88.800 -197.375 89.325 ;
        RECT -197.135 88.775 -196.845 89.940 ;
        RECT -196.605 89.655 -196.435 89.940 ;
        RECT -187.625 90.110 -187.455 90.180 ;
        RECT -186.685 90.110 -186.515 90.180 ;
        RECT -187.625 89.940 -186.515 90.110 ;
        RECT -187.625 89.655 -187.455 89.940 ;
        RECT -196.605 89.325 -195.675 89.655 ;
        RECT -188.385 89.325 -187.455 89.655 ;
        RECT -196.605 88.800 -196.435 89.325 ;
        RECT -187.625 88.800 -187.455 89.325 ;
        RECT -187.215 88.775 -186.925 89.940 ;
        RECT -186.685 89.655 -186.515 89.940 ;
        RECT -177.705 90.110 -177.535 90.180 ;
        RECT -176.765 90.110 -176.595 90.180 ;
        RECT -177.705 89.940 -176.595 90.110 ;
        RECT -177.705 89.655 -177.535 89.940 ;
        RECT -186.685 89.325 -185.755 89.655 ;
        RECT -178.465 89.325 -177.535 89.655 ;
        RECT -186.685 88.800 -186.515 89.325 ;
        RECT -177.705 88.800 -177.535 89.325 ;
        RECT -177.295 88.775 -177.005 89.940 ;
        RECT -176.765 89.655 -176.595 89.940 ;
        RECT -167.785 90.110 -167.615 90.180 ;
        RECT -166.845 90.110 -166.675 90.180 ;
        RECT -167.785 89.940 -166.675 90.110 ;
        RECT -167.785 89.655 -167.615 89.940 ;
        RECT -176.765 89.325 -175.835 89.655 ;
        RECT -168.545 89.325 -167.615 89.655 ;
        RECT -176.765 88.800 -176.595 89.325 ;
        RECT -167.785 88.800 -167.615 89.325 ;
        RECT -167.375 88.775 -167.085 89.940 ;
        RECT -166.845 89.655 -166.675 89.940 ;
        RECT -157.865 90.110 -157.695 90.180 ;
        RECT -156.925 90.110 -156.755 90.180 ;
        RECT -157.865 89.940 -156.755 90.110 ;
        RECT -157.865 89.655 -157.695 89.940 ;
        RECT -166.845 89.325 -165.915 89.655 ;
        RECT -158.625 89.325 -157.695 89.655 ;
        RECT -166.845 88.800 -166.675 89.325 ;
        RECT -157.865 88.800 -157.695 89.325 ;
        RECT -157.455 88.775 -157.165 89.940 ;
        RECT -156.925 89.655 -156.755 89.940 ;
        RECT -147.945 90.110 -147.775 90.180 ;
        RECT -147.005 90.110 -146.835 90.180 ;
        RECT -147.945 89.940 -146.835 90.110 ;
        RECT -147.945 89.655 -147.775 89.940 ;
        RECT -156.925 89.325 -155.995 89.655 ;
        RECT -148.705 89.325 -147.775 89.655 ;
        RECT -156.925 88.800 -156.755 89.325 ;
        RECT -147.945 88.800 -147.775 89.325 ;
        RECT -147.535 88.775 -147.245 89.940 ;
        RECT -147.005 89.655 -146.835 89.940 ;
        RECT -138.025 90.110 -137.855 90.180 ;
        RECT -137.085 90.110 -136.915 90.180 ;
        RECT -138.025 89.940 -136.915 90.110 ;
        RECT -138.025 89.655 -137.855 89.940 ;
        RECT -147.005 89.325 -146.075 89.655 ;
        RECT -138.785 89.325 -137.855 89.655 ;
        RECT -147.005 88.800 -146.835 89.325 ;
        RECT -138.025 88.800 -137.855 89.325 ;
        RECT -137.615 88.775 -137.325 89.940 ;
        RECT -137.085 89.655 -136.915 89.940 ;
        RECT -128.105 90.110 -127.935 90.180 ;
        RECT -127.165 90.110 -126.995 90.180 ;
        RECT -128.105 89.940 -126.995 90.110 ;
        RECT -128.105 89.655 -127.935 89.940 ;
        RECT -137.085 89.325 -136.155 89.655 ;
        RECT -128.865 89.325 -127.935 89.655 ;
        RECT -137.085 88.800 -136.915 89.325 ;
        RECT -128.105 88.800 -127.935 89.325 ;
        RECT -127.695 88.775 -127.405 89.940 ;
        RECT -127.165 89.655 -126.995 89.940 ;
        RECT -118.185 90.110 -118.015 90.180 ;
        RECT -117.245 90.110 -117.075 90.180 ;
        RECT -118.185 89.940 -117.075 90.110 ;
        RECT -118.185 89.655 -118.015 89.940 ;
        RECT -127.165 89.325 -126.235 89.655 ;
        RECT -118.945 89.325 -118.015 89.655 ;
        RECT -127.165 88.800 -126.995 89.325 ;
        RECT -118.185 88.800 -118.015 89.325 ;
        RECT -117.775 88.775 -117.485 89.940 ;
        RECT -117.245 89.655 -117.075 89.940 ;
        RECT -108.265 90.110 -108.095 90.180 ;
        RECT -107.325 90.110 -107.155 90.180 ;
        RECT -108.265 89.940 -107.155 90.110 ;
        RECT -108.265 89.655 -108.095 89.940 ;
        RECT -117.245 89.325 -116.315 89.655 ;
        RECT -109.025 89.325 -108.095 89.655 ;
        RECT -117.245 88.800 -117.075 89.325 ;
        RECT -108.265 88.800 -108.095 89.325 ;
        RECT -107.855 88.775 -107.565 89.940 ;
        RECT -107.325 89.655 -107.155 89.940 ;
        RECT -98.345 90.110 -98.175 90.180 ;
        RECT -97.405 90.110 -97.235 90.180 ;
        RECT -98.345 89.940 -97.235 90.110 ;
        RECT -98.345 89.655 -98.175 89.940 ;
        RECT -107.325 89.325 -106.395 89.655 ;
        RECT -99.105 89.325 -98.175 89.655 ;
        RECT -107.325 88.800 -107.155 89.325 ;
        RECT -98.345 88.800 -98.175 89.325 ;
        RECT -97.935 88.775 -97.645 89.940 ;
        RECT -97.405 89.655 -97.235 89.940 ;
        RECT -88.425 90.110 -88.255 90.180 ;
        RECT -87.485 90.110 -87.315 90.180 ;
        RECT -88.425 89.940 -87.315 90.110 ;
        RECT -88.425 89.655 -88.255 89.940 ;
        RECT -97.405 89.325 -96.475 89.655 ;
        RECT -89.185 89.325 -88.255 89.655 ;
        RECT -97.405 88.800 -97.235 89.325 ;
        RECT -88.425 88.800 -88.255 89.325 ;
        RECT -88.015 88.775 -87.725 89.940 ;
        RECT -87.485 89.655 -87.315 89.940 ;
        RECT -78.505 90.110 -78.335 90.180 ;
        RECT -77.565 90.110 -77.395 90.180 ;
        RECT -78.505 89.940 -77.395 90.110 ;
        RECT -78.505 89.655 -78.335 89.940 ;
        RECT -87.485 89.325 -86.555 89.655 ;
        RECT -79.265 89.325 -78.335 89.655 ;
        RECT -87.485 88.800 -87.315 89.325 ;
        RECT -78.505 88.800 -78.335 89.325 ;
        RECT -78.095 88.775 -77.805 89.940 ;
        RECT -77.565 89.655 -77.395 89.940 ;
        RECT -68.585 90.110 -68.415 90.180 ;
        RECT -67.645 90.110 -67.475 90.180 ;
        RECT -68.585 89.940 -67.475 90.110 ;
        RECT -68.585 89.655 -68.415 89.940 ;
        RECT -77.565 89.325 -76.635 89.655 ;
        RECT -69.345 89.325 -68.415 89.655 ;
        RECT -77.565 88.800 -77.395 89.325 ;
        RECT -68.585 88.800 -68.415 89.325 ;
        RECT -68.175 88.775 -67.885 89.940 ;
        RECT -67.645 89.655 -67.475 89.940 ;
        RECT -58.665 90.110 -58.495 90.180 ;
        RECT -57.725 90.110 -57.555 90.180 ;
        RECT -58.665 89.940 -57.555 90.110 ;
        RECT -58.665 89.655 -58.495 89.940 ;
        RECT -67.645 89.325 -66.715 89.655 ;
        RECT -59.425 89.325 -58.495 89.655 ;
        RECT -67.645 88.800 -67.475 89.325 ;
        RECT -58.665 88.800 -58.495 89.325 ;
        RECT -58.255 88.775 -57.965 89.940 ;
        RECT -57.725 89.655 -57.555 89.940 ;
        RECT -48.745 90.110 -48.575 90.180 ;
        RECT -47.805 90.110 -47.635 90.180 ;
        RECT -48.745 89.940 -47.635 90.110 ;
        RECT -48.745 89.655 -48.575 89.940 ;
        RECT -57.725 89.325 -56.795 89.655 ;
        RECT -49.505 89.325 -48.575 89.655 ;
        RECT -57.725 88.800 -57.555 89.325 ;
        RECT -48.745 88.800 -48.575 89.325 ;
        RECT -48.335 88.775 -48.045 89.940 ;
        RECT -47.805 89.655 -47.635 89.940 ;
        RECT -38.825 90.110 -38.655 90.180 ;
        RECT -37.885 90.110 -37.715 90.180 ;
        RECT -38.825 89.940 -37.715 90.110 ;
        RECT -38.825 89.655 -38.655 89.940 ;
        RECT -47.805 89.325 -46.875 89.655 ;
        RECT -39.585 89.325 -38.655 89.655 ;
        RECT -47.805 88.800 -47.635 89.325 ;
        RECT -38.825 88.800 -38.655 89.325 ;
        RECT -38.415 88.775 -38.125 89.940 ;
        RECT -37.885 89.655 -37.715 89.940 ;
        RECT -28.905 90.110 -28.735 90.180 ;
        RECT -27.965 90.110 -27.795 90.180 ;
        RECT -28.905 89.940 -27.795 90.110 ;
        RECT -28.905 89.655 -28.735 89.940 ;
        RECT -37.885 89.325 -36.955 89.655 ;
        RECT -29.665 89.325 -28.735 89.655 ;
        RECT -37.885 88.800 -37.715 89.325 ;
        RECT -28.905 88.800 -28.735 89.325 ;
        RECT -28.495 88.775 -28.205 89.940 ;
        RECT -27.965 89.655 -27.795 89.940 ;
        RECT -18.985 90.110 -18.815 90.180 ;
        RECT -18.045 90.110 -17.875 90.180 ;
        RECT -18.985 89.940 -17.875 90.110 ;
        RECT -18.985 89.655 -18.815 89.940 ;
        RECT -27.965 89.325 -27.035 89.655 ;
        RECT -19.745 89.325 -18.815 89.655 ;
        RECT -27.965 88.800 -27.795 89.325 ;
        RECT -18.985 88.800 -18.815 89.325 ;
        RECT -18.575 88.775 -18.285 89.940 ;
        RECT -18.045 89.655 -17.875 89.940 ;
        RECT -9.065 90.110 -8.895 90.180 ;
        RECT -8.125 90.110 -7.955 90.180 ;
        RECT -9.065 89.940 -7.955 90.110 ;
        RECT -9.065 89.655 -8.895 89.940 ;
        RECT -18.045 89.325 -17.115 89.655 ;
        RECT -9.825 89.325 -8.895 89.655 ;
        RECT -18.045 88.800 -17.875 89.325 ;
        RECT -9.065 88.800 -8.895 89.325 ;
        RECT -8.655 88.775 -8.365 89.940 ;
        RECT -8.125 89.655 -7.955 89.940 ;
        RECT 0.855 90.110 1.025 90.180 ;
        RECT 1.795 90.110 1.965 90.180 ;
        RECT 0.855 89.940 1.965 90.110 ;
        RECT 0.855 89.655 1.025 89.940 ;
        RECT -8.125 89.325 -7.195 89.655 ;
        RECT 0.095 89.325 1.025 89.655 ;
        RECT -8.125 88.800 -7.955 89.325 ;
        RECT 0.855 88.800 1.025 89.325 ;
        RECT 1.265 88.775 1.555 89.940 ;
        RECT 1.795 89.655 1.965 89.940 ;
        RECT 10.775 90.110 10.945 90.180 ;
        RECT 11.715 90.110 11.885 90.180 ;
        RECT 10.775 89.940 11.885 90.110 ;
        RECT 10.775 89.655 10.945 89.940 ;
        RECT 1.795 89.325 2.725 89.655 ;
        RECT 10.015 89.325 10.945 89.655 ;
        RECT 1.795 88.800 1.965 89.325 ;
        RECT 10.775 88.800 10.945 89.325 ;
        RECT 11.185 88.775 11.475 89.940 ;
        RECT 11.715 89.655 11.885 89.940 ;
        RECT 20.695 90.110 20.865 90.180 ;
        RECT 21.635 90.110 21.805 90.180 ;
        RECT 20.695 89.940 21.805 90.110 ;
        RECT 20.695 89.655 20.865 89.940 ;
        RECT 11.715 89.325 12.645 89.655 ;
        RECT 19.935 89.325 20.865 89.655 ;
        RECT 11.715 88.800 11.885 89.325 ;
        RECT 20.695 88.800 20.865 89.325 ;
        RECT 21.105 88.775 21.395 89.940 ;
        RECT 21.635 89.655 21.805 89.940 ;
        RECT 21.635 89.325 22.565 89.655 ;
        RECT 21.635 88.800 21.805 89.325 ;
        RECT -283.885 10.940 -283.715 11.090 ;
        RECT -282.945 10.940 -282.775 11.090 ;
        RECT -283.885 10.770 -282.775 10.940 ;
        RECT -283.885 10.565 -283.715 10.770 ;
        RECT -284.645 10.235 -283.715 10.565 ;
        RECT -283.885 9.710 -283.715 10.235 ;
        RECT -283.475 9.605 -283.185 10.770 ;
        RECT -282.945 10.565 -282.775 10.770 ;
        RECT -273.965 10.940 -273.795 11.090 ;
        RECT -273.025 10.940 -272.855 11.090 ;
        RECT -273.965 10.770 -272.855 10.940 ;
        RECT -273.965 10.565 -273.795 10.770 ;
        RECT -282.945 10.235 -282.015 10.565 ;
        RECT -274.725 10.235 -273.795 10.565 ;
        RECT -282.945 9.710 -282.775 10.235 ;
        RECT -273.965 9.710 -273.795 10.235 ;
        RECT -273.555 9.605 -273.265 10.770 ;
        RECT -273.025 10.565 -272.855 10.770 ;
        RECT -264.045 10.940 -263.875 11.090 ;
        RECT -263.105 10.940 -262.935 11.090 ;
        RECT -264.045 10.770 -262.935 10.940 ;
        RECT -264.045 10.565 -263.875 10.770 ;
        RECT -273.025 10.235 -272.095 10.565 ;
        RECT -264.805 10.235 -263.875 10.565 ;
        RECT -273.025 9.710 -272.855 10.235 ;
        RECT -264.045 9.710 -263.875 10.235 ;
        RECT -263.635 9.605 -263.345 10.770 ;
        RECT -263.105 10.565 -262.935 10.770 ;
        RECT -254.125 10.940 -253.955 11.090 ;
        RECT -253.185 10.940 -253.015 11.090 ;
        RECT -254.125 10.770 -253.015 10.940 ;
        RECT -254.125 10.565 -253.955 10.770 ;
        RECT -263.105 10.235 -262.175 10.565 ;
        RECT -254.885 10.235 -253.955 10.565 ;
        RECT -263.105 9.710 -262.935 10.235 ;
        RECT -254.125 9.710 -253.955 10.235 ;
        RECT -253.715 9.605 -253.425 10.770 ;
        RECT -253.185 10.565 -253.015 10.770 ;
        RECT -244.205 10.940 -244.035 11.090 ;
        RECT -243.265 10.940 -243.095 11.090 ;
        RECT -244.205 10.770 -243.095 10.940 ;
        RECT -244.205 10.565 -244.035 10.770 ;
        RECT -253.185 10.235 -252.255 10.565 ;
        RECT -244.965 10.235 -244.035 10.565 ;
        RECT -253.185 9.710 -253.015 10.235 ;
        RECT -244.205 9.710 -244.035 10.235 ;
        RECT -243.795 9.605 -243.505 10.770 ;
        RECT -243.265 10.565 -243.095 10.770 ;
        RECT -234.285 10.940 -234.115 11.090 ;
        RECT -233.345 10.940 -233.175 11.090 ;
        RECT -234.285 10.770 -233.175 10.940 ;
        RECT -234.285 10.565 -234.115 10.770 ;
        RECT -243.265 10.235 -242.335 10.565 ;
        RECT -235.045 10.235 -234.115 10.565 ;
        RECT -243.265 9.710 -243.095 10.235 ;
        RECT -234.285 9.710 -234.115 10.235 ;
        RECT -233.875 9.605 -233.585 10.770 ;
        RECT -233.345 10.565 -233.175 10.770 ;
        RECT -224.365 10.940 -224.195 11.090 ;
        RECT -223.425 10.940 -223.255 11.090 ;
        RECT -224.365 10.770 -223.255 10.940 ;
        RECT -224.365 10.565 -224.195 10.770 ;
        RECT -233.345 10.235 -232.415 10.565 ;
        RECT -225.125 10.235 -224.195 10.565 ;
        RECT -233.345 9.710 -233.175 10.235 ;
        RECT -224.365 9.710 -224.195 10.235 ;
        RECT -223.955 9.605 -223.665 10.770 ;
        RECT -223.425 10.565 -223.255 10.770 ;
        RECT -214.445 10.940 -214.275 11.090 ;
        RECT -213.505 10.940 -213.335 11.090 ;
        RECT -214.445 10.770 -213.335 10.940 ;
        RECT -214.445 10.565 -214.275 10.770 ;
        RECT -223.425 10.235 -222.495 10.565 ;
        RECT -215.205 10.235 -214.275 10.565 ;
        RECT -223.425 9.710 -223.255 10.235 ;
        RECT -214.445 9.710 -214.275 10.235 ;
        RECT -214.035 9.605 -213.745 10.770 ;
        RECT -213.505 10.565 -213.335 10.770 ;
        RECT -204.525 10.940 -204.355 11.090 ;
        RECT -203.585 10.940 -203.415 11.090 ;
        RECT -204.525 10.770 -203.415 10.940 ;
        RECT -204.525 10.565 -204.355 10.770 ;
        RECT -213.505 10.235 -212.575 10.565 ;
        RECT -205.285 10.235 -204.355 10.565 ;
        RECT -213.505 9.710 -213.335 10.235 ;
        RECT -204.525 9.710 -204.355 10.235 ;
        RECT -204.115 9.605 -203.825 10.770 ;
        RECT -203.585 10.565 -203.415 10.770 ;
        RECT -194.605 10.940 -194.435 11.090 ;
        RECT -193.665 10.940 -193.495 11.090 ;
        RECT -194.605 10.770 -193.495 10.940 ;
        RECT -194.605 10.565 -194.435 10.770 ;
        RECT -203.585 10.235 -202.655 10.565 ;
        RECT -195.365 10.235 -194.435 10.565 ;
        RECT -203.585 9.710 -203.415 10.235 ;
        RECT -194.605 9.710 -194.435 10.235 ;
        RECT -194.195 9.605 -193.905 10.770 ;
        RECT -193.665 10.565 -193.495 10.770 ;
        RECT -184.685 10.940 -184.515 11.090 ;
        RECT -183.745 10.940 -183.575 11.090 ;
        RECT -184.685 10.770 -183.575 10.940 ;
        RECT -184.685 10.565 -184.515 10.770 ;
        RECT -193.665 10.235 -192.735 10.565 ;
        RECT -185.445 10.235 -184.515 10.565 ;
        RECT -193.665 9.710 -193.495 10.235 ;
        RECT -184.685 9.710 -184.515 10.235 ;
        RECT -184.275 9.605 -183.985 10.770 ;
        RECT -183.745 10.565 -183.575 10.770 ;
        RECT -174.765 10.940 -174.595 11.090 ;
        RECT -173.825 10.940 -173.655 11.090 ;
        RECT -174.765 10.770 -173.655 10.940 ;
        RECT -174.765 10.565 -174.595 10.770 ;
        RECT -183.745 10.235 -182.815 10.565 ;
        RECT -175.525 10.235 -174.595 10.565 ;
        RECT -183.745 9.710 -183.575 10.235 ;
        RECT -174.765 9.710 -174.595 10.235 ;
        RECT -174.355 9.605 -174.065 10.770 ;
        RECT -173.825 10.565 -173.655 10.770 ;
        RECT -164.845 10.940 -164.675 11.090 ;
        RECT -163.905 10.940 -163.735 11.090 ;
        RECT -164.845 10.770 -163.735 10.940 ;
        RECT -164.845 10.565 -164.675 10.770 ;
        RECT -173.825 10.235 -172.895 10.565 ;
        RECT -165.605 10.235 -164.675 10.565 ;
        RECT -173.825 9.710 -173.655 10.235 ;
        RECT -164.845 9.710 -164.675 10.235 ;
        RECT -164.435 9.605 -164.145 10.770 ;
        RECT -163.905 10.565 -163.735 10.770 ;
        RECT -154.925 10.940 -154.755 11.090 ;
        RECT -153.985 10.940 -153.815 11.090 ;
        RECT -154.925 10.770 -153.815 10.940 ;
        RECT -154.925 10.565 -154.755 10.770 ;
        RECT -163.905 10.235 -162.975 10.565 ;
        RECT -155.685 10.235 -154.755 10.565 ;
        RECT -163.905 9.710 -163.735 10.235 ;
        RECT -154.925 9.710 -154.755 10.235 ;
        RECT -154.515 9.605 -154.225 10.770 ;
        RECT -153.985 10.565 -153.815 10.770 ;
        RECT -145.005 10.940 -144.835 11.090 ;
        RECT -144.065 10.940 -143.895 11.090 ;
        RECT -145.005 10.770 -143.895 10.940 ;
        RECT -145.005 10.565 -144.835 10.770 ;
        RECT -153.985 10.235 -153.055 10.565 ;
        RECT -145.765 10.235 -144.835 10.565 ;
        RECT -153.985 9.710 -153.815 10.235 ;
        RECT -145.005 9.710 -144.835 10.235 ;
        RECT -144.595 9.605 -144.305 10.770 ;
        RECT -144.065 10.565 -143.895 10.770 ;
        RECT -135.085 10.940 -134.915 11.090 ;
        RECT -134.145 10.940 -133.975 11.090 ;
        RECT -135.085 10.770 -133.975 10.940 ;
        RECT -135.085 10.565 -134.915 10.770 ;
        RECT -144.065 10.235 -143.135 10.565 ;
        RECT -135.845 10.235 -134.915 10.565 ;
        RECT -144.065 9.710 -143.895 10.235 ;
        RECT -135.085 9.710 -134.915 10.235 ;
        RECT -134.675 9.605 -134.385 10.770 ;
        RECT -134.145 10.565 -133.975 10.770 ;
        RECT -125.165 10.940 -124.995 11.090 ;
        RECT -124.225 10.940 -124.055 11.090 ;
        RECT -125.165 10.770 -124.055 10.940 ;
        RECT -125.165 10.565 -124.995 10.770 ;
        RECT -134.145 10.235 -133.215 10.565 ;
        RECT -125.925 10.235 -124.995 10.565 ;
        RECT -134.145 9.710 -133.975 10.235 ;
        RECT -125.165 9.710 -124.995 10.235 ;
        RECT -124.755 9.605 -124.465 10.770 ;
        RECT -124.225 10.565 -124.055 10.770 ;
        RECT -115.245 10.940 -115.075 11.090 ;
        RECT -114.305 10.940 -114.135 11.090 ;
        RECT -115.245 10.770 -114.135 10.940 ;
        RECT -115.245 10.565 -115.075 10.770 ;
        RECT -124.225 10.235 -123.295 10.565 ;
        RECT -116.005 10.235 -115.075 10.565 ;
        RECT -124.225 9.710 -124.055 10.235 ;
        RECT -115.245 9.710 -115.075 10.235 ;
        RECT -114.835 9.605 -114.545 10.770 ;
        RECT -114.305 10.565 -114.135 10.770 ;
        RECT -105.325 10.940 -105.155 11.090 ;
        RECT -104.385 10.940 -104.215 11.090 ;
        RECT -105.325 10.770 -104.215 10.940 ;
        RECT -105.325 10.565 -105.155 10.770 ;
        RECT -114.305 10.235 -113.375 10.565 ;
        RECT -106.085 10.235 -105.155 10.565 ;
        RECT -114.305 9.710 -114.135 10.235 ;
        RECT -105.325 9.710 -105.155 10.235 ;
        RECT -104.915 9.605 -104.625 10.770 ;
        RECT -104.385 10.565 -104.215 10.770 ;
        RECT -95.405 10.940 -95.235 11.090 ;
        RECT -94.465 10.940 -94.295 11.090 ;
        RECT -95.405 10.770 -94.295 10.940 ;
        RECT -95.405 10.565 -95.235 10.770 ;
        RECT -104.385 10.235 -103.455 10.565 ;
        RECT -96.165 10.235 -95.235 10.565 ;
        RECT -104.385 9.710 -104.215 10.235 ;
        RECT -95.405 9.710 -95.235 10.235 ;
        RECT -94.995 9.605 -94.705 10.770 ;
        RECT -94.465 10.565 -94.295 10.770 ;
        RECT -85.485 10.940 -85.315 11.090 ;
        RECT -84.545 10.940 -84.375 11.090 ;
        RECT -85.485 10.770 -84.375 10.940 ;
        RECT -85.485 10.565 -85.315 10.770 ;
        RECT -94.465 10.235 -93.535 10.565 ;
        RECT -86.245 10.235 -85.315 10.565 ;
        RECT -94.465 9.710 -94.295 10.235 ;
        RECT -85.485 9.710 -85.315 10.235 ;
        RECT -85.075 9.605 -84.785 10.770 ;
        RECT -84.545 10.565 -84.375 10.770 ;
        RECT -75.565 10.940 -75.395 11.090 ;
        RECT -74.625 10.940 -74.455 11.090 ;
        RECT -75.565 10.770 -74.455 10.940 ;
        RECT -75.565 10.565 -75.395 10.770 ;
        RECT -84.545 10.235 -83.615 10.565 ;
        RECT -76.325 10.235 -75.395 10.565 ;
        RECT -84.545 9.710 -84.375 10.235 ;
        RECT -75.565 9.710 -75.395 10.235 ;
        RECT -75.155 9.605 -74.865 10.770 ;
        RECT -74.625 10.565 -74.455 10.770 ;
        RECT -65.645 10.940 -65.475 11.090 ;
        RECT -64.705 10.940 -64.535 11.090 ;
        RECT -65.645 10.770 -64.535 10.940 ;
        RECT -65.645 10.565 -65.475 10.770 ;
        RECT -74.625 10.235 -73.695 10.565 ;
        RECT -66.405 10.235 -65.475 10.565 ;
        RECT -74.625 9.710 -74.455 10.235 ;
        RECT -65.645 9.710 -65.475 10.235 ;
        RECT -65.235 9.605 -64.945 10.770 ;
        RECT -64.705 10.565 -64.535 10.770 ;
        RECT -55.725 10.940 -55.555 11.090 ;
        RECT -54.785 10.940 -54.615 11.090 ;
        RECT -55.725 10.770 -54.615 10.940 ;
        RECT -55.725 10.565 -55.555 10.770 ;
        RECT -64.705 10.235 -63.775 10.565 ;
        RECT -56.485 10.235 -55.555 10.565 ;
        RECT -64.705 9.710 -64.535 10.235 ;
        RECT -55.725 9.710 -55.555 10.235 ;
        RECT -55.315 9.605 -55.025 10.770 ;
        RECT -54.785 10.565 -54.615 10.770 ;
        RECT -45.805 10.940 -45.635 11.090 ;
        RECT -44.865 10.940 -44.695 11.090 ;
        RECT -45.805 10.770 -44.695 10.940 ;
        RECT -45.805 10.565 -45.635 10.770 ;
        RECT -54.785 10.235 -53.855 10.565 ;
        RECT -46.565 10.235 -45.635 10.565 ;
        RECT -54.785 9.710 -54.615 10.235 ;
        RECT -45.805 9.710 -45.635 10.235 ;
        RECT -45.395 9.605 -45.105 10.770 ;
        RECT -44.865 10.565 -44.695 10.770 ;
        RECT -35.885 10.940 -35.715 11.090 ;
        RECT -34.945 10.940 -34.775 11.090 ;
        RECT -35.885 10.770 -34.775 10.940 ;
        RECT -35.885 10.565 -35.715 10.770 ;
        RECT -44.865 10.235 -43.935 10.565 ;
        RECT -36.645 10.235 -35.715 10.565 ;
        RECT -44.865 9.710 -44.695 10.235 ;
        RECT -35.885 9.710 -35.715 10.235 ;
        RECT -35.475 9.605 -35.185 10.770 ;
        RECT -34.945 10.565 -34.775 10.770 ;
        RECT -25.965 10.940 -25.795 11.090 ;
        RECT -25.025 10.940 -24.855 11.090 ;
        RECT -25.965 10.770 -24.855 10.940 ;
        RECT -25.965 10.565 -25.795 10.770 ;
        RECT -34.945 10.235 -34.015 10.565 ;
        RECT -26.725 10.235 -25.795 10.565 ;
        RECT -34.945 9.710 -34.775 10.235 ;
        RECT -25.965 9.710 -25.795 10.235 ;
        RECT -25.555 9.605 -25.265 10.770 ;
        RECT -25.025 10.565 -24.855 10.770 ;
        RECT -16.045 10.940 -15.875 11.090 ;
        RECT -15.105 10.940 -14.935 11.090 ;
        RECT -16.045 10.770 -14.935 10.940 ;
        RECT -16.045 10.565 -15.875 10.770 ;
        RECT -25.025 10.235 -24.095 10.565 ;
        RECT -16.805 10.235 -15.875 10.565 ;
        RECT -25.025 9.710 -24.855 10.235 ;
        RECT -16.045 9.710 -15.875 10.235 ;
        RECT -15.635 9.605 -15.345 10.770 ;
        RECT -15.105 10.565 -14.935 10.770 ;
        RECT -6.125 10.940 -5.955 11.090 ;
        RECT -5.185 10.940 -5.015 11.090 ;
        RECT -6.125 10.770 -5.015 10.940 ;
        RECT -6.125 10.565 -5.955 10.770 ;
        RECT -15.105 10.235 -14.175 10.565 ;
        RECT -6.885 10.235 -5.955 10.565 ;
        RECT -15.105 9.710 -14.935 10.235 ;
        RECT -6.125 9.710 -5.955 10.235 ;
        RECT -5.715 9.605 -5.425 10.770 ;
        RECT -5.185 10.565 -5.015 10.770 ;
        RECT 3.795 10.940 3.965 11.090 ;
        RECT 4.735 10.940 4.905 11.090 ;
        RECT 3.795 10.770 4.905 10.940 ;
        RECT 3.795 10.565 3.965 10.770 ;
        RECT -5.185 10.235 -4.255 10.565 ;
        RECT 3.035 10.235 3.965 10.565 ;
        RECT -5.185 9.710 -5.015 10.235 ;
        RECT 3.795 9.710 3.965 10.235 ;
        RECT 4.205 9.605 4.495 10.770 ;
        RECT 4.735 10.565 4.905 10.770 ;
        RECT 13.715 10.940 13.885 11.090 ;
        RECT 14.655 10.940 14.825 11.090 ;
        RECT 13.715 10.770 14.825 10.940 ;
        RECT 13.715 10.565 13.885 10.770 ;
        RECT 4.735 10.235 5.665 10.565 ;
        RECT 12.955 10.235 13.885 10.565 ;
        RECT 4.735 9.710 4.905 10.235 ;
        RECT 13.715 9.710 13.885 10.235 ;
        RECT 14.125 9.605 14.415 10.770 ;
        RECT 14.655 10.565 14.825 10.770 ;
        RECT 23.635 10.940 23.805 11.090 ;
        RECT 23.635 10.770 24.420 10.940 ;
        RECT 23.635 10.565 23.805 10.770 ;
        RECT 14.655 10.235 15.585 10.565 ;
        RECT 22.875 10.235 23.805 10.565 ;
        RECT 14.655 9.710 14.825 10.235 ;
        RECT 23.635 9.710 23.805 10.235 ;
        RECT 24.045 9.605 24.335 10.770 ;
        RECT -289.900 9.195 -286.680 9.365 ;
        RECT -279.980 9.195 -276.760 9.365 ;
        RECT -270.060 9.195 -266.840 9.365 ;
        RECT -260.140 9.195 -256.920 9.365 ;
        RECT -250.220 9.195 -247.000 9.365 ;
        RECT -240.300 9.195 -237.080 9.365 ;
        RECT -230.380 9.195 -227.160 9.365 ;
        RECT -220.460 9.195 -217.240 9.365 ;
        RECT -210.540 9.195 -207.320 9.365 ;
        RECT -200.620 9.195 -197.400 9.365 ;
        RECT -190.700 9.195 -187.480 9.365 ;
        RECT -180.780 9.195 -177.560 9.365 ;
        RECT -170.860 9.195 -167.640 9.365 ;
        RECT -160.940 9.195 -157.720 9.365 ;
        RECT -151.020 9.195 -147.800 9.365 ;
        RECT -141.100 9.195 -137.880 9.365 ;
        RECT -131.180 9.195 -127.960 9.365 ;
        RECT -121.260 9.195 -118.040 9.365 ;
        RECT -111.340 9.195 -108.120 9.365 ;
        RECT -101.420 9.195 -98.200 9.365 ;
        RECT -91.500 9.195 -88.280 9.365 ;
        RECT -81.580 9.195 -78.360 9.365 ;
        RECT -71.660 9.195 -68.440 9.365 ;
        RECT -61.740 9.195 -58.520 9.365 ;
        RECT -51.820 9.195 -48.600 9.365 ;
        RECT -41.900 9.195 -38.680 9.365 ;
        RECT -31.980 9.195 -28.760 9.365 ;
        RECT -22.060 9.195 -18.840 9.365 ;
        RECT -12.140 9.195 -8.920 9.365 ;
        RECT -2.220 9.195 1.000 9.365 ;
        RECT 7.700 9.195 10.920 9.365 ;
        RECT 17.620 9.195 20.840 9.365 ;
        RECT -289.815 8.055 -289.555 9.195 ;
        RECT -288.885 8.055 -288.605 9.195 ;
        RECT -288.435 8.030 -288.145 9.195 ;
        RECT -287.975 8.055 -287.695 9.195 ;
        RECT -287.025 8.055 -286.765 9.195 ;
        RECT -279.895 8.055 -279.635 9.195 ;
        RECT -278.965 8.055 -278.685 9.195 ;
        RECT -278.515 8.030 -278.225 9.195 ;
        RECT -278.055 8.055 -277.775 9.195 ;
        RECT -277.105 8.055 -276.845 9.195 ;
        RECT -269.975 8.055 -269.715 9.195 ;
        RECT -269.045 8.055 -268.765 9.195 ;
        RECT -268.595 8.030 -268.305 9.195 ;
        RECT -268.135 8.055 -267.855 9.195 ;
        RECT -267.185 8.055 -266.925 9.195 ;
        RECT -260.055 8.055 -259.795 9.195 ;
        RECT -259.125 8.055 -258.845 9.195 ;
        RECT -258.675 8.030 -258.385 9.195 ;
        RECT -258.215 8.055 -257.935 9.195 ;
        RECT -257.265 8.055 -257.005 9.195 ;
        RECT -250.135 8.055 -249.875 9.195 ;
        RECT -249.205 8.055 -248.925 9.195 ;
        RECT -248.755 8.030 -248.465 9.195 ;
        RECT -248.295 8.055 -248.015 9.195 ;
        RECT -247.345 8.055 -247.085 9.195 ;
        RECT -240.215 8.055 -239.955 9.195 ;
        RECT -239.285 8.055 -239.005 9.195 ;
        RECT -238.835 8.030 -238.545 9.195 ;
        RECT -238.375 8.055 -238.095 9.195 ;
        RECT -237.425 8.055 -237.165 9.195 ;
        RECT -230.295 8.055 -230.035 9.195 ;
        RECT -229.365 8.055 -229.085 9.195 ;
        RECT -228.915 8.030 -228.625 9.195 ;
        RECT -228.455 8.055 -228.175 9.195 ;
        RECT -227.505 8.055 -227.245 9.195 ;
        RECT -220.375 8.055 -220.115 9.195 ;
        RECT -219.445 8.055 -219.165 9.195 ;
        RECT -218.995 8.030 -218.705 9.195 ;
        RECT -218.535 8.055 -218.255 9.195 ;
        RECT -217.585 8.055 -217.325 9.195 ;
        RECT -210.455 8.055 -210.195 9.195 ;
        RECT -209.525 8.055 -209.245 9.195 ;
        RECT -209.075 8.030 -208.785 9.195 ;
        RECT -208.615 8.055 -208.335 9.195 ;
        RECT -207.665 8.055 -207.405 9.195 ;
        RECT -200.535 8.055 -200.275 9.195 ;
        RECT -199.605 8.055 -199.325 9.195 ;
        RECT -199.155 8.030 -198.865 9.195 ;
        RECT -198.695 8.055 -198.415 9.195 ;
        RECT -197.745 8.055 -197.485 9.195 ;
        RECT -190.615 8.055 -190.355 9.195 ;
        RECT -189.685 8.055 -189.405 9.195 ;
        RECT -189.235 8.030 -188.945 9.195 ;
        RECT -188.775 8.055 -188.495 9.195 ;
        RECT -187.825 8.055 -187.565 9.195 ;
        RECT -180.695 8.055 -180.435 9.195 ;
        RECT -179.765 8.055 -179.485 9.195 ;
        RECT -179.315 8.030 -179.025 9.195 ;
        RECT -178.855 8.055 -178.575 9.195 ;
        RECT -177.905 8.055 -177.645 9.195 ;
        RECT -170.775 8.055 -170.515 9.195 ;
        RECT -169.845 8.055 -169.565 9.195 ;
        RECT -169.395 8.030 -169.105 9.195 ;
        RECT -168.935 8.055 -168.655 9.195 ;
        RECT -167.985 8.055 -167.725 9.195 ;
        RECT -160.855 8.055 -160.595 9.195 ;
        RECT -159.925 8.055 -159.645 9.195 ;
        RECT -159.475 8.030 -159.185 9.195 ;
        RECT -159.015 8.055 -158.735 9.195 ;
        RECT -158.065 8.055 -157.805 9.195 ;
        RECT -150.935 8.055 -150.675 9.195 ;
        RECT -150.005 8.055 -149.725 9.195 ;
        RECT -149.555 8.030 -149.265 9.195 ;
        RECT -149.095 8.055 -148.815 9.195 ;
        RECT -148.145 8.055 -147.885 9.195 ;
        RECT -141.015 8.055 -140.755 9.195 ;
        RECT -140.085 8.055 -139.805 9.195 ;
        RECT -139.635 8.030 -139.345 9.195 ;
        RECT -139.175 8.055 -138.895 9.195 ;
        RECT -138.225 8.055 -137.965 9.195 ;
        RECT -131.095 8.055 -130.835 9.195 ;
        RECT -130.165 8.055 -129.885 9.195 ;
        RECT -129.715 8.030 -129.425 9.195 ;
        RECT -129.255 8.055 -128.975 9.195 ;
        RECT -128.305 8.055 -128.045 9.195 ;
        RECT -121.175 8.055 -120.915 9.195 ;
        RECT -120.245 8.055 -119.965 9.195 ;
        RECT -119.795 8.030 -119.505 9.195 ;
        RECT -119.335 8.055 -119.055 9.195 ;
        RECT -118.385 8.055 -118.125 9.195 ;
        RECT -111.255 8.055 -110.995 9.195 ;
        RECT -110.325 8.055 -110.045 9.195 ;
        RECT -109.875 8.030 -109.585 9.195 ;
        RECT -109.415 8.055 -109.135 9.195 ;
        RECT -108.465 8.055 -108.205 9.195 ;
        RECT -101.335 8.055 -101.075 9.195 ;
        RECT -100.405 8.055 -100.125 9.195 ;
        RECT -99.955 8.030 -99.665 9.195 ;
        RECT -99.495 8.055 -99.215 9.195 ;
        RECT -98.545 8.055 -98.285 9.195 ;
        RECT -91.415 8.055 -91.155 9.195 ;
        RECT -90.485 8.055 -90.205 9.195 ;
        RECT -90.035 8.030 -89.745 9.195 ;
        RECT -89.575 8.055 -89.295 9.195 ;
        RECT -88.625 8.055 -88.365 9.195 ;
        RECT -81.495 8.055 -81.235 9.195 ;
        RECT -80.565 8.055 -80.285 9.195 ;
        RECT -80.115 8.030 -79.825 9.195 ;
        RECT -79.655 8.055 -79.375 9.195 ;
        RECT -78.705 8.055 -78.445 9.195 ;
        RECT -71.575 8.055 -71.315 9.195 ;
        RECT -70.645 8.055 -70.365 9.195 ;
        RECT -70.195 8.030 -69.905 9.195 ;
        RECT -69.735 8.055 -69.455 9.195 ;
        RECT -68.785 8.055 -68.525 9.195 ;
        RECT -61.655 8.055 -61.395 9.195 ;
        RECT -60.725 8.055 -60.445 9.195 ;
        RECT -60.275 8.030 -59.985 9.195 ;
        RECT -59.815 8.055 -59.535 9.195 ;
        RECT -58.865 8.055 -58.605 9.195 ;
        RECT -51.735 8.055 -51.475 9.195 ;
        RECT -50.805 8.055 -50.525 9.195 ;
        RECT -50.355 8.030 -50.065 9.195 ;
        RECT -49.895 8.055 -49.615 9.195 ;
        RECT -48.945 8.055 -48.685 9.195 ;
        RECT -41.815 8.055 -41.555 9.195 ;
        RECT -40.885 8.055 -40.605 9.195 ;
        RECT -40.435 8.030 -40.145 9.195 ;
        RECT -39.975 8.055 -39.695 9.195 ;
        RECT -39.025 8.055 -38.765 9.195 ;
        RECT -31.895 8.055 -31.635 9.195 ;
        RECT -30.965 8.055 -30.685 9.195 ;
        RECT -30.515 8.030 -30.225 9.195 ;
        RECT -30.055 8.055 -29.775 9.195 ;
        RECT -29.105 8.055 -28.845 9.195 ;
        RECT -21.975 8.055 -21.715 9.195 ;
        RECT -21.045 8.055 -20.765 9.195 ;
        RECT -20.595 8.030 -20.305 9.195 ;
        RECT -20.135 8.055 -19.855 9.195 ;
        RECT -19.185 8.055 -18.925 9.195 ;
        RECT -12.055 8.055 -11.795 9.195 ;
        RECT -11.125 8.055 -10.845 9.195 ;
        RECT -10.675 8.030 -10.385 9.195 ;
        RECT -10.215 8.055 -9.935 9.195 ;
        RECT -9.265 8.055 -9.005 9.195 ;
        RECT -2.135 8.055 -1.875 9.195 ;
        RECT -1.205 8.055 -0.925 9.195 ;
        RECT -0.755 8.030 -0.465 9.195 ;
        RECT -0.295 8.055 -0.015 9.195 ;
        RECT 0.655 8.055 0.915 9.195 ;
        RECT 7.785 8.055 8.045 9.195 ;
        RECT 8.715 8.055 8.995 9.195 ;
        RECT 9.165 8.030 9.455 9.195 ;
        RECT 9.625 8.055 9.905 9.195 ;
        RECT 10.575 8.055 10.835 9.195 ;
        RECT 17.705 8.055 17.965 9.195 ;
        RECT 18.635 8.055 18.915 9.195 ;
        RECT 19.085 8.030 19.375 9.195 ;
        RECT 19.545 8.055 19.825 9.195 ;
        RECT 20.495 8.055 20.755 9.195 ;
        RECT -284.855 6.645 -284.595 7.785 ;
        RECT -283.925 6.645 -283.645 7.785 ;
        RECT -283.475 6.645 -283.185 7.810 ;
        RECT -283.015 6.645 -282.735 7.785 ;
        RECT -282.065 6.645 -281.805 7.785 ;
        RECT -274.935 6.645 -274.675 7.785 ;
        RECT -274.005 6.645 -273.725 7.785 ;
        RECT -273.555 6.645 -273.265 7.810 ;
        RECT -273.095 6.645 -272.815 7.785 ;
        RECT -272.145 6.645 -271.885 7.785 ;
        RECT -265.015 6.645 -264.755 7.785 ;
        RECT -264.085 6.645 -263.805 7.785 ;
        RECT -263.635 6.645 -263.345 7.810 ;
        RECT -263.175 6.645 -262.895 7.785 ;
        RECT -262.225 6.645 -261.965 7.785 ;
        RECT -255.095 6.645 -254.835 7.785 ;
        RECT -254.165 6.645 -253.885 7.785 ;
        RECT -253.715 6.645 -253.425 7.810 ;
        RECT -253.255 6.645 -252.975 7.785 ;
        RECT -252.305 6.645 -252.045 7.785 ;
        RECT -245.175 6.645 -244.915 7.785 ;
        RECT -244.245 6.645 -243.965 7.785 ;
        RECT -243.795 6.645 -243.505 7.810 ;
        RECT -243.335 6.645 -243.055 7.785 ;
        RECT -242.385 6.645 -242.125 7.785 ;
        RECT -235.255 6.645 -234.995 7.785 ;
        RECT -234.325 6.645 -234.045 7.785 ;
        RECT -233.875 6.645 -233.585 7.810 ;
        RECT -233.415 6.645 -233.135 7.785 ;
        RECT -232.465 6.645 -232.205 7.785 ;
        RECT -225.335 6.645 -225.075 7.785 ;
        RECT -224.405 6.645 -224.125 7.785 ;
        RECT -223.955 6.645 -223.665 7.810 ;
        RECT -223.495 6.645 -223.215 7.785 ;
        RECT -222.545 6.645 -222.285 7.785 ;
        RECT -215.415 6.645 -215.155 7.785 ;
        RECT -214.485 6.645 -214.205 7.785 ;
        RECT -214.035 6.645 -213.745 7.810 ;
        RECT -213.575 6.645 -213.295 7.785 ;
        RECT -212.625 6.645 -212.365 7.785 ;
        RECT -205.495 6.645 -205.235 7.785 ;
        RECT -204.565 6.645 -204.285 7.785 ;
        RECT -204.115 6.645 -203.825 7.810 ;
        RECT -203.655 6.645 -203.375 7.785 ;
        RECT -202.705 6.645 -202.445 7.785 ;
        RECT -195.575 6.645 -195.315 7.785 ;
        RECT -194.645 6.645 -194.365 7.785 ;
        RECT -194.195 6.645 -193.905 7.810 ;
        RECT -193.735 6.645 -193.455 7.785 ;
        RECT -192.785 6.645 -192.525 7.785 ;
        RECT -185.655 6.645 -185.395 7.785 ;
        RECT -184.725 6.645 -184.445 7.785 ;
        RECT -184.275 6.645 -183.985 7.810 ;
        RECT -183.815 6.645 -183.535 7.785 ;
        RECT -182.865 6.645 -182.605 7.785 ;
        RECT -175.735 6.645 -175.475 7.785 ;
        RECT -174.805 6.645 -174.525 7.785 ;
        RECT -174.355 6.645 -174.065 7.810 ;
        RECT -173.895 6.645 -173.615 7.785 ;
        RECT -172.945 6.645 -172.685 7.785 ;
        RECT -165.815 6.645 -165.555 7.785 ;
        RECT -164.885 6.645 -164.605 7.785 ;
        RECT -164.435 6.645 -164.145 7.810 ;
        RECT -163.975 6.645 -163.695 7.785 ;
        RECT -163.025 6.645 -162.765 7.785 ;
        RECT -155.895 6.645 -155.635 7.785 ;
        RECT -154.965 6.645 -154.685 7.785 ;
        RECT -154.515 6.645 -154.225 7.810 ;
        RECT -154.055 6.645 -153.775 7.785 ;
        RECT -153.105 6.645 -152.845 7.785 ;
        RECT -145.975 6.645 -145.715 7.785 ;
        RECT -145.045 6.645 -144.765 7.785 ;
        RECT -144.595 6.645 -144.305 7.810 ;
        RECT -144.135 6.645 -143.855 7.785 ;
        RECT -143.185 6.645 -142.925 7.785 ;
        RECT -136.055 6.645 -135.795 7.785 ;
        RECT -135.125 6.645 -134.845 7.785 ;
        RECT -134.675 6.645 -134.385 7.810 ;
        RECT -134.215 6.645 -133.935 7.785 ;
        RECT -133.265 6.645 -133.005 7.785 ;
        RECT -126.135 6.645 -125.875 7.785 ;
        RECT -125.205 6.645 -124.925 7.785 ;
        RECT -124.755 6.645 -124.465 7.810 ;
        RECT -124.295 6.645 -124.015 7.785 ;
        RECT -123.345 6.645 -123.085 7.785 ;
        RECT -116.215 6.645 -115.955 7.785 ;
        RECT -115.285 6.645 -115.005 7.785 ;
        RECT -114.835 6.645 -114.545 7.810 ;
        RECT -114.375 6.645 -114.095 7.785 ;
        RECT -113.425 6.645 -113.165 7.785 ;
        RECT -106.295 6.645 -106.035 7.785 ;
        RECT -105.365 6.645 -105.085 7.785 ;
        RECT -104.915 6.645 -104.625 7.810 ;
        RECT -104.455 6.645 -104.175 7.785 ;
        RECT -103.505 6.645 -103.245 7.785 ;
        RECT -96.375 6.645 -96.115 7.785 ;
        RECT -95.445 6.645 -95.165 7.785 ;
        RECT -94.995 6.645 -94.705 7.810 ;
        RECT -94.535 6.645 -94.255 7.785 ;
        RECT -93.585 6.645 -93.325 7.785 ;
        RECT -86.455 6.645 -86.195 7.785 ;
        RECT -85.525 6.645 -85.245 7.785 ;
        RECT -85.075 6.645 -84.785 7.810 ;
        RECT -84.615 6.645 -84.335 7.785 ;
        RECT -83.665 6.645 -83.405 7.785 ;
        RECT -76.535 6.645 -76.275 7.785 ;
        RECT -75.605 6.645 -75.325 7.785 ;
        RECT -75.155 6.645 -74.865 7.810 ;
        RECT -74.695 6.645 -74.415 7.785 ;
        RECT -73.745 6.645 -73.485 7.785 ;
        RECT -66.615 6.645 -66.355 7.785 ;
        RECT -65.685 6.645 -65.405 7.785 ;
        RECT -65.235 6.645 -64.945 7.810 ;
        RECT -64.775 6.645 -64.495 7.785 ;
        RECT -63.825 6.645 -63.565 7.785 ;
        RECT -56.695 6.645 -56.435 7.785 ;
        RECT -55.765 6.645 -55.485 7.785 ;
        RECT -55.315 6.645 -55.025 7.810 ;
        RECT -54.855 6.645 -54.575 7.785 ;
        RECT -53.905 6.645 -53.645 7.785 ;
        RECT -46.775 6.645 -46.515 7.785 ;
        RECT -45.845 6.645 -45.565 7.785 ;
        RECT -45.395 6.645 -45.105 7.810 ;
        RECT -44.935 6.645 -44.655 7.785 ;
        RECT -43.985 6.645 -43.725 7.785 ;
        RECT -36.855 6.645 -36.595 7.785 ;
        RECT -35.925 6.645 -35.645 7.785 ;
        RECT -35.475 6.645 -35.185 7.810 ;
        RECT -35.015 6.645 -34.735 7.785 ;
        RECT -34.065 6.645 -33.805 7.785 ;
        RECT -26.935 6.645 -26.675 7.785 ;
        RECT -26.005 6.645 -25.725 7.785 ;
        RECT -25.555 6.645 -25.265 7.810 ;
        RECT -25.095 6.645 -24.815 7.785 ;
        RECT -24.145 6.645 -23.885 7.785 ;
        RECT -17.015 6.645 -16.755 7.785 ;
        RECT -16.085 6.645 -15.805 7.785 ;
        RECT -15.635 6.645 -15.345 7.810 ;
        RECT -15.175 6.645 -14.895 7.785 ;
        RECT -14.225 6.645 -13.965 7.785 ;
        RECT -7.095 6.645 -6.835 7.785 ;
        RECT -6.165 6.645 -5.885 7.785 ;
        RECT -5.715 6.645 -5.425 7.810 ;
        RECT -5.255 6.645 -4.975 7.785 ;
        RECT -4.305 6.645 -4.045 7.785 ;
        RECT 2.825 6.645 3.085 7.785 ;
        RECT 3.755 6.645 4.035 7.785 ;
        RECT 4.205 6.645 4.495 7.810 ;
        RECT 4.665 6.645 4.945 7.785 ;
        RECT 5.615 6.645 5.875 7.785 ;
        RECT 12.745 6.645 13.005 7.785 ;
        RECT 13.675 6.645 13.955 7.785 ;
        RECT 14.125 6.645 14.415 7.810 ;
        RECT 14.585 6.645 14.865 7.785 ;
        RECT 15.535 6.645 15.795 7.785 ;
        RECT 22.665 6.645 22.925 7.785 ;
        RECT 23.595 6.645 23.875 7.785 ;
        RECT 24.045 6.645 24.335 7.810 ;
        RECT -284.940 6.475 -281.720 6.645 ;
        RECT -275.020 6.475 -271.800 6.645 ;
        RECT -265.100 6.475 -261.880 6.645 ;
        RECT -255.180 6.475 -251.960 6.645 ;
        RECT -245.260 6.475 -242.040 6.645 ;
        RECT -235.340 6.475 -232.120 6.645 ;
        RECT -225.420 6.475 -222.200 6.645 ;
        RECT -215.500 6.475 -212.280 6.645 ;
        RECT -205.580 6.475 -202.360 6.645 ;
        RECT -195.660 6.475 -192.440 6.645 ;
        RECT -185.740 6.475 -182.520 6.645 ;
        RECT -175.820 6.475 -172.600 6.645 ;
        RECT -165.900 6.475 -162.680 6.645 ;
        RECT -155.980 6.475 -152.760 6.645 ;
        RECT -146.060 6.475 -142.840 6.645 ;
        RECT -136.140 6.475 -132.920 6.645 ;
        RECT -126.220 6.475 -123.000 6.645 ;
        RECT -116.300 6.475 -113.080 6.645 ;
        RECT -106.380 6.475 -103.160 6.645 ;
        RECT -96.460 6.475 -93.240 6.645 ;
        RECT -86.540 6.475 -83.320 6.645 ;
        RECT -76.620 6.475 -73.400 6.645 ;
        RECT -66.700 6.475 -63.480 6.645 ;
        RECT -56.780 6.475 -53.560 6.645 ;
        RECT -46.860 6.475 -43.640 6.645 ;
        RECT -36.940 6.475 -33.720 6.645 ;
        RECT -27.020 6.475 -23.800 6.645 ;
        RECT -17.100 6.475 -13.880 6.645 ;
        RECT -7.180 6.475 -3.960 6.645 ;
        RECT 2.740 6.475 5.960 6.645 ;
        RECT 12.660 6.475 15.880 6.645 ;
        RECT 22.580 6.475 24.420 6.645 ;
        RECT -288.845 6.060 -288.675 6.130 ;
        RECT -287.905 6.060 -287.735 6.130 ;
        RECT -288.845 5.890 -287.735 6.060 ;
        RECT -288.845 5.605 -288.675 5.890 ;
        RECT -289.605 5.275 -288.675 5.605 ;
        RECT -288.845 4.750 -288.675 5.275 ;
        RECT -288.435 4.725 -288.145 5.890 ;
        RECT -287.905 5.605 -287.735 5.890 ;
        RECT -278.925 6.060 -278.755 6.130 ;
        RECT -277.985 6.060 -277.815 6.130 ;
        RECT -278.925 5.890 -277.815 6.060 ;
        RECT -278.925 5.605 -278.755 5.890 ;
        RECT -287.905 5.275 -286.975 5.605 ;
        RECT -279.685 5.275 -278.755 5.605 ;
        RECT -287.905 4.750 -287.735 5.275 ;
        RECT -278.925 4.750 -278.755 5.275 ;
        RECT -278.515 4.725 -278.225 5.890 ;
        RECT -277.985 5.605 -277.815 5.890 ;
        RECT -269.005 6.060 -268.835 6.130 ;
        RECT -268.065 6.060 -267.895 6.130 ;
        RECT -269.005 5.890 -267.895 6.060 ;
        RECT -269.005 5.605 -268.835 5.890 ;
        RECT -277.985 5.275 -277.055 5.605 ;
        RECT -269.765 5.275 -268.835 5.605 ;
        RECT -277.985 4.750 -277.815 5.275 ;
        RECT -269.005 4.750 -268.835 5.275 ;
        RECT -268.595 4.725 -268.305 5.890 ;
        RECT -268.065 5.605 -267.895 5.890 ;
        RECT -259.085 6.060 -258.915 6.130 ;
        RECT -258.145 6.060 -257.975 6.130 ;
        RECT -259.085 5.890 -257.975 6.060 ;
        RECT -259.085 5.605 -258.915 5.890 ;
        RECT -268.065 5.275 -267.135 5.605 ;
        RECT -259.845 5.275 -258.915 5.605 ;
        RECT -268.065 4.750 -267.895 5.275 ;
        RECT -259.085 4.750 -258.915 5.275 ;
        RECT -258.675 4.725 -258.385 5.890 ;
        RECT -258.145 5.605 -257.975 5.890 ;
        RECT -249.165 6.060 -248.995 6.130 ;
        RECT -248.225 6.060 -248.055 6.130 ;
        RECT -249.165 5.890 -248.055 6.060 ;
        RECT -249.165 5.605 -248.995 5.890 ;
        RECT -258.145 5.275 -257.215 5.605 ;
        RECT -249.925 5.275 -248.995 5.605 ;
        RECT -258.145 4.750 -257.975 5.275 ;
        RECT -249.165 4.750 -248.995 5.275 ;
        RECT -248.755 4.725 -248.465 5.890 ;
        RECT -248.225 5.605 -248.055 5.890 ;
        RECT -239.245 6.060 -239.075 6.130 ;
        RECT -238.305 6.060 -238.135 6.130 ;
        RECT -239.245 5.890 -238.135 6.060 ;
        RECT -239.245 5.605 -239.075 5.890 ;
        RECT -248.225 5.275 -247.295 5.605 ;
        RECT -240.005 5.275 -239.075 5.605 ;
        RECT -248.225 4.750 -248.055 5.275 ;
        RECT -239.245 4.750 -239.075 5.275 ;
        RECT -238.835 4.725 -238.545 5.890 ;
        RECT -238.305 5.605 -238.135 5.890 ;
        RECT -229.325 6.060 -229.155 6.130 ;
        RECT -228.385 6.060 -228.215 6.130 ;
        RECT -229.325 5.890 -228.215 6.060 ;
        RECT -229.325 5.605 -229.155 5.890 ;
        RECT -238.305 5.275 -237.375 5.605 ;
        RECT -230.085 5.275 -229.155 5.605 ;
        RECT -238.305 4.750 -238.135 5.275 ;
        RECT -229.325 4.750 -229.155 5.275 ;
        RECT -228.915 4.725 -228.625 5.890 ;
        RECT -228.385 5.605 -228.215 5.890 ;
        RECT -219.405 6.060 -219.235 6.130 ;
        RECT -218.465 6.060 -218.295 6.130 ;
        RECT -219.405 5.890 -218.295 6.060 ;
        RECT -219.405 5.605 -219.235 5.890 ;
        RECT -228.385 5.275 -227.455 5.605 ;
        RECT -220.165 5.275 -219.235 5.605 ;
        RECT -228.385 4.750 -228.215 5.275 ;
        RECT -219.405 4.750 -219.235 5.275 ;
        RECT -218.995 4.725 -218.705 5.890 ;
        RECT -218.465 5.605 -218.295 5.890 ;
        RECT -209.485 6.060 -209.315 6.130 ;
        RECT -208.545 6.060 -208.375 6.130 ;
        RECT -209.485 5.890 -208.375 6.060 ;
        RECT -209.485 5.605 -209.315 5.890 ;
        RECT -218.465 5.275 -217.535 5.605 ;
        RECT -210.245 5.275 -209.315 5.605 ;
        RECT -218.465 4.750 -218.295 5.275 ;
        RECT -209.485 4.750 -209.315 5.275 ;
        RECT -209.075 4.725 -208.785 5.890 ;
        RECT -208.545 5.605 -208.375 5.890 ;
        RECT -199.565 6.060 -199.395 6.130 ;
        RECT -198.625 6.060 -198.455 6.130 ;
        RECT -199.565 5.890 -198.455 6.060 ;
        RECT -199.565 5.605 -199.395 5.890 ;
        RECT -208.545 5.275 -207.615 5.605 ;
        RECT -200.325 5.275 -199.395 5.605 ;
        RECT -208.545 4.750 -208.375 5.275 ;
        RECT -199.565 4.750 -199.395 5.275 ;
        RECT -199.155 4.725 -198.865 5.890 ;
        RECT -198.625 5.605 -198.455 5.890 ;
        RECT -189.645 6.060 -189.475 6.130 ;
        RECT -188.705 6.060 -188.535 6.130 ;
        RECT -189.645 5.890 -188.535 6.060 ;
        RECT -189.645 5.605 -189.475 5.890 ;
        RECT -198.625 5.275 -197.695 5.605 ;
        RECT -190.405 5.275 -189.475 5.605 ;
        RECT -198.625 4.750 -198.455 5.275 ;
        RECT -189.645 4.750 -189.475 5.275 ;
        RECT -189.235 4.725 -188.945 5.890 ;
        RECT -188.705 5.605 -188.535 5.890 ;
        RECT -179.725 6.060 -179.555 6.130 ;
        RECT -178.785 6.060 -178.615 6.130 ;
        RECT -179.725 5.890 -178.615 6.060 ;
        RECT -179.725 5.605 -179.555 5.890 ;
        RECT -188.705 5.275 -187.775 5.605 ;
        RECT -180.485 5.275 -179.555 5.605 ;
        RECT -188.705 4.750 -188.535 5.275 ;
        RECT -179.725 4.750 -179.555 5.275 ;
        RECT -179.315 4.725 -179.025 5.890 ;
        RECT -178.785 5.605 -178.615 5.890 ;
        RECT -169.805 6.060 -169.635 6.130 ;
        RECT -168.865 6.060 -168.695 6.130 ;
        RECT -169.805 5.890 -168.695 6.060 ;
        RECT -169.805 5.605 -169.635 5.890 ;
        RECT -178.785 5.275 -177.855 5.605 ;
        RECT -170.565 5.275 -169.635 5.605 ;
        RECT -178.785 4.750 -178.615 5.275 ;
        RECT -169.805 4.750 -169.635 5.275 ;
        RECT -169.395 4.725 -169.105 5.890 ;
        RECT -168.865 5.605 -168.695 5.890 ;
        RECT -159.885 6.060 -159.715 6.130 ;
        RECT -158.945 6.060 -158.775 6.130 ;
        RECT -159.885 5.890 -158.775 6.060 ;
        RECT -159.885 5.605 -159.715 5.890 ;
        RECT -168.865 5.275 -167.935 5.605 ;
        RECT -160.645 5.275 -159.715 5.605 ;
        RECT -168.865 4.750 -168.695 5.275 ;
        RECT -159.885 4.750 -159.715 5.275 ;
        RECT -159.475 4.725 -159.185 5.890 ;
        RECT -158.945 5.605 -158.775 5.890 ;
        RECT -149.965 6.060 -149.795 6.130 ;
        RECT -149.025 6.060 -148.855 6.130 ;
        RECT -149.965 5.890 -148.855 6.060 ;
        RECT -149.965 5.605 -149.795 5.890 ;
        RECT -158.945 5.275 -158.015 5.605 ;
        RECT -150.725 5.275 -149.795 5.605 ;
        RECT -158.945 4.750 -158.775 5.275 ;
        RECT -149.965 4.750 -149.795 5.275 ;
        RECT -149.555 4.725 -149.265 5.890 ;
        RECT -149.025 5.605 -148.855 5.890 ;
        RECT -140.045 6.060 -139.875 6.130 ;
        RECT -139.105 6.060 -138.935 6.130 ;
        RECT -140.045 5.890 -138.935 6.060 ;
        RECT -140.045 5.605 -139.875 5.890 ;
        RECT -149.025 5.275 -148.095 5.605 ;
        RECT -140.805 5.275 -139.875 5.605 ;
        RECT -149.025 4.750 -148.855 5.275 ;
        RECT -140.045 4.750 -139.875 5.275 ;
        RECT -139.635 4.725 -139.345 5.890 ;
        RECT -139.105 5.605 -138.935 5.890 ;
        RECT -130.125 6.060 -129.955 6.130 ;
        RECT -129.185 6.060 -129.015 6.130 ;
        RECT -130.125 5.890 -129.015 6.060 ;
        RECT -130.125 5.605 -129.955 5.890 ;
        RECT -139.105 5.275 -138.175 5.605 ;
        RECT -130.885 5.275 -129.955 5.605 ;
        RECT -139.105 4.750 -138.935 5.275 ;
        RECT -130.125 4.750 -129.955 5.275 ;
        RECT -129.715 4.725 -129.425 5.890 ;
        RECT -129.185 5.605 -129.015 5.890 ;
        RECT -120.205 6.060 -120.035 6.130 ;
        RECT -119.265 6.060 -119.095 6.130 ;
        RECT -120.205 5.890 -119.095 6.060 ;
        RECT -120.205 5.605 -120.035 5.890 ;
        RECT -129.185 5.275 -128.255 5.605 ;
        RECT -120.965 5.275 -120.035 5.605 ;
        RECT -129.185 4.750 -129.015 5.275 ;
        RECT -120.205 4.750 -120.035 5.275 ;
        RECT -119.795 4.725 -119.505 5.890 ;
        RECT -119.265 5.605 -119.095 5.890 ;
        RECT -110.285 6.060 -110.115 6.130 ;
        RECT -109.345 6.060 -109.175 6.130 ;
        RECT -110.285 5.890 -109.175 6.060 ;
        RECT -110.285 5.605 -110.115 5.890 ;
        RECT -119.265 5.275 -118.335 5.605 ;
        RECT -111.045 5.275 -110.115 5.605 ;
        RECT -119.265 4.750 -119.095 5.275 ;
        RECT -110.285 4.750 -110.115 5.275 ;
        RECT -109.875 4.725 -109.585 5.890 ;
        RECT -109.345 5.605 -109.175 5.890 ;
        RECT -100.365 6.060 -100.195 6.130 ;
        RECT -99.425 6.060 -99.255 6.130 ;
        RECT -100.365 5.890 -99.255 6.060 ;
        RECT -100.365 5.605 -100.195 5.890 ;
        RECT -109.345 5.275 -108.415 5.605 ;
        RECT -101.125 5.275 -100.195 5.605 ;
        RECT -109.345 4.750 -109.175 5.275 ;
        RECT -100.365 4.750 -100.195 5.275 ;
        RECT -99.955 4.725 -99.665 5.890 ;
        RECT -99.425 5.605 -99.255 5.890 ;
        RECT -90.445 6.060 -90.275 6.130 ;
        RECT -89.505 6.060 -89.335 6.130 ;
        RECT -90.445 5.890 -89.335 6.060 ;
        RECT -90.445 5.605 -90.275 5.890 ;
        RECT -99.425 5.275 -98.495 5.605 ;
        RECT -91.205 5.275 -90.275 5.605 ;
        RECT -99.425 4.750 -99.255 5.275 ;
        RECT -90.445 4.750 -90.275 5.275 ;
        RECT -90.035 4.725 -89.745 5.890 ;
        RECT -89.505 5.605 -89.335 5.890 ;
        RECT -80.525 6.060 -80.355 6.130 ;
        RECT -79.585 6.060 -79.415 6.130 ;
        RECT -80.525 5.890 -79.415 6.060 ;
        RECT -80.525 5.605 -80.355 5.890 ;
        RECT -89.505 5.275 -88.575 5.605 ;
        RECT -81.285 5.275 -80.355 5.605 ;
        RECT -89.505 4.750 -89.335 5.275 ;
        RECT -80.525 4.750 -80.355 5.275 ;
        RECT -80.115 4.725 -79.825 5.890 ;
        RECT -79.585 5.605 -79.415 5.890 ;
        RECT -70.605 6.060 -70.435 6.130 ;
        RECT -69.665 6.060 -69.495 6.130 ;
        RECT -70.605 5.890 -69.495 6.060 ;
        RECT -70.605 5.605 -70.435 5.890 ;
        RECT -79.585 5.275 -78.655 5.605 ;
        RECT -71.365 5.275 -70.435 5.605 ;
        RECT -79.585 4.750 -79.415 5.275 ;
        RECT -70.605 4.750 -70.435 5.275 ;
        RECT -70.195 4.725 -69.905 5.890 ;
        RECT -69.665 5.605 -69.495 5.890 ;
        RECT -60.685 6.060 -60.515 6.130 ;
        RECT -59.745 6.060 -59.575 6.130 ;
        RECT -60.685 5.890 -59.575 6.060 ;
        RECT -60.685 5.605 -60.515 5.890 ;
        RECT -69.665 5.275 -68.735 5.605 ;
        RECT -61.445 5.275 -60.515 5.605 ;
        RECT -69.665 4.750 -69.495 5.275 ;
        RECT -60.685 4.750 -60.515 5.275 ;
        RECT -60.275 4.725 -59.985 5.890 ;
        RECT -59.745 5.605 -59.575 5.890 ;
        RECT -50.765 6.060 -50.595 6.130 ;
        RECT -49.825 6.060 -49.655 6.130 ;
        RECT -50.765 5.890 -49.655 6.060 ;
        RECT -50.765 5.605 -50.595 5.890 ;
        RECT -59.745 5.275 -58.815 5.605 ;
        RECT -51.525 5.275 -50.595 5.605 ;
        RECT -59.745 4.750 -59.575 5.275 ;
        RECT -50.765 4.750 -50.595 5.275 ;
        RECT -50.355 4.725 -50.065 5.890 ;
        RECT -49.825 5.605 -49.655 5.890 ;
        RECT -40.845 6.060 -40.675 6.130 ;
        RECT -39.905 6.060 -39.735 6.130 ;
        RECT -40.845 5.890 -39.735 6.060 ;
        RECT -40.845 5.605 -40.675 5.890 ;
        RECT -49.825 5.275 -48.895 5.605 ;
        RECT -41.605 5.275 -40.675 5.605 ;
        RECT -49.825 4.750 -49.655 5.275 ;
        RECT -40.845 4.750 -40.675 5.275 ;
        RECT -40.435 4.725 -40.145 5.890 ;
        RECT -39.905 5.605 -39.735 5.890 ;
        RECT -30.925 6.060 -30.755 6.130 ;
        RECT -29.985 6.060 -29.815 6.130 ;
        RECT -30.925 5.890 -29.815 6.060 ;
        RECT -30.925 5.605 -30.755 5.890 ;
        RECT -39.905 5.275 -38.975 5.605 ;
        RECT -31.685 5.275 -30.755 5.605 ;
        RECT -39.905 4.750 -39.735 5.275 ;
        RECT -30.925 4.750 -30.755 5.275 ;
        RECT -30.515 4.725 -30.225 5.890 ;
        RECT -29.985 5.605 -29.815 5.890 ;
        RECT -21.005 6.060 -20.835 6.130 ;
        RECT -20.065 6.060 -19.895 6.130 ;
        RECT -21.005 5.890 -19.895 6.060 ;
        RECT -21.005 5.605 -20.835 5.890 ;
        RECT -29.985 5.275 -29.055 5.605 ;
        RECT -21.765 5.275 -20.835 5.605 ;
        RECT -29.985 4.750 -29.815 5.275 ;
        RECT -21.005 4.750 -20.835 5.275 ;
        RECT -20.595 4.725 -20.305 5.890 ;
        RECT -20.065 5.605 -19.895 5.890 ;
        RECT -11.085 6.060 -10.915 6.130 ;
        RECT -10.145 6.060 -9.975 6.130 ;
        RECT -11.085 5.890 -9.975 6.060 ;
        RECT -11.085 5.605 -10.915 5.890 ;
        RECT -20.065 5.275 -19.135 5.605 ;
        RECT -11.845 5.275 -10.915 5.605 ;
        RECT -20.065 4.750 -19.895 5.275 ;
        RECT -11.085 4.750 -10.915 5.275 ;
        RECT -10.675 4.725 -10.385 5.890 ;
        RECT -10.145 5.605 -9.975 5.890 ;
        RECT -1.165 6.060 -0.995 6.130 ;
        RECT -0.225 6.060 -0.055 6.130 ;
        RECT -1.165 5.890 -0.055 6.060 ;
        RECT -1.165 5.605 -0.995 5.890 ;
        RECT -10.145 5.275 -9.215 5.605 ;
        RECT -1.925 5.275 -0.995 5.605 ;
        RECT -10.145 4.750 -9.975 5.275 ;
        RECT -1.165 4.750 -0.995 5.275 ;
        RECT -0.755 4.725 -0.465 5.890 ;
        RECT -0.225 5.605 -0.055 5.890 ;
        RECT 8.755 6.060 8.925 6.130 ;
        RECT 9.695 6.060 9.865 6.130 ;
        RECT 8.755 5.890 9.865 6.060 ;
        RECT 8.755 5.605 8.925 5.890 ;
        RECT -0.225 5.275 0.705 5.605 ;
        RECT 7.995 5.275 8.925 5.605 ;
        RECT -0.225 4.750 -0.055 5.275 ;
        RECT 8.755 4.750 8.925 5.275 ;
        RECT 9.165 4.725 9.455 5.890 ;
        RECT 9.695 5.605 9.865 5.890 ;
        RECT 18.675 6.060 18.845 6.130 ;
        RECT 19.615 6.060 19.785 6.130 ;
        RECT 18.675 5.890 19.785 6.060 ;
        RECT 18.675 5.605 18.845 5.890 ;
        RECT 9.695 5.275 10.625 5.605 ;
        RECT 17.915 5.275 18.845 5.605 ;
        RECT 9.695 4.750 9.865 5.275 ;
        RECT 18.675 4.750 18.845 5.275 ;
        RECT 19.085 4.725 19.375 5.890 ;
        RECT 19.615 5.605 19.785 5.890 ;
        RECT 19.615 5.275 20.545 5.605 ;
        RECT 19.615 4.750 19.785 5.275 ;
        RECT -283.525 -78.010 -283.355 -77.860 ;
        RECT -282.585 -78.010 -282.415 -77.860 ;
        RECT -283.525 -78.180 -282.415 -78.010 ;
        RECT -283.525 -78.385 -283.355 -78.180 ;
        RECT -284.285 -78.715 -283.355 -78.385 ;
        RECT -283.525 -79.240 -283.355 -78.715 ;
        RECT -283.115 -79.345 -282.825 -78.180 ;
        RECT -282.585 -78.385 -282.415 -78.180 ;
        RECT -273.605 -78.010 -273.435 -77.860 ;
        RECT -272.665 -78.010 -272.495 -77.860 ;
        RECT -273.605 -78.180 -272.495 -78.010 ;
        RECT -273.605 -78.385 -273.435 -78.180 ;
        RECT -282.585 -78.715 -281.655 -78.385 ;
        RECT -274.365 -78.715 -273.435 -78.385 ;
        RECT -282.585 -79.240 -282.415 -78.715 ;
        RECT -273.605 -79.240 -273.435 -78.715 ;
        RECT -273.195 -79.345 -272.905 -78.180 ;
        RECT -272.665 -78.385 -272.495 -78.180 ;
        RECT -263.685 -78.010 -263.515 -77.860 ;
        RECT -262.745 -78.010 -262.575 -77.860 ;
        RECT -263.685 -78.180 -262.575 -78.010 ;
        RECT -263.685 -78.385 -263.515 -78.180 ;
        RECT -272.665 -78.715 -271.735 -78.385 ;
        RECT -264.445 -78.715 -263.515 -78.385 ;
        RECT -272.665 -79.240 -272.495 -78.715 ;
        RECT -263.685 -79.240 -263.515 -78.715 ;
        RECT -263.275 -79.345 -262.985 -78.180 ;
        RECT -262.745 -78.385 -262.575 -78.180 ;
        RECT -253.765 -78.010 -253.595 -77.860 ;
        RECT -252.825 -78.010 -252.655 -77.860 ;
        RECT -253.765 -78.180 -252.655 -78.010 ;
        RECT -253.765 -78.385 -253.595 -78.180 ;
        RECT -262.745 -78.715 -261.815 -78.385 ;
        RECT -254.525 -78.715 -253.595 -78.385 ;
        RECT -262.745 -79.240 -262.575 -78.715 ;
        RECT -253.765 -79.240 -253.595 -78.715 ;
        RECT -253.355 -79.345 -253.065 -78.180 ;
        RECT -252.825 -78.385 -252.655 -78.180 ;
        RECT -243.845 -78.010 -243.675 -77.860 ;
        RECT -242.905 -78.010 -242.735 -77.860 ;
        RECT -243.845 -78.180 -242.735 -78.010 ;
        RECT -243.845 -78.385 -243.675 -78.180 ;
        RECT -252.825 -78.715 -251.895 -78.385 ;
        RECT -244.605 -78.715 -243.675 -78.385 ;
        RECT -252.825 -79.240 -252.655 -78.715 ;
        RECT -243.845 -79.240 -243.675 -78.715 ;
        RECT -243.435 -79.345 -243.145 -78.180 ;
        RECT -242.905 -78.385 -242.735 -78.180 ;
        RECT -233.925 -78.010 -233.755 -77.860 ;
        RECT -232.985 -78.010 -232.815 -77.860 ;
        RECT -233.925 -78.180 -232.815 -78.010 ;
        RECT -233.925 -78.385 -233.755 -78.180 ;
        RECT -242.905 -78.715 -241.975 -78.385 ;
        RECT -234.685 -78.715 -233.755 -78.385 ;
        RECT -242.905 -79.240 -242.735 -78.715 ;
        RECT -233.925 -79.240 -233.755 -78.715 ;
        RECT -233.515 -79.345 -233.225 -78.180 ;
        RECT -232.985 -78.385 -232.815 -78.180 ;
        RECT -224.005 -78.010 -223.835 -77.860 ;
        RECT -223.065 -78.010 -222.895 -77.860 ;
        RECT -224.005 -78.180 -222.895 -78.010 ;
        RECT -224.005 -78.385 -223.835 -78.180 ;
        RECT -232.985 -78.715 -232.055 -78.385 ;
        RECT -224.765 -78.715 -223.835 -78.385 ;
        RECT -232.985 -79.240 -232.815 -78.715 ;
        RECT -224.005 -79.240 -223.835 -78.715 ;
        RECT -223.595 -79.345 -223.305 -78.180 ;
        RECT -223.065 -78.385 -222.895 -78.180 ;
        RECT -214.085 -78.010 -213.915 -77.860 ;
        RECT -213.145 -78.010 -212.975 -77.860 ;
        RECT -214.085 -78.180 -212.975 -78.010 ;
        RECT -214.085 -78.385 -213.915 -78.180 ;
        RECT -223.065 -78.715 -222.135 -78.385 ;
        RECT -214.845 -78.715 -213.915 -78.385 ;
        RECT -223.065 -79.240 -222.895 -78.715 ;
        RECT -214.085 -79.240 -213.915 -78.715 ;
        RECT -213.675 -79.345 -213.385 -78.180 ;
        RECT -213.145 -78.385 -212.975 -78.180 ;
        RECT -204.165 -78.010 -203.995 -77.860 ;
        RECT -203.225 -78.010 -203.055 -77.860 ;
        RECT -204.165 -78.180 -203.055 -78.010 ;
        RECT -204.165 -78.385 -203.995 -78.180 ;
        RECT -213.145 -78.715 -212.215 -78.385 ;
        RECT -204.925 -78.715 -203.995 -78.385 ;
        RECT -213.145 -79.240 -212.975 -78.715 ;
        RECT -204.165 -79.240 -203.995 -78.715 ;
        RECT -203.755 -79.345 -203.465 -78.180 ;
        RECT -203.225 -78.385 -203.055 -78.180 ;
        RECT -194.245 -78.010 -194.075 -77.860 ;
        RECT -193.305 -78.010 -193.135 -77.860 ;
        RECT -194.245 -78.180 -193.135 -78.010 ;
        RECT -194.245 -78.385 -194.075 -78.180 ;
        RECT -203.225 -78.715 -202.295 -78.385 ;
        RECT -195.005 -78.715 -194.075 -78.385 ;
        RECT -203.225 -79.240 -203.055 -78.715 ;
        RECT -194.245 -79.240 -194.075 -78.715 ;
        RECT -193.835 -79.345 -193.545 -78.180 ;
        RECT -193.305 -78.385 -193.135 -78.180 ;
        RECT -184.325 -78.010 -184.155 -77.860 ;
        RECT -183.385 -78.010 -183.215 -77.860 ;
        RECT -184.325 -78.180 -183.215 -78.010 ;
        RECT -184.325 -78.385 -184.155 -78.180 ;
        RECT -193.305 -78.715 -192.375 -78.385 ;
        RECT -185.085 -78.715 -184.155 -78.385 ;
        RECT -193.305 -79.240 -193.135 -78.715 ;
        RECT -184.325 -79.240 -184.155 -78.715 ;
        RECT -183.915 -79.345 -183.625 -78.180 ;
        RECT -183.385 -78.385 -183.215 -78.180 ;
        RECT -174.405 -78.010 -174.235 -77.860 ;
        RECT -173.465 -78.010 -173.295 -77.860 ;
        RECT -174.405 -78.180 -173.295 -78.010 ;
        RECT -174.405 -78.385 -174.235 -78.180 ;
        RECT -183.385 -78.715 -182.455 -78.385 ;
        RECT -175.165 -78.715 -174.235 -78.385 ;
        RECT -183.385 -79.240 -183.215 -78.715 ;
        RECT -174.405 -79.240 -174.235 -78.715 ;
        RECT -173.995 -79.345 -173.705 -78.180 ;
        RECT -173.465 -78.385 -173.295 -78.180 ;
        RECT -164.485 -78.010 -164.315 -77.860 ;
        RECT -163.545 -78.010 -163.375 -77.860 ;
        RECT -164.485 -78.180 -163.375 -78.010 ;
        RECT -164.485 -78.385 -164.315 -78.180 ;
        RECT -173.465 -78.715 -172.535 -78.385 ;
        RECT -165.245 -78.715 -164.315 -78.385 ;
        RECT -173.465 -79.240 -173.295 -78.715 ;
        RECT -164.485 -79.240 -164.315 -78.715 ;
        RECT -164.075 -79.345 -163.785 -78.180 ;
        RECT -163.545 -78.385 -163.375 -78.180 ;
        RECT -154.565 -78.010 -154.395 -77.860 ;
        RECT -153.625 -78.010 -153.455 -77.860 ;
        RECT -154.565 -78.180 -153.455 -78.010 ;
        RECT -154.565 -78.385 -154.395 -78.180 ;
        RECT -163.545 -78.715 -162.615 -78.385 ;
        RECT -155.325 -78.715 -154.395 -78.385 ;
        RECT -163.545 -79.240 -163.375 -78.715 ;
        RECT -154.565 -79.240 -154.395 -78.715 ;
        RECT -154.155 -79.345 -153.865 -78.180 ;
        RECT -153.625 -78.385 -153.455 -78.180 ;
        RECT -144.645 -78.010 -144.475 -77.860 ;
        RECT -143.705 -78.010 -143.535 -77.860 ;
        RECT -144.645 -78.180 -143.535 -78.010 ;
        RECT -144.645 -78.385 -144.475 -78.180 ;
        RECT -153.625 -78.715 -152.695 -78.385 ;
        RECT -145.405 -78.715 -144.475 -78.385 ;
        RECT -153.625 -79.240 -153.455 -78.715 ;
        RECT -144.645 -79.240 -144.475 -78.715 ;
        RECT -144.235 -79.345 -143.945 -78.180 ;
        RECT -143.705 -78.385 -143.535 -78.180 ;
        RECT -134.725 -78.010 -134.555 -77.860 ;
        RECT -133.785 -78.010 -133.615 -77.860 ;
        RECT -134.725 -78.180 -133.615 -78.010 ;
        RECT -134.725 -78.385 -134.555 -78.180 ;
        RECT -143.705 -78.715 -142.775 -78.385 ;
        RECT -135.485 -78.715 -134.555 -78.385 ;
        RECT -143.705 -79.240 -143.535 -78.715 ;
        RECT -134.725 -79.240 -134.555 -78.715 ;
        RECT -134.315 -79.345 -134.025 -78.180 ;
        RECT -133.785 -78.385 -133.615 -78.180 ;
        RECT -124.805 -78.010 -124.635 -77.860 ;
        RECT -123.865 -78.010 -123.695 -77.860 ;
        RECT -124.805 -78.180 -123.695 -78.010 ;
        RECT -124.805 -78.385 -124.635 -78.180 ;
        RECT -133.785 -78.715 -132.855 -78.385 ;
        RECT -125.565 -78.715 -124.635 -78.385 ;
        RECT -133.785 -79.240 -133.615 -78.715 ;
        RECT -124.805 -79.240 -124.635 -78.715 ;
        RECT -124.395 -79.345 -124.105 -78.180 ;
        RECT -123.865 -78.385 -123.695 -78.180 ;
        RECT -114.885 -78.010 -114.715 -77.860 ;
        RECT -113.945 -78.010 -113.775 -77.860 ;
        RECT -114.885 -78.180 -113.775 -78.010 ;
        RECT -114.885 -78.385 -114.715 -78.180 ;
        RECT -123.865 -78.715 -122.935 -78.385 ;
        RECT -115.645 -78.715 -114.715 -78.385 ;
        RECT -123.865 -79.240 -123.695 -78.715 ;
        RECT -114.885 -79.240 -114.715 -78.715 ;
        RECT -114.475 -79.345 -114.185 -78.180 ;
        RECT -113.945 -78.385 -113.775 -78.180 ;
        RECT -104.965 -78.010 -104.795 -77.860 ;
        RECT -104.025 -78.010 -103.855 -77.860 ;
        RECT -104.965 -78.180 -103.855 -78.010 ;
        RECT -104.965 -78.385 -104.795 -78.180 ;
        RECT -113.945 -78.715 -113.015 -78.385 ;
        RECT -105.725 -78.715 -104.795 -78.385 ;
        RECT -113.945 -79.240 -113.775 -78.715 ;
        RECT -104.965 -79.240 -104.795 -78.715 ;
        RECT -104.555 -79.345 -104.265 -78.180 ;
        RECT -104.025 -78.385 -103.855 -78.180 ;
        RECT -95.045 -78.010 -94.875 -77.860 ;
        RECT -94.105 -78.010 -93.935 -77.860 ;
        RECT -95.045 -78.180 -93.935 -78.010 ;
        RECT -95.045 -78.385 -94.875 -78.180 ;
        RECT -104.025 -78.715 -103.095 -78.385 ;
        RECT -95.805 -78.715 -94.875 -78.385 ;
        RECT -104.025 -79.240 -103.855 -78.715 ;
        RECT -95.045 -79.240 -94.875 -78.715 ;
        RECT -94.635 -79.345 -94.345 -78.180 ;
        RECT -94.105 -78.385 -93.935 -78.180 ;
        RECT -85.125 -78.010 -84.955 -77.860 ;
        RECT -84.185 -78.010 -84.015 -77.860 ;
        RECT -85.125 -78.180 -84.015 -78.010 ;
        RECT -85.125 -78.385 -84.955 -78.180 ;
        RECT -94.105 -78.715 -93.175 -78.385 ;
        RECT -85.885 -78.715 -84.955 -78.385 ;
        RECT -94.105 -79.240 -93.935 -78.715 ;
        RECT -85.125 -79.240 -84.955 -78.715 ;
        RECT -84.715 -79.345 -84.425 -78.180 ;
        RECT -84.185 -78.385 -84.015 -78.180 ;
        RECT -75.205 -78.010 -75.035 -77.860 ;
        RECT -74.265 -78.010 -74.095 -77.860 ;
        RECT -75.205 -78.180 -74.095 -78.010 ;
        RECT -75.205 -78.385 -75.035 -78.180 ;
        RECT -84.185 -78.715 -83.255 -78.385 ;
        RECT -75.965 -78.715 -75.035 -78.385 ;
        RECT -84.185 -79.240 -84.015 -78.715 ;
        RECT -75.205 -79.240 -75.035 -78.715 ;
        RECT -74.795 -79.345 -74.505 -78.180 ;
        RECT -74.265 -78.385 -74.095 -78.180 ;
        RECT -65.285 -78.010 -65.115 -77.860 ;
        RECT -64.345 -78.010 -64.175 -77.860 ;
        RECT -65.285 -78.180 -64.175 -78.010 ;
        RECT -65.285 -78.385 -65.115 -78.180 ;
        RECT -74.265 -78.715 -73.335 -78.385 ;
        RECT -66.045 -78.715 -65.115 -78.385 ;
        RECT -74.265 -79.240 -74.095 -78.715 ;
        RECT -65.285 -79.240 -65.115 -78.715 ;
        RECT -64.875 -79.345 -64.585 -78.180 ;
        RECT -64.345 -78.385 -64.175 -78.180 ;
        RECT -55.365 -78.010 -55.195 -77.860 ;
        RECT -54.425 -78.010 -54.255 -77.860 ;
        RECT -55.365 -78.180 -54.255 -78.010 ;
        RECT -55.365 -78.385 -55.195 -78.180 ;
        RECT -64.345 -78.715 -63.415 -78.385 ;
        RECT -56.125 -78.715 -55.195 -78.385 ;
        RECT -64.345 -79.240 -64.175 -78.715 ;
        RECT -55.365 -79.240 -55.195 -78.715 ;
        RECT -54.955 -79.345 -54.665 -78.180 ;
        RECT -54.425 -78.385 -54.255 -78.180 ;
        RECT -45.445 -78.010 -45.275 -77.860 ;
        RECT -44.505 -78.010 -44.335 -77.860 ;
        RECT -45.445 -78.180 -44.335 -78.010 ;
        RECT -45.445 -78.385 -45.275 -78.180 ;
        RECT -54.425 -78.715 -53.495 -78.385 ;
        RECT -46.205 -78.715 -45.275 -78.385 ;
        RECT -54.425 -79.240 -54.255 -78.715 ;
        RECT -45.445 -79.240 -45.275 -78.715 ;
        RECT -45.035 -79.345 -44.745 -78.180 ;
        RECT -44.505 -78.385 -44.335 -78.180 ;
        RECT -35.525 -78.010 -35.355 -77.860 ;
        RECT -34.585 -78.010 -34.415 -77.860 ;
        RECT -35.525 -78.180 -34.415 -78.010 ;
        RECT -35.525 -78.385 -35.355 -78.180 ;
        RECT -44.505 -78.715 -43.575 -78.385 ;
        RECT -36.285 -78.715 -35.355 -78.385 ;
        RECT -44.505 -79.240 -44.335 -78.715 ;
        RECT -35.525 -79.240 -35.355 -78.715 ;
        RECT -35.115 -79.345 -34.825 -78.180 ;
        RECT -34.585 -78.385 -34.415 -78.180 ;
        RECT -25.605 -78.010 -25.435 -77.860 ;
        RECT -24.665 -78.010 -24.495 -77.860 ;
        RECT -25.605 -78.180 -24.495 -78.010 ;
        RECT -25.605 -78.385 -25.435 -78.180 ;
        RECT -34.585 -78.715 -33.655 -78.385 ;
        RECT -26.365 -78.715 -25.435 -78.385 ;
        RECT -34.585 -79.240 -34.415 -78.715 ;
        RECT -25.605 -79.240 -25.435 -78.715 ;
        RECT -25.195 -79.345 -24.905 -78.180 ;
        RECT -24.665 -78.385 -24.495 -78.180 ;
        RECT -15.685 -78.010 -15.515 -77.860 ;
        RECT -14.745 -78.010 -14.575 -77.860 ;
        RECT -15.685 -78.180 -14.575 -78.010 ;
        RECT -15.685 -78.385 -15.515 -78.180 ;
        RECT -24.665 -78.715 -23.735 -78.385 ;
        RECT -16.445 -78.715 -15.515 -78.385 ;
        RECT -24.665 -79.240 -24.495 -78.715 ;
        RECT -15.685 -79.240 -15.515 -78.715 ;
        RECT -15.275 -79.345 -14.985 -78.180 ;
        RECT -14.745 -78.385 -14.575 -78.180 ;
        RECT -5.765 -78.010 -5.595 -77.860 ;
        RECT -4.825 -78.010 -4.655 -77.860 ;
        RECT -5.765 -78.180 -4.655 -78.010 ;
        RECT -5.765 -78.385 -5.595 -78.180 ;
        RECT -14.745 -78.715 -13.815 -78.385 ;
        RECT -6.525 -78.715 -5.595 -78.385 ;
        RECT -14.745 -79.240 -14.575 -78.715 ;
        RECT -5.765 -79.240 -5.595 -78.715 ;
        RECT -5.355 -79.345 -5.065 -78.180 ;
        RECT -4.825 -78.385 -4.655 -78.180 ;
        RECT 4.155 -78.010 4.325 -77.860 ;
        RECT 5.095 -78.010 5.265 -77.860 ;
        RECT 4.155 -78.180 5.265 -78.010 ;
        RECT 4.155 -78.385 4.325 -78.180 ;
        RECT -4.825 -78.715 -3.895 -78.385 ;
        RECT 3.395 -78.715 4.325 -78.385 ;
        RECT -4.825 -79.240 -4.655 -78.715 ;
        RECT 4.155 -79.240 4.325 -78.715 ;
        RECT 4.565 -79.345 4.855 -78.180 ;
        RECT 5.095 -78.385 5.265 -78.180 ;
        RECT 14.075 -78.010 14.245 -77.860 ;
        RECT 15.015 -78.010 15.185 -77.860 ;
        RECT 14.075 -78.180 15.185 -78.010 ;
        RECT 14.075 -78.385 14.245 -78.180 ;
        RECT 5.095 -78.715 6.025 -78.385 ;
        RECT 13.315 -78.715 14.245 -78.385 ;
        RECT 5.095 -79.240 5.265 -78.715 ;
        RECT 14.075 -79.240 14.245 -78.715 ;
        RECT 14.485 -79.345 14.775 -78.180 ;
        RECT 15.015 -78.385 15.185 -78.180 ;
        RECT 23.995 -78.010 24.165 -77.860 ;
        RECT 23.995 -78.180 24.780 -78.010 ;
        RECT 23.995 -78.385 24.165 -78.180 ;
        RECT 15.015 -78.715 15.945 -78.385 ;
        RECT 23.235 -78.715 24.165 -78.385 ;
        RECT 15.015 -79.240 15.185 -78.715 ;
        RECT 23.995 -79.240 24.165 -78.715 ;
        RECT 24.405 -79.345 24.695 -78.180 ;
        RECT -289.540 -79.755 -286.320 -79.585 ;
        RECT -279.620 -79.755 -276.400 -79.585 ;
        RECT -269.700 -79.755 -266.480 -79.585 ;
        RECT -259.780 -79.755 -256.560 -79.585 ;
        RECT -249.860 -79.755 -246.640 -79.585 ;
        RECT -239.940 -79.755 -236.720 -79.585 ;
        RECT -230.020 -79.755 -226.800 -79.585 ;
        RECT -220.100 -79.755 -216.880 -79.585 ;
        RECT -210.180 -79.755 -206.960 -79.585 ;
        RECT -200.260 -79.755 -197.040 -79.585 ;
        RECT -190.340 -79.755 -187.120 -79.585 ;
        RECT -180.420 -79.755 -177.200 -79.585 ;
        RECT -170.500 -79.755 -167.280 -79.585 ;
        RECT -160.580 -79.755 -157.360 -79.585 ;
        RECT -150.660 -79.755 -147.440 -79.585 ;
        RECT -140.740 -79.755 -137.520 -79.585 ;
        RECT -130.820 -79.755 -127.600 -79.585 ;
        RECT -120.900 -79.755 -117.680 -79.585 ;
        RECT -110.980 -79.755 -107.760 -79.585 ;
        RECT -101.060 -79.755 -97.840 -79.585 ;
        RECT -91.140 -79.755 -87.920 -79.585 ;
        RECT -81.220 -79.755 -78.000 -79.585 ;
        RECT -71.300 -79.755 -68.080 -79.585 ;
        RECT -61.380 -79.755 -58.160 -79.585 ;
        RECT -51.460 -79.755 -48.240 -79.585 ;
        RECT -41.540 -79.755 -38.320 -79.585 ;
        RECT -31.620 -79.755 -28.400 -79.585 ;
        RECT -21.700 -79.755 -18.480 -79.585 ;
        RECT -11.780 -79.755 -8.560 -79.585 ;
        RECT -1.860 -79.755 1.360 -79.585 ;
        RECT 8.060 -79.755 11.280 -79.585 ;
        RECT 17.980 -79.755 21.200 -79.585 ;
        RECT -289.455 -80.895 -289.195 -79.755 ;
        RECT -288.525 -80.895 -288.245 -79.755 ;
        RECT -288.075 -80.920 -287.785 -79.755 ;
        RECT -287.615 -80.895 -287.335 -79.755 ;
        RECT -286.665 -80.895 -286.405 -79.755 ;
        RECT -279.535 -80.895 -279.275 -79.755 ;
        RECT -278.605 -80.895 -278.325 -79.755 ;
        RECT -278.155 -80.920 -277.865 -79.755 ;
        RECT -277.695 -80.895 -277.415 -79.755 ;
        RECT -276.745 -80.895 -276.485 -79.755 ;
        RECT -269.615 -80.895 -269.355 -79.755 ;
        RECT -268.685 -80.895 -268.405 -79.755 ;
        RECT -268.235 -80.920 -267.945 -79.755 ;
        RECT -267.775 -80.895 -267.495 -79.755 ;
        RECT -266.825 -80.895 -266.565 -79.755 ;
        RECT -259.695 -80.895 -259.435 -79.755 ;
        RECT -258.765 -80.895 -258.485 -79.755 ;
        RECT -258.315 -80.920 -258.025 -79.755 ;
        RECT -257.855 -80.895 -257.575 -79.755 ;
        RECT -256.905 -80.895 -256.645 -79.755 ;
        RECT -249.775 -80.895 -249.515 -79.755 ;
        RECT -248.845 -80.895 -248.565 -79.755 ;
        RECT -248.395 -80.920 -248.105 -79.755 ;
        RECT -247.935 -80.895 -247.655 -79.755 ;
        RECT -246.985 -80.895 -246.725 -79.755 ;
        RECT -239.855 -80.895 -239.595 -79.755 ;
        RECT -238.925 -80.895 -238.645 -79.755 ;
        RECT -238.475 -80.920 -238.185 -79.755 ;
        RECT -238.015 -80.895 -237.735 -79.755 ;
        RECT -237.065 -80.895 -236.805 -79.755 ;
        RECT -229.935 -80.895 -229.675 -79.755 ;
        RECT -229.005 -80.895 -228.725 -79.755 ;
        RECT -228.555 -80.920 -228.265 -79.755 ;
        RECT -228.095 -80.895 -227.815 -79.755 ;
        RECT -227.145 -80.895 -226.885 -79.755 ;
        RECT -220.015 -80.895 -219.755 -79.755 ;
        RECT -219.085 -80.895 -218.805 -79.755 ;
        RECT -218.635 -80.920 -218.345 -79.755 ;
        RECT -218.175 -80.895 -217.895 -79.755 ;
        RECT -217.225 -80.895 -216.965 -79.755 ;
        RECT -210.095 -80.895 -209.835 -79.755 ;
        RECT -209.165 -80.895 -208.885 -79.755 ;
        RECT -208.715 -80.920 -208.425 -79.755 ;
        RECT -208.255 -80.895 -207.975 -79.755 ;
        RECT -207.305 -80.895 -207.045 -79.755 ;
        RECT -200.175 -80.895 -199.915 -79.755 ;
        RECT -199.245 -80.895 -198.965 -79.755 ;
        RECT -198.795 -80.920 -198.505 -79.755 ;
        RECT -198.335 -80.895 -198.055 -79.755 ;
        RECT -197.385 -80.895 -197.125 -79.755 ;
        RECT -190.255 -80.895 -189.995 -79.755 ;
        RECT -189.325 -80.895 -189.045 -79.755 ;
        RECT -188.875 -80.920 -188.585 -79.755 ;
        RECT -188.415 -80.895 -188.135 -79.755 ;
        RECT -187.465 -80.895 -187.205 -79.755 ;
        RECT -180.335 -80.895 -180.075 -79.755 ;
        RECT -179.405 -80.895 -179.125 -79.755 ;
        RECT -178.955 -80.920 -178.665 -79.755 ;
        RECT -178.495 -80.895 -178.215 -79.755 ;
        RECT -177.545 -80.895 -177.285 -79.755 ;
        RECT -170.415 -80.895 -170.155 -79.755 ;
        RECT -169.485 -80.895 -169.205 -79.755 ;
        RECT -169.035 -80.920 -168.745 -79.755 ;
        RECT -168.575 -80.895 -168.295 -79.755 ;
        RECT -167.625 -80.895 -167.365 -79.755 ;
        RECT -160.495 -80.895 -160.235 -79.755 ;
        RECT -159.565 -80.895 -159.285 -79.755 ;
        RECT -159.115 -80.920 -158.825 -79.755 ;
        RECT -158.655 -80.895 -158.375 -79.755 ;
        RECT -157.705 -80.895 -157.445 -79.755 ;
        RECT -150.575 -80.895 -150.315 -79.755 ;
        RECT -149.645 -80.895 -149.365 -79.755 ;
        RECT -149.195 -80.920 -148.905 -79.755 ;
        RECT -148.735 -80.895 -148.455 -79.755 ;
        RECT -147.785 -80.895 -147.525 -79.755 ;
        RECT -140.655 -80.895 -140.395 -79.755 ;
        RECT -139.725 -80.895 -139.445 -79.755 ;
        RECT -139.275 -80.920 -138.985 -79.755 ;
        RECT -138.815 -80.895 -138.535 -79.755 ;
        RECT -137.865 -80.895 -137.605 -79.755 ;
        RECT -130.735 -80.895 -130.475 -79.755 ;
        RECT -129.805 -80.895 -129.525 -79.755 ;
        RECT -129.355 -80.920 -129.065 -79.755 ;
        RECT -128.895 -80.895 -128.615 -79.755 ;
        RECT -127.945 -80.895 -127.685 -79.755 ;
        RECT -120.815 -80.895 -120.555 -79.755 ;
        RECT -119.885 -80.895 -119.605 -79.755 ;
        RECT -119.435 -80.920 -119.145 -79.755 ;
        RECT -118.975 -80.895 -118.695 -79.755 ;
        RECT -118.025 -80.895 -117.765 -79.755 ;
        RECT -110.895 -80.895 -110.635 -79.755 ;
        RECT -109.965 -80.895 -109.685 -79.755 ;
        RECT -109.515 -80.920 -109.225 -79.755 ;
        RECT -109.055 -80.895 -108.775 -79.755 ;
        RECT -108.105 -80.895 -107.845 -79.755 ;
        RECT -100.975 -80.895 -100.715 -79.755 ;
        RECT -100.045 -80.895 -99.765 -79.755 ;
        RECT -99.595 -80.920 -99.305 -79.755 ;
        RECT -99.135 -80.895 -98.855 -79.755 ;
        RECT -98.185 -80.895 -97.925 -79.755 ;
        RECT -91.055 -80.895 -90.795 -79.755 ;
        RECT -90.125 -80.895 -89.845 -79.755 ;
        RECT -89.675 -80.920 -89.385 -79.755 ;
        RECT -89.215 -80.895 -88.935 -79.755 ;
        RECT -88.265 -80.895 -88.005 -79.755 ;
        RECT -81.135 -80.895 -80.875 -79.755 ;
        RECT -80.205 -80.895 -79.925 -79.755 ;
        RECT -79.755 -80.920 -79.465 -79.755 ;
        RECT -79.295 -80.895 -79.015 -79.755 ;
        RECT -78.345 -80.895 -78.085 -79.755 ;
        RECT -71.215 -80.895 -70.955 -79.755 ;
        RECT -70.285 -80.895 -70.005 -79.755 ;
        RECT -69.835 -80.920 -69.545 -79.755 ;
        RECT -69.375 -80.895 -69.095 -79.755 ;
        RECT -68.425 -80.895 -68.165 -79.755 ;
        RECT -61.295 -80.895 -61.035 -79.755 ;
        RECT -60.365 -80.895 -60.085 -79.755 ;
        RECT -59.915 -80.920 -59.625 -79.755 ;
        RECT -59.455 -80.895 -59.175 -79.755 ;
        RECT -58.505 -80.895 -58.245 -79.755 ;
        RECT -51.375 -80.895 -51.115 -79.755 ;
        RECT -50.445 -80.895 -50.165 -79.755 ;
        RECT -49.995 -80.920 -49.705 -79.755 ;
        RECT -49.535 -80.895 -49.255 -79.755 ;
        RECT -48.585 -80.895 -48.325 -79.755 ;
        RECT -41.455 -80.895 -41.195 -79.755 ;
        RECT -40.525 -80.895 -40.245 -79.755 ;
        RECT -40.075 -80.920 -39.785 -79.755 ;
        RECT -39.615 -80.895 -39.335 -79.755 ;
        RECT -38.665 -80.895 -38.405 -79.755 ;
        RECT -31.535 -80.895 -31.275 -79.755 ;
        RECT -30.605 -80.895 -30.325 -79.755 ;
        RECT -30.155 -80.920 -29.865 -79.755 ;
        RECT -29.695 -80.895 -29.415 -79.755 ;
        RECT -28.745 -80.895 -28.485 -79.755 ;
        RECT -21.615 -80.895 -21.355 -79.755 ;
        RECT -20.685 -80.895 -20.405 -79.755 ;
        RECT -20.235 -80.920 -19.945 -79.755 ;
        RECT -19.775 -80.895 -19.495 -79.755 ;
        RECT -18.825 -80.895 -18.565 -79.755 ;
        RECT -11.695 -80.895 -11.435 -79.755 ;
        RECT -10.765 -80.895 -10.485 -79.755 ;
        RECT -10.315 -80.920 -10.025 -79.755 ;
        RECT -9.855 -80.895 -9.575 -79.755 ;
        RECT -8.905 -80.895 -8.645 -79.755 ;
        RECT -1.775 -80.895 -1.515 -79.755 ;
        RECT -0.845 -80.895 -0.565 -79.755 ;
        RECT -0.395 -80.920 -0.105 -79.755 ;
        RECT 0.065 -80.895 0.345 -79.755 ;
        RECT 1.015 -80.895 1.275 -79.755 ;
        RECT 8.145 -80.895 8.405 -79.755 ;
        RECT 9.075 -80.895 9.355 -79.755 ;
        RECT 9.525 -80.920 9.815 -79.755 ;
        RECT 9.985 -80.895 10.265 -79.755 ;
        RECT 10.935 -80.895 11.195 -79.755 ;
        RECT 18.065 -80.895 18.325 -79.755 ;
        RECT 18.995 -80.895 19.275 -79.755 ;
        RECT 19.445 -80.920 19.735 -79.755 ;
        RECT 19.905 -80.895 20.185 -79.755 ;
        RECT 20.855 -80.895 21.115 -79.755 ;
        RECT -284.495 -82.305 -284.235 -81.165 ;
        RECT -283.565 -82.305 -283.285 -81.165 ;
        RECT -283.115 -82.305 -282.825 -81.140 ;
        RECT -282.655 -82.305 -282.375 -81.165 ;
        RECT -281.705 -82.305 -281.445 -81.165 ;
        RECT -274.575 -82.305 -274.315 -81.165 ;
        RECT -273.645 -82.305 -273.365 -81.165 ;
        RECT -273.195 -82.305 -272.905 -81.140 ;
        RECT -272.735 -82.305 -272.455 -81.165 ;
        RECT -271.785 -82.305 -271.525 -81.165 ;
        RECT -264.655 -82.305 -264.395 -81.165 ;
        RECT -263.725 -82.305 -263.445 -81.165 ;
        RECT -263.275 -82.305 -262.985 -81.140 ;
        RECT -262.815 -82.305 -262.535 -81.165 ;
        RECT -261.865 -82.305 -261.605 -81.165 ;
        RECT -254.735 -82.305 -254.475 -81.165 ;
        RECT -253.805 -82.305 -253.525 -81.165 ;
        RECT -253.355 -82.305 -253.065 -81.140 ;
        RECT -252.895 -82.305 -252.615 -81.165 ;
        RECT -251.945 -82.305 -251.685 -81.165 ;
        RECT -244.815 -82.305 -244.555 -81.165 ;
        RECT -243.885 -82.305 -243.605 -81.165 ;
        RECT -243.435 -82.305 -243.145 -81.140 ;
        RECT -242.975 -82.305 -242.695 -81.165 ;
        RECT -242.025 -82.305 -241.765 -81.165 ;
        RECT -234.895 -82.305 -234.635 -81.165 ;
        RECT -233.965 -82.305 -233.685 -81.165 ;
        RECT -233.515 -82.305 -233.225 -81.140 ;
        RECT -233.055 -82.305 -232.775 -81.165 ;
        RECT -232.105 -82.305 -231.845 -81.165 ;
        RECT -224.975 -82.305 -224.715 -81.165 ;
        RECT -224.045 -82.305 -223.765 -81.165 ;
        RECT -223.595 -82.305 -223.305 -81.140 ;
        RECT -223.135 -82.305 -222.855 -81.165 ;
        RECT -222.185 -82.305 -221.925 -81.165 ;
        RECT -215.055 -82.305 -214.795 -81.165 ;
        RECT -214.125 -82.305 -213.845 -81.165 ;
        RECT -213.675 -82.305 -213.385 -81.140 ;
        RECT -213.215 -82.305 -212.935 -81.165 ;
        RECT -212.265 -82.305 -212.005 -81.165 ;
        RECT -205.135 -82.305 -204.875 -81.165 ;
        RECT -204.205 -82.305 -203.925 -81.165 ;
        RECT -203.755 -82.305 -203.465 -81.140 ;
        RECT -203.295 -82.305 -203.015 -81.165 ;
        RECT -202.345 -82.305 -202.085 -81.165 ;
        RECT -195.215 -82.305 -194.955 -81.165 ;
        RECT -194.285 -82.305 -194.005 -81.165 ;
        RECT -193.835 -82.305 -193.545 -81.140 ;
        RECT -193.375 -82.305 -193.095 -81.165 ;
        RECT -192.425 -82.305 -192.165 -81.165 ;
        RECT -185.295 -82.305 -185.035 -81.165 ;
        RECT -184.365 -82.305 -184.085 -81.165 ;
        RECT -183.915 -82.305 -183.625 -81.140 ;
        RECT -183.455 -82.305 -183.175 -81.165 ;
        RECT -182.505 -82.305 -182.245 -81.165 ;
        RECT -175.375 -82.305 -175.115 -81.165 ;
        RECT -174.445 -82.305 -174.165 -81.165 ;
        RECT -173.995 -82.305 -173.705 -81.140 ;
        RECT -173.535 -82.305 -173.255 -81.165 ;
        RECT -172.585 -82.305 -172.325 -81.165 ;
        RECT -165.455 -82.305 -165.195 -81.165 ;
        RECT -164.525 -82.305 -164.245 -81.165 ;
        RECT -164.075 -82.305 -163.785 -81.140 ;
        RECT -163.615 -82.305 -163.335 -81.165 ;
        RECT -162.665 -82.305 -162.405 -81.165 ;
        RECT -155.535 -82.305 -155.275 -81.165 ;
        RECT -154.605 -82.305 -154.325 -81.165 ;
        RECT -154.155 -82.305 -153.865 -81.140 ;
        RECT -153.695 -82.305 -153.415 -81.165 ;
        RECT -152.745 -82.305 -152.485 -81.165 ;
        RECT -145.615 -82.305 -145.355 -81.165 ;
        RECT -144.685 -82.305 -144.405 -81.165 ;
        RECT -144.235 -82.305 -143.945 -81.140 ;
        RECT -143.775 -82.305 -143.495 -81.165 ;
        RECT -142.825 -82.305 -142.565 -81.165 ;
        RECT -135.695 -82.305 -135.435 -81.165 ;
        RECT -134.765 -82.305 -134.485 -81.165 ;
        RECT -134.315 -82.305 -134.025 -81.140 ;
        RECT -133.855 -82.305 -133.575 -81.165 ;
        RECT -132.905 -82.305 -132.645 -81.165 ;
        RECT -125.775 -82.305 -125.515 -81.165 ;
        RECT -124.845 -82.305 -124.565 -81.165 ;
        RECT -124.395 -82.305 -124.105 -81.140 ;
        RECT -123.935 -82.305 -123.655 -81.165 ;
        RECT -122.985 -82.305 -122.725 -81.165 ;
        RECT -115.855 -82.305 -115.595 -81.165 ;
        RECT -114.925 -82.305 -114.645 -81.165 ;
        RECT -114.475 -82.305 -114.185 -81.140 ;
        RECT -114.015 -82.305 -113.735 -81.165 ;
        RECT -113.065 -82.305 -112.805 -81.165 ;
        RECT -105.935 -82.305 -105.675 -81.165 ;
        RECT -105.005 -82.305 -104.725 -81.165 ;
        RECT -104.555 -82.305 -104.265 -81.140 ;
        RECT -104.095 -82.305 -103.815 -81.165 ;
        RECT -103.145 -82.305 -102.885 -81.165 ;
        RECT -96.015 -82.305 -95.755 -81.165 ;
        RECT -95.085 -82.305 -94.805 -81.165 ;
        RECT -94.635 -82.305 -94.345 -81.140 ;
        RECT -94.175 -82.305 -93.895 -81.165 ;
        RECT -93.225 -82.305 -92.965 -81.165 ;
        RECT -86.095 -82.305 -85.835 -81.165 ;
        RECT -85.165 -82.305 -84.885 -81.165 ;
        RECT -84.715 -82.305 -84.425 -81.140 ;
        RECT -84.255 -82.305 -83.975 -81.165 ;
        RECT -83.305 -82.305 -83.045 -81.165 ;
        RECT -76.175 -82.305 -75.915 -81.165 ;
        RECT -75.245 -82.305 -74.965 -81.165 ;
        RECT -74.795 -82.305 -74.505 -81.140 ;
        RECT -74.335 -82.305 -74.055 -81.165 ;
        RECT -73.385 -82.305 -73.125 -81.165 ;
        RECT -66.255 -82.305 -65.995 -81.165 ;
        RECT -65.325 -82.305 -65.045 -81.165 ;
        RECT -64.875 -82.305 -64.585 -81.140 ;
        RECT -64.415 -82.305 -64.135 -81.165 ;
        RECT -63.465 -82.305 -63.205 -81.165 ;
        RECT -56.335 -82.305 -56.075 -81.165 ;
        RECT -55.405 -82.305 -55.125 -81.165 ;
        RECT -54.955 -82.305 -54.665 -81.140 ;
        RECT -54.495 -82.305 -54.215 -81.165 ;
        RECT -53.545 -82.305 -53.285 -81.165 ;
        RECT -46.415 -82.305 -46.155 -81.165 ;
        RECT -45.485 -82.305 -45.205 -81.165 ;
        RECT -45.035 -82.305 -44.745 -81.140 ;
        RECT -44.575 -82.305 -44.295 -81.165 ;
        RECT -43.625 -82.305 -43.365 -81.165 ;
        RECT -36.495 -82.305 -36.235 -81.165 ;
        RECT -35.565 -82.305 -35.285 -81.165 ;
        RECT -35.115 -82.305 -34.825 -81.140 ;
        RECT -34.655 -82.305 -34.375 -81.165 ;
        RECT -33.705 -82.305 -33.445 -81.165 ;
        RECT -26.575 -82.305 -26.315 -81.165 ;
        RECT -25.645 -82.305 -25.365 -81.165 ;
        RECT -25.195 -82.305 -24.905 -81.140 ;
        RECT -24.735 -82.305 -24.455 -81.165 ;
        RECT -23.785 -82.305 -23.525 -81.165 ;
        RECT -16.655 -82.305 -16.395 -81.165 ;
        RECT -15.725 -82.305 -15.445 -81.165 ;
        RECT -15.275 -82.305 -14.985 -81.140 ;
        RECT -14.815 -82.305 -14.535 -81.165 ;
        RECT -13.865 -82.305 -13.605 -81.165 ;
        RECT -6.735 -82.305 -6.475 -81.165 ;
        RECT -5.805 -82.305 -5.525 -81.165 ;
        RECT -5.355 -82.305 -5.065 -81.140 ;
        RECT -4.895 -82.305 -4.615 -81.165 ;
        RECT -3.945 -82.305 -3.685 -81.165 ;
        RECT 3.185 -82.305 3.445 -81.165 ;
        RECT 4.115 -82.305 4.395 -81.165 ;
        RECT 4.565 -82.305 4.855 -81.140 ;
        RECT 5.025 -82.305 5.305 -81.165 ;
        RECT 5.975 -82.305 6.235 -81.165 ;
        RECT 13.105 -82.305 13.365 -81.165 ;
        RECT 14.035 -82.305 14.315 -81.165 ;
        RECT 14.485 -82.305 14.775 -81.140 ;
        RECT 14.945 -82.305 15.225 -81.165 ;
        RECT 15.895 -82.305 16.155 -81.165 ;
        RECT 23.025 -82.305 23.285 -81.165 ;
        RECT 23.955 -82.305 24.235 -81.165 ;
        RECT 24.405 -82.305 24.695 -81.140 ;
        RECT -284.580 -82.475 -281.360 -82.305 ;
        RECT -274.660 -82.475 -271.440 -82.305 ;
        RECT -264.740 -82.475 -261.520 -82.305 ;
        RECT -254.820 -82.475 -251.600 -82.305 ;
        RECT -244.900 -82.475 -241.680 -82.305 ;
        RECT -234.980 -82.475 -231.760 -82.305 ;
        RECT -225.060 -82.475 -221.840 -82.305 ;
        RECT -215.140 -82.475 -211.920 -82.305 ;
        RECT -205.220 -82.475 -202.000 -82.305 ;
        RECT -195.300 -82.475 -192.080 -82.305 ;
        RECT -185.380 -82.475 -182.160 -82.305 ;
        RECT -175.460 -82.475 -172.240 -82.305 ;
        RECT -165.540 -82.475 -162.320 -82.305 ;
        RECT -155.620 -82.475 -152.400 -82.305 ;
        RECT -145.700 -82.475 -142.480 -82.305 ;
        RECT -135.780 -82.475 -132.560 -82.305 ;
        RECT -125.860 -82.475 -122.640 -82.305 ;
        RECT -115.940 -82.475 -112.720 -82.305 ;
        RECT -106.020 -82.475 -102.800 -82.305 ;
        RECT -96.100 -82.475 -92.880 -82.305 ;
        RECT -86.180 -82.475 -82.960 -82.305 ;
        RECT -76.260 -82.475 -73.040 -82.305 ;
        RECT -66.340 -82.475 -63.120 -82.305 ;
        RECT -56.420 -82.475 -53.200 -82.305 ;
        RECT -46.500 -82.475 -43.280 -82.305 ;
        RECT -36.580 -82.475 -33.360 -82.305 ;
        RECT -26.660 -82.475 -23.440 -82.305 ;
        RECT -16.740 -82.475 -13.520 -82.305 ;
        RECT -6.820 -82.475 -3.600 -82.305 ;
        RECT 3.100 -82.475 6.320 -82.305 ;
        RECT 13.020 -82.475 16.240 -82.305 ;
        RECT 22.940 -82.475 24.780 -82.305 ;
        RECT -288.485 -82.890 -288.315 -82.820 ;
        RECT -287.545 -82.890 -287.375 -82.820 ;
        RECT -288.485 -83.060 -287.375 -82.890 ;
        RECT -288.485 -83.345 -288.315 -83.060 ;
        RECT -289.245 -83.675 -288.315 -83.345 ;
        RECT -288.485 -84.200 -288.315 -83.675 ;
        RECT -288.075 -84.225 -287.785 -83.060 ;
        RECT -287.545 -83.345 -287.375 -83.060 ;
        RECT -278.565 -82.890 -278.395 -82.820 ;
        RECT -277.625 -82.890 -277.455 -82.820 ;
        RECT -278.565 -83.060 -277.455 -82.890 ;
        RECT -278.565 -83.345 -278.395 -83.060 ;
        RECT -287.545 -83.675 -286.615 -83.345 ;
        RECT -279.325 -83.675 -278.395 -83.345 ;
        RECT -287.545 -84.200 -287.375 -83.675 ;
        RECT -278.565 -84.200 -278.395 -83.675 ;
        RECT -278.155 -84.225 -277.865 -83.060 ;
        RECT -277.625 -83.345 -277.455 -83.060 ;
        RECT -268.645 -82.890 -268.475 -82.820 ;
        RECT -267.705 -82.890 -267.535 -82.820 ;
        RECT -268.645 -83.060 -267.535 -82.890 ;
        RECT -268.645 -83.345 -268.475 -83.060 ;
        RECT -277.625 -83.675 -276.695 -83.345 ;
        RECT -269.405 -83.675 -268.475 -83.345 ;
        RECT -277.625 -84.200 -277.455 -83.675 ;
        RECT -268.645 -84.200 -268.475 -83.675 ;
        RECT -268.235 -84.225 -267.945 -83.060 ;
        RECT -267.705 -83.345 -267.535 -83.060 ;
        RECT -258.725 -82.890 -258.555 -82.820 ;
        RECT -257.785 -82.890 -257.615 -82.820 ;
        RECT -258.725 -83.060 -257.615 -82.890 ;
        RECT -258.725 -83.345 -258.555 -83.060 ;
        RECT -267.705 -83.675 -266.775 -83.345 ;
        RECT -259.485 -83.675 -258.555 -83.345 ;
        RECT -267.705 -84.200 -267.535 -83.675 ;
        RECT -258.725 -84.200 -258.555 -83.675 ;
        RECT -258.315 -84.225 -258.025 -83.060 ;
        RECT -257.785 -83.345 -257.615 -83.060 ;
        RECT -248.805 -82.890 -248.635 -82.820 ;
        RECT -247.865 -82.890 -247.695 -82.820 ;
        RECT -248.805 -83.060 -247.695 -82.890 ;
        RECT -248.805 -83.345 -248.635 -83.060 ;
        RECT -257.785 -83.675 -256.855 -83.345 ;
        RECT -249.565 -83.675 -248.635 -83.345 ;
        RECT -257.785 -84.200 -257.615 -83.675 ;
        RECT -248.805 -84.200 -248.635 -83.675 ;
        RECT -248.395 -84.225 -248.105 -83.060 ;
        RECT -247.865 -83.345 -247.695 -83.060 ;
        RECT -238.885 -82.890 -238.715 -82.820 ;
        RECT -237.945 -82.890 -237.775 -82.820 ;
        RECT -238.885 -83.060 -237.775 -82.890 ;
        RECT -238.885 -83.345 -238.715 -83.060 ;
        RECT -247.865 -83.675 -246.935 -83.345 ;
        RECT -239.645 -83.675 -238.715 -83.345 ;
        RECT -247.865 -84.200 -247.695 -83.675 ;
        RECT -238.885 -84.200 -238.715 -83.675 ;
        RECT -238.475 -84.225 -238.185 -83.060 ;
        RECT -237.945 -83.345 -237.775 -83.060 ;
        RECT -228.965 -82.890 -228.795 -82.820 ;
        RECT -228.025 -82.890 -227.855 -82.820 ;
        RECT -228.965 -83.060 -227.855 -82.890 ;
        RECT -228.965 -83.345 -228.795 -83.060 ;
        RECT -237.945 -83.675 -237.015 -83.345 ;
        RECT -229.725 -83.675 -228.795 -83.345 ;
        RECT -237.945 -84.200 -237.775 -83.675 ;
        RECT -228.965 -84.200 -228.795 -83.675 ;
        RECT -228.555 -84.225 -228.265 -83.060 ;
        RECT -228.025 -83.345 -227.855 -83.060 ;
        RECT -219.045 -82.890 -218.875 -82.820 ;
        RECT -218.105 -82.890 -217.935 -82.820 ;
        RECT -219.045 -83.060 -217.935 -82.890 ;
        RECT -219.045 -83.345 -218.875 -83.060 ;
        RECT -228.025 -83.675 -227.095 -83.345 ;
        RECT -219.805 -83.675 -218.875 -83.345 ;
        RECT -228.025 -84.200 -227.855 -83.675 ;
        RECT -219.045 -84.200 -218.875 -83.675 ;
        RECT -218.635 -84.225 -218.345 -83.060 ;
        RECT -218.105 -83.345 -217.935 -83.060 ;
        RECT -209.125 -82.890 -208.955 -82.820 ;
        RECT -208.185 -82.890 -208.015 -82.820 ;
        RECT -209.125 -83.060 -208.015 -82.890 ;
        RECT -209.125 -83.345 -208.955 -83.060 ;
        RECT -218.105 -83.675 -217.175 -83.345 ;
        RECT -209.885 -83.675 -208.955 -83.345 ;
        RECT -218.105 -84.200 -217.935 -83.675 ;
        RECT -209.125 -84.200 -208.955 -83.675 ;
        RECT -208.715 -84.225 -208.425 -83.060 ;
        RECT -208.185 -83.345 -208.015 -83.060 ;
        RECT -199.205 -82.890 -199.035 -82.820 ;
        RECT -198.265 -82.890 -198.095 -82.820 ;
        RECT -199.205 -83.060 -198.095 -82.890 ;
        RECT -199.205 -83.345 -199.035 -83.060 ;
        RECT -208.185 -83.675 -207.255 -83.345 ;
        RECT -199.965 -83.675 -199.035 -83.345 ;
        RECT -208.185 -84.200 -208.015 -83.675 ;
        RECT -199.205 -84.200 -199.035 -83.675 ;
        RECT -198.795 -84.225 -198.505 -83.060 ;
        RECT -198.265 -83.345 -198.095 -83.060 ;
        RECT -189.285 -82.890 -189.115 -82.820 ;
        RECT -188.345 -82.890 -188.175 -82.820 ;
        RECT -189.285 -83.060 -188.175 -82.890 ;
        RECT -189.285 -83.345 -189.115 -83.060 ;
        RECT -198.265 -83.675 -197.335 -83.345 ;
        RECT -190.045 -83.675 -189.115 -83.345 ;
        RECT -198.265 -84.200 -198.095 -83.675 ;
        RECT -189.285 -84.200 -189.115 -83.675 ;
        RECT -188.875 -84.225 -188.585 -83.060 ;
        RECT -188.345 -83.345 -188.175 -83.060 ;
        RECT -179.365 -82.890 -179.195 -82.820 ;
        RECT -178.425 -82.890 -178.255 -82.820 ;
        RECT -179.365 -83.060 -178.255 -82.890 ;
        RECT -179.365 -83.345 -179.195 -83.060 ;
        RECT -188.345 -83.675 -187.415 -83.345 ;
        RECT -180.125 -83.675 -179.195 -83.345 ;
        RECT -188.345 -84.200 -188.175 -83.675 ;
        RECT -179.365 -84.200 -179.195 -83.675 ;
        RECT -178.955 -84.225 -178.665 -83.060 ;
        RECT -178.425 -83.345 -178.255 -83.060 ;
        RECT -169.445 -82.890 -169.275 -82.820 ;
        RECT -168.505 -82.890 -168.335 -82.820 ;
        RECT -169.445 -83.060 -168.335 -82.890 ;
        RECT -169.445 -83.345 -169.275 -83.060 ;
        RECT -178.425 -83.675 -177.495 -83.345 ;
        RECT -170.205 -83.675 -169.275 -83.345 ;
        RECT -178.425 -84.200 -178.255 -83.675 ;
        RECT -169.445 -84.200 -169.275 -83.675 ;
        RECT -169.035 -84.225 -168.745 -83.060 ;
        RECT -168.505 -83.345 -168.335 -83.060 ;
        RECT -159.525 -82.890 -159.355 -82.820 ;
        RECT -158.585 -82.890 -158.415 -82.820 ;
        RECT -159.525 -83.060 -158.415 -82.890 ;
        RECT -159.525 -83.345 -159.355 -83.060 ;
        RECT -168.505 -83.675 -167.575 -83.345 ;
        RECT -160.285 -83.675 -159.355 -83.345 ;
        RECT -168.505 -84.200 -168.335 -83.675 ;
        RECT -159.525 -84.200 -159.355 -83.675 ;
        RECT -159.115 -84.225 -158.825 -83.060 ;
        RECT -158.585 -83.345 -158.415 -83.060 ;
        RECT -149.605 -82.890 -149.435 -82.820 ;
        RECT -148.665 -82.890 -148.495 -82.820 ;
        RECT -149.605 -83.060 -148.495 -82.890 ;
        RECT -149.605 -83.345 -149.435 -83.060 ;
        RECT -158.585 -83.675 -157.655 -83.345 ;
        RECT -150.365 -83.675 -149.435 -83.345 ;
        RECT -158.585 -84.200 -158.415 -83.675 ;
        RECT -149.605 -84.200 -149.435 -83.675 ;
        RECT -149.195 -84.225 -148.905 -83.060 ;
        RECT -148.665 -83.345 -148.495 -83.060 ;
        RECT -139.685 -82.890 -139.515 -82.820 ;
        RECT -138.745 -82.890 -138.575 -82.820 ;
        RECT -139.685 -83.060 -138.575 -82.890 ;
        RECT -139.685 -83.345 -139.515 -83.060 ;
        RECT -148.665 -83.675 -147.735 -83.345 ;
        RECT -140.445 -83.675 -139.515 -83.345 ;
        RECT -148.665 -84.200 -148.495 -83.675 ;
        RECT -139.685 -84.200 -139.515 -83.675 ;
        RECT -139.275 -84.225 -138.985 -83.060 ;
        RECT -138.745 -83.345 -138.575 -83.060 ;
        RECT -129.765 -82.890 -129.595 -82.820 ;
        RECT -128.825 -82.890 -128.655 -82.820 ;
        RECT -129.765 -83.060 -128.655 -82.890 ;
        RECT -129.765 -83.345 -129.595 -83.060 ;
        RECT -138.745 -83.675 -137.815 -83.345 ;
        RECT -130.525 -83.675 -129.595 -83.345 ;
        RECT -138.745 -84.200 -138.575 -83.675 ;
        RECT -129.765 -84.200 -129.595 -83.675 ;
        RECT -129.355 -84.225 -129.065 -83.060 ;
        RECT -128.825 -83.345 -128.655 -83.060 ;
        RECT -119.845 -82.890 -119.675 -82.820 ;
        RECT -118.905 -82.890 -118.735 -82.820 ;
        RECT -119.845 -83.060 -118.735 -82.890 ;
        RECT -119.845 -83.345 -119.675 -83.060 ;
        RECT -128.825 -83.675 -127.895 -83.345 ;
        RECT -120.605 -83.675 -119.675 -83.345 ;
        RECT -128.825 -84.200 -128.655 -83.675 ;
        RECT -119.845 -84.200 -119.675 -83.675 ;
        RECT -119.435 -84.225 -119.145 -83.060 ;
        RECT -118.905 -83.345 -118.735 -83.060 ;
        RECT -109.925 -82.890 -109.755 -82.820 ;
        RECT -108.985 -82.890 -108.815 -82.820 ;
        RECT -109.925 -83.060 -108.815 -82.890 ;
        RECT -109.925 -83.345 -109.755 -83.060 ;
        RECT -118.905 -83.675 -117.975 -83.345 ;
        RECT -110.685 -83.675 -109.755 -83.345 ;
        RECT -118.905 -84.200 -118.735 -83.675 ;
        RECT -109.925 -84.200 -109.755 -83.675 ;
        RECT -109.515 -84.225 -109.225 -83.060 ;
        RECT -108.985 -83.345 -108.815 -83.060 ;
        RECT -100.005 -82.890 -99.835 -82.820 ;
        RECT -99.065 -82.890 -98.895 -82.820 ;
        RECT -100.005 -83.060 -98.895 -82.890 ;
        RECT -100.005 -83.345 -99.835 -83.060 ;
        RECT -108.985 -83.675 -108.055 -83.345 ;
        RECT -100.765 -83.675 -99.835 -83.345 ;
        RECT -108.985 -84.200 -108.815 -83.675 ;
        RECT -100.005 -84.200 -99.835 -83.675 ;
        RECT -99.595 -84.225 -99.305 -83.060 ;
        RECT -99.065 -83.345 -98.895 -83.060 ;
        RECT -90.085 -82.890 -89.915 -82.820 ;
        RECT -89.145 -82.890 -88.975 -82.820 ;
        RECT -90.085 -83.060 -88.975 -82.890 ;
        RECT -90.085 -83.345 -89.915 -83.060 ;
        RECT -99.065 -83.675 -98.135 -83.345 ;
        RECT -90.845 -83.675 -89.915 -83.345 ;
        RECT -99.065 -84.200 -98.895 -83.675 ;
        RECT -90.085 -84.200 -89.915 -83.675 ;
        RECT -89.675 -84.225 -89.385 -83.060 ;
        RECT -89.145 -83.345 -88.975 -83.060 ;
        RECT -80.165 -82.890 -79.995 -82.820 ;
        RECT -79.225 -82.890 -79.055 -82.820 ;
        RECT -80.165 -83.060 -79.055 -82.890 ;
        RECT -80.165 -83.345 -79.995 -83.060 ;
        RECT -89.145 -83.675 -88.215 -83.345 ;
        RECT -80.925 -83.675 -79.995 -83.345 ;
        RECT -89.145 -84.200 -88.975 -83.675 ;
        RECT -80.165 -84.200 -79.995 -83.675 ;
        RECT -79.755 -84.225 -79.465 -83.060 ;
        RECT -79.225 -83.345 -79.055 -83.060 ;
        RECT -70.245 -82.890 -70.075 -82.820 ;
        RECT -69.305 -82.890 -69.135 -82.820 ;
        RECT -70.245 -83.060 -69.135 -82.890 ;
        RECT -70.245 -83.345 -70.075 -83.060 ;
        RECT -79.225 -83.675 -78.295 -83.345 ;
        RECT -71.005 -83.675 -70.075 -83.345 ;
        RECT -79.225 -84.200 -79.055 -83.675 ;
        RECT -70.245 -84.200 -70.075 -83.675 ;
        RECT -69.835 -84.225 -69.545 -83.060 ;
        RECT -69.305 -83.345 -69.135 -83.060 ;
        RECT -60.325 -82.890 -60.155 -82.820 ;
        RECT -59.385 -82.890 -59.215 -82.820 ;
        RECT -60.325 -83.060 -59.215 -82.890 ;
        RECT -60.325 -83.345 -60.155 -83.060 ;
        RECT -69.305 -83.675 -68.375 -83.345 ;
        RECT -61.085 -83.675 -60.155 -83.345 ;
        RECT -69.305 -84.200 -69.135 -83.675 ;
        RECT -60.325 -84.200 -60.155 -83.675 ;
        RECT -59.915 -84.225 -59.625 -83.060 ;
        RECT -59.385 -83.345 -59.215 -83.060 ;
        RECT -50.405 -82.890 -50.235 -82.820 ;
        RECT -49.465 -82.890 -49.295 -82.820 ;
        RECT -50.405 -83.060 -49.295 -82.890 ;
        RECT -50.405 -83.345 -50.235 -83.060 ;
        RECT -59.385 -83.675 -58.455 -83.345 ;
        RECT -51.165 -83.675 -50.235 -83.345 ;
        RECT -59.385 -84.200 -59.215 -83.675 ;
        RECT -50.405 -84.200 -50.235 -83.675 ;
        RECT -49.995 -84.225 -49.705 -83.060 ;
        RECT -49.465 -83.345 -49.295 -83.060 ;
        RECT -40.485 -82.890 -40.315 -82.820 ;
        RECT -39.545 -82.890 -39.375 -82.820 ;
        RECT -40.485 -83.060 -39.375 -82.890 ;
        RECT -40.485 -83.345 -40.315 -83.060 ;
        RECT -49.465 -83.675 -48.535 -83.345 ;
        RECT -41.245 -83.675 -40.315 -83.345 ;
        RECT -49.465 -84.200 -49.295 -83.675 ;
        RECT -40.485 -84.200 -40.315 -83.675 ;
        RECT -40.075 -84.225 -39.785 -83.060 ;
        RECT -39.545 -83.345 -39.375 -83.060 ;
        RECT -30.565 -82.890 -30.395 -82.820 ;
        RECT -29.625 -82.890 -29.455 -82.820 ;
        RECT -30.565 -83.060 -29.455 -82.890 ;
        RECT -30.565 -83.345 -30.395 -83.060 ;
        RECT -39.545 -83.675 -38.615 -83.345 ;
        RECT -31.325 -83.675 -30.395 -83.345 ;
        RECT -39.545 -84.200 -39.375 -83.675 ;
        RECT -30.565 -84.200 -30.395 -83.675 ;
        RECT -30.155 -84.225 -29.865 -83.060 ;
        RECT -29.625 -83.345 -29.455 -83.060 ;
        RECT -20.645 -82.890 -20.475 -82.820 ;
        RECT -19.705 -82.890 -19.535 -82.820 ;
        RECT -20.645 -83.060 -19.535 -82.890 ;
        RECT -20.645 -83.345 -20.475 -83.060 ;
        RECT -29.625 -83.675 -28.695 -83.345 ;
        RECT -21.405 -83.675 -20.475 -83.345 ;
        RECT -29.625 -84.200 -29.455 -83.675 ;
        RECT -20.645 -84.200 -20.475 -83.675 ;
        RECT -20.235 -84.225 -19.945 -83.060 ;
        RECT -19.705 -83.345 -19.535 -83.060 ;
        RECT -10.725 -82.890 -10.555 -82.820 ;
        RECT -9.785 -82.890 -9.615 -82.820 ;
        RECT -10.725 -83.060 -9.615 -82.890 ;
        RECT -10.725 -83.345 -10.555 -83.060 ;
        RECT -19.705 -83.675 -18.775 -83.345 ;
        RECT -11.485 -83.675 -10.555 -83.345 ;
        RECT -19.705 -84.200 -19.535 -83.675 ;
        RECT -10.725 -84.200 -10.555 -83.675 ;
        RECT -10.315 -84.225 -10.025 -83.060 ;
        RECT -9.785 -83.345 -9.615 -83.060 ;
        RECT -0.805 -82.890 -0.635 -82.820 ;
        RECT 0.135 -82.890 0.305 -82.820 ;
        RECT -0.805 -83.060 0.305 -82.890 ;
        RECT -0.805 -83.345 -0.635 -83.060 ;
        RECT -9.785 -83.675 -8.855 -83.345 ;
        RECT -1.565 -83.675 -0.635 -83.345 ;
        RECT -9.785 -84.200 -9.615 -83.675 ;
        RECT -0.805 -84.200 -0.635 -83.675 ;
        RECT -0.395 -84.225 -0.105 -83.060 ;
        RECT 0.135 -83.345 0.305 -83.060 ;
        RECT 9.115 -82.890 9.285 -82.820 ;
        RECT 10.055 -82.890 10.225 -82.820 ;
        RECT 9.115 -83.060 10.225 -82.890 ;
        RECT 9.115 -83.345 9.285 -83.060 ;
        RECT 0.135 -83.675 1.065 -83.345 ;
        RECT 8.355 -83.675 9.285 -83.345 ;
        RECT 0.135 -84.200 0.305 -83.675 ;
        RECT 9.115 -84.200 9.285 -83.675 ;
        RECT 9.525 -84.225 9.815 -83.060 ;
        RECT 10.055 -83.345 10.225 -83.060 ;
        RECT 19.035 -82.890 19.205 -82.820 ;
        RECT 19.975 -82.890 20.145 -82.820 ;
        RECT 19.035 -83.060 20.145 -82.890 ;
        RECT 19.035 -83.345 19.205 -83.060 ;
        RECT 10.055 -83.675 10.985 -83.345 ;
        RECT 18.275 -83.675 19.205 -83.345 ;
        RECT 10.055 -84.200 10.225 -83.675 ;
        RECT 19.035 -84.200 19.205 -83.675 ;
        RECT 19.445 -84.225 19.735 -83.060 ;
        RECT 19.975 -83.345 20.145 -83.060 ;
        RECT 19.975 -83.675 20.905 -83.345 ;
        RECT 19.975 -84.200 20.145 -83.675 ;
        RECT -285.285 -172.590 -285.115 -172.440 ;
        RECT -284.345 -172.590 -284.175 -172.440 ;
        RECT -285.285 -172.760 -284.175 -172.590 ;
        RECT -285.285 -172.965 -285.115 -172.760 ;
        RECT -286.045 -173.295 -285.115 -172.965 ;
        RECT -285.285 -173.820 -285.115 -173.295 ;
        RECT -284.875 -173.925 -284.585 -172.760 ;
        RECT -284.345 -172.965 -284.175 -172.760 ;
        RECT -275.365 -172.590 -275.195 -172.440 ;
        RECT -274.425 -172.590 -274.255 -172.440 ;
        RECT -275.365 -172.760 -274.255 -172.590 ;
        RECT -275.365 -172.965 -275.195 -172.760 ;
        RECT -284.345 -173.295 -283.415 -172.965 ;
        RECT -276.125 -173.295 -275.195 -172.965 ;
        RECT -284.345 -173.820 -284.175 -173.295 ;
        RECT -275.365 -173.820 -275.195 -173.295 ;
        RECT -274.955 -173.925 -274.665 -172.760 ;
        RECT -274.425 -172.965 -274.255 -172.760 ;
        RECT -265.445 -172.590 -265.275 -172.440 ;
        RECT -264.505 -172.590 -264.335 -172.440 ;
        RECT -265.445 -172.760 -264.335 -172.590 ;
        RECT -265.445 -172.965 -265.275 -172.760 ;
        RECT -274.425 -173.295 -273.495 -172.965 ;
        RECT -266.205 -173.295 -265.275 -172.965 ;
        RECT -274.425 -173.820 -274.255 -173.295 ;
        RECT -265.445 -173.820 -265.275 -173.295 ;
        RECT -265.035 -173.925 -264.745 -172.760 ;
        RECT -264.505 -172.965 -264.335 -172.760 ;
        RECT -255.525 -172.590 -255.355 -172.440 ;
        RECT -254.585 -172.590 -254.415 -172.440 ;
        RECT -255.525 -172.760 -254.415 -172.590 ;
        RECT -255.525 -172.965 -255.355 -172.760 ;
        RECT -264.505 -173.295 -263.575 -172.965 ;
        RECT -256.285 -173.295 -255.355 -172.965 ;
        RECT -264.505 -173.820 -264.335 -173.295 ;
        RECT -255.525 -173.820 -255.355 -173.295 ;
        RECT -255.115 -173.925 -254.825 -172.760 ;
        RECT -254.585 -172.965 -254.415 -172.760 ;
        RECT -245.605 -172.590 -245.435 -172.440 ;
        RECT -244.665 -172.590 -244.495 -172.440 ;
        RECT -245.605 -172.760 -244.495 -172.590 ;
        RECT -245.605 -172.965 -245.435 -172.760 ;
        RECT -254.585 -173.295 -253.655 -172.965 ;
        RECT -246.365 -173.295 -245.435 -172.965 ;
        RECT -254.585 -173.820 -254.415 -173.295 ;
        RECT -245.605 -173.820 -245.435 -173.295 ;
        RECT -245.195 -173.925 -244.905 -172.760 ;
        RECT -244.665 -172.965 -244.495 -172.760 ;
        RECT -235.685 -172.590 -235.515 -172.440 ;
        RECT -234.745 -172.590 -234.575 -172.440 ;
        RECT -235.685 -172.760 -234.575 -172.590 ;
        RECT -235.685 -172.965 -235.515 -172.760 ;
        RECT -244.665 -173.295 -243.735 -172.965 ;
        RECT -236.445 -173.295 -235.515 -172.965 ;
        RECT -244.665 -173.820 -244.495 -173.295 ;
        RECT -235.685 -173.820 -235.515 -173.295 ;
        RECT -235.275 -173.925 -234.985 -172.760 ;
        RECT -234.745 -172.965 -234.575 -172.760 ;
        RECT -225.765 -172.590 -225.595 -172.440 ;
        RECT -224.825 -172.590 -224.655 -172.440 ;
        RECT -225.765 -172.760 -224.655 -172.590 ;
        RECT -225.765 -172.965 -225.595 -172.760 ;
        RECT -234.745 -173.295 -233.815 -172.965 ;
        RECT -226.525 -173.295 -225.595 -172.965 ;
        RECT -234.745 -173.820 -234.575 -173.295 ;
        RECT -225.765 -173.820 -225.595 -173.295 ;
        RECT -225.355 -173.925 -225.065 -172.760 ;
        RECT -224.825 -172.965 -224.655 -172.760 ;
        RECT -215.845 -172.590 -215.675 -172.440 ;
        RECT -214.905 -172.590 -214.735 -172.440 ;
        RECT -215.845 -172.760 -214.735 -172.590 ;
        RECT -215.845 -172.965 -215.675 -172.760 ;
        RECT -224.825 -173.295 -223.895 -172.965 ;
        RECT -216.605 -173.295 -215.675 -172.965 ;
        RECT -224.825 -173.820 -224.655 -173.295 ;
        RECT -215.845 -173.820 -215.675 -173.295 ;
        RECT -215.435 -173.925 -215.145 -172.760 ;
        RECT -214.905 -172.965 -214.735 -172.760 ;
        RECT -205.925 -172.590 -205.755 -172.440 ;
        RECT -204.985 -172.590 -204.815 -172.440 ;
        RECT -205.925 -172.760 -204.815 -172.590 ;
        RECT -205.925 -172.965 -205.755 -172.760 ;
        RECT -214.905 -173.295 -213.975 -172.965 ;
        RECT -206.685 -173.295 -205.755 -172.965 ;
        RECT -214.905 -173.820 -214.735 -173.295 ;
        RECT -205.925 -173.820 -205.755 -173.295 ;
        RECT -205.515 -173.925 -205.225 -172.760 ;
        RECT -204.985 -172.965 -204.815 -172.760 ;
        RECT -196.005 -172.590 -195.835 -172.440 ;
        RECT -195.065 -172.590 -194.895 -172.440 ;
        RECT -196.005 -172.760 -194.895 -172.590 ;
        RECT -196.005 -172.965 -195.835 -172.760 ;
        RECT -204.985 -173.295 -204.055 -172.965 ;
        RECT -196.765 -173.295 -195.835 -172.965 ;
        RECT -204.985 -173.820 -204.815 -173.295 ;
        RECT -196.005 -173.820 -195.835 -173.295 ;
        RECT -195.595 -173.925 -195.305 -172.760 ;
        RECT -195.065 -172.965 -194.895 -172.760 ;
        RECT -186.085 -172.590 -185.915 -172.440 ;
        RECT -185.145 -172.590 -184.975 -172.440 ;
        RECT -186.085 -172.760 -184.975 -172.590 ;
        RECT -186.085 -172.965 -185.915 -172.760 ;
        RECT -195.065 -173.295 -194.135 -172.965 ;
        RECT -186.845 -173.295 -185.915 -172.965 ;
        RECT -195.065 -173.820 -194.895 -173.295 ;
        RECT -186.085 -173.820 -185.915 -173.295 ;
        RECT -185.675 -173.925 -185.385 -172.760 ;
        RECT -185.145 -172.965 -184.975 -172.760 ;
        RECT -176.165 -172.590 -175.995 -172.440 ;
        RECT -175.225 -172.590 -175.055 -172.440 ;
        RECT -176.165 -172.760 -175.055 -172.590 ;
        RECT -176.165 -172.965 -175.995 -172.760 ;
        RECT -185.145 -173.295 -184.215 -172.965 ;
        RECT -176.925 -173.295 -175.995 -172.965 ;
        RECT -185.145 -173.820 -184.975 -173.295 ;
        RECT -176.165 -173.820 -175.995 -173.295 ;
        RECT -175.755 -173.925 -175.465 -172.760 ;
        RECT -175.225 -172.965 -175.055 -172.760 ;
        RECT -166.245 -172.590 -166.075 -172.440 ;
        RECT -165.305 -172.590 -165.135 -172.440 ;
        RECT -166.245 -172.760 -165.135 -172.590 ;
        RECT -166.245 -172.965 -166.075 -172.760 ;
        RECT -175.225 -173.295 -174.295 -172.965 ;
        RECT -167.005 -173.295 -166.075 -172.965 ;
        RECT -175.225 -173.820 -175.055 -173.295 ;
        RECT -166.245 -173.820 -166.075 -173.295 ;
        RECT -165.835 -173.925 -165.545 -172.760 ;
        RECT -165.305 -172.965 -165.135 -172.760 ;
        RECT -156.325 -172.590 -156.155 -172.440 ;
        RECT -155.385 -172.590 -155.215 -172.440 ;
        RECT -156.325 -172.760 -155.215 -172.590 ;
        RECT -156.325 -172.965 -156.155 -172.760 ;
        RECT -165.305 -173.295 -164.375 -172.965 ;
        RECT -157.085 -173.295 -156.155 -172.965 ;
        RECT -165.305 -173.820 -165.135 -173.295 ;
        RECT -156.325 -173.820 -156.155 -173.295 ;
        RECT -155.915 -173.925 -155.625 -172.760 ;
        RECT -155.385 -172.965 -155.215 -172.760 ;
        RECT -146.405 -172.590 -146.235 -172.440 ;
        RECT -145.465 -172.590 -145.295 -172.440 ;
        RECT -146.405 -172.760 -145.295 -172.590 ;
        RECT -146.405 -172.965 -146.235 -172.760 ;
        RECT -155.385 -173.295 -154.455 -172.965 ;
        RECT -147.165 -173.295 -146.235 -172.965 ;
        RECT -155.385 -173.820 -155.215 -173.295 ;
        RECT -146.405 -173.820 -146.235 -173.295 ;
        RECT -145.995 -173.925 -145.705 -172.760 ;
        RECT -145.465 -172.965 -145.295 -172.760 ;
        RECT -136.485 -172.590 -136.315 -172.440 ;
        RECT -135.545 -172.590 -135.375 -172.440 ;
        RECT -136.485 -172.760 -135.375 -172.590 ;
        RECT -136.485 -172.965 -136.315 -172.760 ;
        RECT -145.465 -173.295 -144.535 -172.965 ;
        RECT -137.245 -173.295 -136.315 -172.965 ;
        RECT -145.465 -173.820 -145.295 -173.295 ;
        RECT -136.485 -173.820 -136.315 -173.295 ;
        RECT -136.075 -173.925 -135.785 -172.760 ;
        RECT -135.545 -172.965 -135.375 -172.760 ;
        RECT -126.565 -172.590 -126.395 -172.440 ;
        RECT -125.625 -172.590 -125.455 -172.440 ;
        RECT -126.565 -172.760 -125.455 -172.590 ;
        RECT -126.565 -172.965 -126.395 -172.760 ;
        RECT -135.545 -173.295 -134.615 -172.965 ;
        RECT -127.325 -173.295 -126.395 -172.965 ;
        RECT -135.545 -173.820 -135.375 -173.295 ;
        RECT -126.565 -173.820 -126.395 -173.295 ;
        RECT -126.155 -173.925 -125.865 -172.760 ;
        RECT -125.625 -172.965 -125.455 -172.760 ;
        RECT -116.645 -172.590 -116.475 -172.440 ;
        RECT -115.705 -172.590 -115.535 -172.440 ;
        RECT -116.645 -172.760 -115.535 -172.590 ;
        RECT -116.645 -172.965 -116.475 -172.760 ;
        RECT -125.625 -173.295 -124.695 -172.965 ;
        RECT -117.405 -173.295 -116.475 -172.965 ;
        RECT -125.625 -173.820 -125.455 -173.295 ;
        RECT -116.645 -173.820 -116.475 -173.295 ;
        RECT -116.235 -173.925 -115.945 -172.760 ;
        RECT -115.705 -172.965 -115.535 -172.760 ;
        RECT -106.725 -172.590 -106.555 -172.440 ;
        RECT -105.785 -172.590 -105.615 -172.440 ;
        RECT -106.725 -172.760 -105.615 -172.590 ;
        RECT -106.725 -172.965 -106.555 -172.760 ;
        RECT -115.705 -173.295 -114.775 -172.965 ;
        RECT -107.485 -173.295 -106.555 -172.965 ;
        RECT -115.705 -173.820 -115.535 -173.295 ;
        RECT -106.725 -173.820 -106.555 -173.295 ;
        RECT -106.315 -173.925 -106.025 -172.760 ;
        RECT -105.785 -172.965 -105.615 -172.760 ;
        RECT -96.805 -172.590 -96.635 -172.440 ;
        RECT -95.865 -172.590 -95.695 -172.440 ;
        RECT -96.805 -172.760 -95.695 -172.590 ;
        RECT -96.805 -172.965 -96.635 -172.760 ;
        RECT -105.785 -173.295 -104.855 -172.965 ;
        RECT -97.565 -173.295 -96.635 -172.965 ;
        RECT -105.785 -173.820 -105.615 -173.295 ;
        RECT -96.805 -173.820 -96.635 -173.295 ;
        RECT -96.395 -173.925 -96.105 -172.760 ;
        RECT -95.865 -172.965 -95.695 -172.760 ;
        RECT -86.885 -172.590 -86.715 -172.440 ;
        RECT -85.945 -172.590 -85.775 -172.440 ;
        RECT -86.885 -172.760 -85.775 -172.590 ;
        RECT -86.885 -172.965 -86.715 -172.760 ;
        RECT -95.865 -173.295 -94.935 -172.965 ;
        RECT -87.645 -173.295 -86.715 -172.965 ;
        RECT -95.865 -173.820 -95.695 -173.295 ;
        RECT -86.885 -173.820 -86.715 -173.295 ;
        RECT -86.475 -173.925 -86.185 -172.760 ;
        RECT -85.945 -172.965 -85.775 -172.760 ;
        RECT -76.965 -172.590 -76.795 -172.440 ;
        RECT -76.025 -172.590 -75.855 -172.440 ;
        RECT -76.965 -172.760 -75.855 -172.590 ;
        RECT -76.965 -172.965 -76.795 -172.760 ;
        RECT -85.945 -173.295 -85.015 -172.965 ;
        RECT -77.725 -173.295 -76.795 -172.965 ;
        RECT -85.945 -173.820 -85.775 -173.295 ;
        RECT -76.965 -173.820 -76.795 -173.295 ;
        RECT -76.555 -173.925 -76.265 -172.760 ;
        RECT -76.025 -172.965 -75.855 -172.760 ;
        RECT -67.045 -172.590 -66.875 -172.440 ;
        RECT -66.105 -172.590 -65.935 -172.440 ;
        RECT -67.045 -172.760 -65.935 -172.590 ;
        RECT -67.045 -172.965 -66.875 -172.760 ;
        RECT -76.025 -173.295 -75.095 -172.965 ;
        RECT -67.805 -173.295 -66.875 -172.965 ;
        RECT -76.025 -173.820 -75.855 -173.295 ;
        RECT -67.045 -173.820 -66.875 -173.295 ;
        RECT -66.635 -173.925 -66.345 -172.760 ;
        RECT -66.105 -172.965 -65.935 -172.760 ;
        RECT -57.125 -172.590 -56.955 -172.440 ;
        RECT -56.185 -172.590 -56.015 -172.440 ;
        RECT -57.125 -172.760 -56.015 -172.590 ;
        RECT -57.125 -172.965 -56.955 -172.760 ;
        RECT -66.105 -173.295 -65.175 -172.965 ;
        RECT -57.885 -173.295 -56.955 -172.965 ;
        RECT -66.105 -173.820 -65.935 -173.295 ;
        RECT -57.125 -173.820 -56.955 -173.295 ;
        RECT -56.715 -173.925 -56.425 -172.760 ;
        RECT -56.185 -172.965 -56.015 -172.760 ;
        RECT -47.205 -172.590 -47.035 -172.440 ;
        RECT -46.265 -172.590 -46.095 -172.440 ;
        RECT -47.205 -172.760 -46.095 -172.590 ;
        RECT -47.205 -172.965 -47.035 -172.760 ;
        RECT -56.185 -173.295 -55.255 -172.965 ;
        RECT -47.965 -173.295 -47.035 -172.965 ;
        RECT -56.185 -173.820 -56.015 -173.295 ;
        RECT -47.205 -173.820 -47.035 -173.295 ;
        RECT -46.795 -173.925 -46.505 -172.760 ;
        RECT -46.265 -172.965 -46.095 -172.760 ;
        RECT -37.285 -172.590 -37.115 -172.440 ;
        RECT -36.345 -172.590 -36.175 -172.440 ;
        RECT -37.285 -172.760 -36.175 -172.590 ;
        RECT -37.285 -172.965 -37.115 -172.760 ;
        RECT -46.265 -173.295 -45.335 -172.965 ;
        RECT -38.045 -173.295 -37.115 -172.965 ;
        RECT -46.265 -173.820 -46.095 -173.295 ;
        RECT -37.285 -173.820 -37.115 -173.295 ;
        RECT -36.875 -173.925 -36.585 -172.760 ;
        RECT -36.345 -172.965 -36.175 -172.760 ;
        RECT -27.365 -172.590 -27.195 -172.440 ;
        RECT -26.425 -172.590 -26.255 -172.440 ;
        RECT -27.365 -172.760 -26.255 -172.590 ;
        RECT -27.365 -172.965 -27.195 -172.760 ;
        RECT -36.345 -173.295 -35.415 -172.965 ;
        RECT -28.125 -173.295 -27.195 -172.965 ;
        RECT -36.345 -173.820 -36.175 -173.295 ;
        RECT -27.365 -173.820 -27.195 -173.295 ;
        RECT -26.955 -173.925 -26.665 -172.760 ;
        RECT -26.425 -172.965 -26.255 -172.760 ;
        RECT -17.445 -172.590 -17.275 -172.440 ;
        RECT -16.505 -172.590 -16.335 -172.440 ;
        RECT -17.445 -172.760 -16.335 -172.590 ;
        RECT -17.445 -172.965 -17.275 -172.760 ;
        RECT -26.425 -173.295 -25.495 -172.965 ;
        RECT -18.205 -173.295 -17.275 -172.965 ;
        RECT -26.425 -173.820 -26.255 -173.295 ;
        RECT -17.445 -173.820 -17.275 -173.295 ;
        RECT -17.035 -173.925 -16.745 -172.760 ;
        RECT -16.505 -172.965 -16.335 -172.760 ;
        RECT -7.525 -172.590 -7.355 -172.440 ;
        RECT -6.585 -172.590 -6.415 -172.440 ;
        RECT -7.525 -172.760 -6.415 -172.590 ;
        RECT -7.525 -172.965 -7.355 -172.760 ;
        RECT -16.505 -173.295 -15.575 -172.965 ;
        RECT -8.285 -173.295 -7.355 -172.965 ;
        RECT -16.505 -173.820 -16.335 -173.295 ;
        RECT -7.525 -173.820 -7.355 -173.295 ;
        RECT -7.115 -173.925 -6.825 -172.760 ;
        RECT -6.585 -172.965 -6.415 -172.760 ;
        RECT 2.395 -172.590 2.565 -172.440 ;
        RECT 3.335 -172.590 3.505 -172.440 ;
        RECT 2.395 -172.760 3.505 -172.590 ;
        RECT 2.395 -172.965 2.565 -172.760 ;
        RECT -6.585 -173.295 -5.655 -172.965 ;
        RECT 1.635 -173.295 2.565 -172.965 ;
        RECT -6.585 -173.820 -6.415 -173.295 ;
        RECT 2.395 -173.820 2.565 -173.295 ;
        RECT 2.805 -173.925 3.095 -172.760 ;
        RECT 3.335 -172.965 3.505 -172.760 ;
        RECT 12.315 -172.590 12.485 -172.440 ;
        RECT 13.255 -172.590 13.425 -172.440 ;
        RECT 12.315 -172.760 13.425 -172.590 ;
        RECT 12.315 -172.965 12.485 -172.760 ;
        RECT 3.335 -173.295 4.265 -172.965 ;
        RECT 11.555 -173.295 12.485 -172.965 ;
        RECT 3.335 -173.820 3.505 -173.295 ;
        RECT 12.315 -173.820 12.485 -173.295 ;
        RECT 12.725 -173.925 13.015 -172.760 ;
        RECT 13.255 -172.965 13.425 -172.760 ;
        RECT 22.235 -172.590 22.405 -172.440 ;
        RECT 22.235 -172.760 23.020 -172.590 ;
        RECT 22.235 -172.965 22.405 -172.760 ;
        RECT 13.255 -173.295 14.185 -172.965 ;
        RECT 21.475 -173.295 22.405 -172.965 ;
        RECT 13.255 -173.820 13.425 -173.295 ;
        RECT 22.235 -173.820 22.405 -173.295 ;
        RECT 22.645 -173.925 22.935 -172.760 ;
        RECT -291.300 -174.335 -288.080 -174.165 ;
        RECT -281.380 -174.335 -278.160 -174.165 ;
        RECT -271.460 -174.335 -268.240 -174.165 ;
        RECT -261.540 -174.335 -258.320 -174.165 ;
        RECT -251.620 -174.335 -248.400 -174.165 ;
        RECT -241.700 -174.335 -238.480 -174.165 ;
        RECT -231.780 -174.335 -228.560 -174.165 ;
        RECT -221.860 -174.335 -218.640 -174.165 ;
        RECT -211.940 -174.335 -208.720 -174.165 ;
        RECT -202.020 -174.335 -198.800 -174.165 ;
        RECT -192.100 -174.335 -188.880 -174.165 ;
        RECT -182.180 -174.335 -178.960 -174.165 ;
        RECT -172.260 -174.335 -169.040 -174.165 ;
        RECT -162.340 -174.335 -159.120 -174.165 ;
        RECT -152.420 -174.335 -149.200 -174.165 ;
        RECT -142.500 -174.335 -139.280 -174.165 ;
        RECT -132.580 -174.335 -129.360 -174.165 ;
        RECT -122.660 -174.335 -119.440 -174.165 ;
        RECT -112.740 -174.335 -109.520 -174.165 ;
        RECT -102.820 -174.335 -99.600 -174.165 ;
        RECT -92.900 -174.335 -89.680 -174.165 ;
        RECT -82.980 -174.335 -79.760 -174.165 ;
        RECT -73.060 -174.335 -69.840 -174.165 ;
        RECT -63.140 -174.335 -59.920 -174.165 ;
        RECT -53.220 -174.335 -50.000 -174.165 ;
        RECT -43.300 -174.335 -40.080 -174.165 ;
        RECT -33.380 -174.335 -30.160 -174.165 ;
        RECT -23.460 -174.335 -20.240 -174.165 ;
        RECT -13.540 -174.335 -10.320 -174.165 ;
        RECT -3.620 -174.335 -0.400 -174.165 ;
        RECT 6.300 -174.335 9.520 -174.165 ;
        RECT 16.220 -174.335 19.440 -174.165 ;
        RECT -291.215 -175.475 -290.955 -174.335 ;
        RECT -290.285 -175.475 -290.005 -174.335 ;
        RECT -289.835 -175.500 -289.545 -174.335 ;
        RECT -289.375 -175.475 -289.095 -174.335 ;
        RECT -288.425 -175.475 -288.165 -174.335 ;
        RECT -281.295 -175.475 -281.035 -174.335 ;
        RECT -280.365 -175.475 -280.085 -174.335 ;
        RECT -279.915 -175.500 -279.625 -174.335 ;
        RECT -279.455 -175.475 -279.175 -174.335 ;
        RECT -278.505 -175.475 -278.245 -174.335 ;
        RECT -271.375 -175.475 -271.115 -174.335 ;
        RECT -270.445 -175.475 -270.165 -174.335 ;
        RECT -269.995 -175.500 -269.705 -174.335 ;
        RECT -269.535 -175.475 -269.255 -174.335 ;
        RECT -268.585 -175.475 -268.325 -174.335 ;
        RECT -261.455 -175.475 -261.195 -174.335 ;
        RECT -260.525 -175.475 -260.245 -174.335 ;
        RECT -260.075 -175.500 -259.785 -174.335 ;
        RECT -259.615 -175.475 -259.335 -174.335 ;
        RECT -258.665 -175.475 -258.405 -174.335 ;
        RECT -251.535 -175.475 -251.275 -174.335 ;
        RECT -250.605 -175.475 -250.325 -174.335 ;
        RECT -250.155 -175.500 -249.865 -174.335 ;
        RECT -249.695 -175.475 -249.415 -174.335 ;
        RECT -248.745 -175.475 -248.485 -174.335 ;
        RECT -241.615 -175.475 -241.355 -174.335 ;
        RECT -240.685 -175.475 -240.405 -174.335 ;
        RECT -240.235 -175.500 -239.945 -174.335 ;
        RECT -239.775 -175.475 -239.495 -174.335 ;
        RECT -238.825 -175.475 -238.565 -174.335 ;
        RECT -231.695 -175.475 -231.435 -174.335 ;
        RECT -230.765 -175.475 -230.485 -174.335 ;
        RECT -230.315 -175.500 -230.025 -174.335 ;
        RECT -229.855 -175.475 -229.575 -174.335 ;
        RECT -228.905 -175.475 -228.645 -174.335 ;
        RECT -221.775 -175.475 -221.515 -174.335 ;
        RECT -220.845 -175.475 -220.565 -174.335 ;
        RECT -220.395 -175.500 -220.105 -174.335 ;
        RECT -219.935 -175.475 -219.655 -174.335 ;
        RECT -218.985 -175.475 -218.725 -174.335 ;
        RECT -211.855 -175.475 -211.595 -174.335 ;
        RECT -210.925 -175.475 -210.645 -174.335 ;
        RECT -210.475 -175.500 -210.185 -174.335 ;
        RECT -210.015 -175.475 -209.735 -174.335 ;
        RECT -209.065 -175.475 -208.805 -174.335 ;
        RECT -201.935 -175.475 -201.675 -174.335 ;
        RECT -201.005 -175.475 -200.725 -174.335 ;
        RECT -200.555 -175.500 -200.265 -174.335 ;
        RECT -200.095 -175.475 -199.815 -174.335 ;
        RECT -199.145 -175.475 -198.885 -174.335 ;
        RECT -192.015 -175.475 -191.755 -174.335 ;
        RECT -191.085 -175.475 -190.805 -174.335 ;
        RECT -190.635 -175.500 -190.345 -174.335 ;
        RECT -190.175 -175.475 -189.895 -174.335 ;
        RECT -189.225 -175.475 -188.965 -174.335 ;
        RECT -182.095 -175.475 -181.835 -174.335 ;
        RECT -181.165 -175.475 -180.885 -174.335 ;
        RECT -180.715 -175.500 -180.425 -174.335 ;
        RECT -180.255 -175.475 -179.975 -174.335 ;
        RECT -179.305 -175.475 -179.045 -174.335 ;
        RECT -172.175 -175.475 -171.915 -174.335 ;
        RECT -171.245 -175.475 -170.965 -174.335 ;
        RECT -170.795 -175.500 -170.505 -174.335 ;
        RECT -170.335 -175.475 -170.055 -174.335 ;
        RECT -169.385 -175.475 -169.125 -174.335 ;
        RECT -162.255 -175.475 -161.995 -174.335 ;
        RECT -161.325 -175.475 -161.045 -174.335 ;
        RECT -160.875 -175.500 -160.585 -174.335 ;
        RECT -160.415 -175.475 -160.135 -174.335 ;
        RECT -159.465 -175.475 -159.205 -174.335 ;
        RECT -152.335 -175.475 -152.075 -174.335 ;
        RECT -151.405 -175.475 -151.125 -174.335 ;
        RECT -150.955 -175.500 -150.665 -174.335 ;
        RECT -150.495 -175.475 -150.215 -174.335 ;
        RECT -149.545 -175.475 -149.285 -174.335 ;
        RECT -142.415 -175.475 -142.155 -174.335 ;
        RECT -141.485 -175.475 -141.205 -174.335 ;
        RECT -141.035 -175.500 -140.745 -174.335 ;
        RECT -140.575 -175.475 -140.295 -174.335 ;
        RECT -139.625 -175.475 -139.365 -174.335 ;
        RECT -132.495 -175.475 -132.235 -174.335 ;
        RECT -131.565 -175.475 -131.285 -174.335 ;
        RECT -131.115 -175.500 -130.825 -174.335 ;
        RECT -130.655 -175.475 -130.375 -174.335 ;
        RECT -129.705 -175.475 -129.445 -174.335 ;
        RECT -122.575 -175.475 -122.315 -174.335 ;
        RECT -121.645 -175.475 -121.365 -174.335 ;
        RECT -121.195 -175.500 -120.905 -174.335 ;
        RECT -120.735 -175.475 -120.455 -174.335 ;
        RECT -119.785 -175.475 -119.525 -174.335 ;
        RECT -112.655 -175.475 -112.395 -174.335 ;
        RECT -111.725 -175.475 -111.445 -174.335 ;
        RECT -111.275 -175.500 -110.985 -174.335 ;
        RECT -110.815 -175.475 -110.535 -174.335 ;
        RECT -109.865 -175.475 -109.605 -174.335 ;
        RECT -102.735 -175.475 -102.475 -174.335 ;
        RECT -101.805 -175.475 -101.525 -174.335 ;
        RECT -101.355 -175.500 -101.065 -174.335 ;
        RECT -100.895 -175.475 -100.615 -174.335 ;
        RECT -99.945 -175.475 -99.685 -174.335 ;
        RECT -92.815 -175.475 -92.555 -174.335 ;
        RECT -91.885 -175.475 -91.605 -174.335 ;
        RECT -91.435 -175.500 -91.145 -174.335 ;
        RECT -90.975 -175.475 -90.695 -174.335 ;
        RECT -90.025 -175.475 -89.765 -174.335 ;
        RECT -82.895 -175.475 -82.635 -174.335 ;
        RECT -81.965 -175.475 -81.685 -174.335 ;
        RECT -81.515 -175.500 -81.225 -174.335 ;
        RECT -81.055 -175.475 -80.775 -174.335 ;
        RECT -80.105 -175.475 -79.845 -174.335 ;
        RECT -72.975 -175.475 -72.715 -174.335 ;
        RECT -72.045 -175.475 -71.765 -174.335 ;
        RECT -71.595 -175.500 -71.305 -174.335 ;
        RECT -71.135 -175.475 -70.855 -174.335 ;
        RECT -70.185 -175.475 -69.925 -174.335 ;
        RECT -63.055 -175.475 -62.795 -174.335 ;
        RECT -62.125 -175.475 -61.845 -174.335 ;
        RECT -61.675 -175.500 -61.385 -174.335 ;
        RECT -61.215 -175.475 -60.935 -174.335 ;
        RECT -60.265 -175.475 -60.005 -174.335 ;
        RECT -53.135 -175.475 -52.875 -174.335 ;
        RECT -52.205 -175.475 -51.925 -174.335 ;
        RECT -51.755 -175.500 -51.465 -174.335 ;
        RECT -51.295 -175.475 -51.015 -174.335 ;
        RECT -50.345 -175.475 -50.085 -174.335 ;
        RECT -43.215 -175.475 -42.955 -174.335 ;
        RECT -42.285 -175.475 -42.005 -174.335 ;
        RECT -41.835 -175.500 -41.545 -174.335 ;
        RECT -41.375 -175.475 -41.095 -174.335 ;
        RECT -40.425 -175.475 -40.165 -174.335 ;
        RECT -33.295 -175.475 -33.035 -174.335 ;
        RECT -32.365 -175.475 -32.085 -174.335 ;
        RECT -31.915 -175.500 -31.625 -174.335 ;
        RECT -31.455 -175.475 -31.175 -174.335 ;
        RECT -30.505 -175.475 -30.245 -174.335 ;
        RECT -23.375 -175.475 -23.115 -174.335 ;
        RECT -22.445 -175.475 -22.165 -174.335 ;
        RECT -21.995 -175.500 -21.705 -174.335 ;
        RECT -21.535 -175.475 -21.255 -174.335 ;
        RECT -20.585 -175.475 -20.325 -174.335 ;
        RECT -13.455 -175.475 -13.195 -174.335 ;
        RECT -12.525 -175.475 -12.245 -174.335 ;
        RECT -12.075 -175.500 -11.785 -174.335 ;
        RECT -11.615 -175.475 -11.335 -174.335 ;
        RECT -10.665 -175.475 -10.405 -174.335 ;
        RECT -3.535 -175.475 -3.275 -174.335 ;
        RECT -2.605 -175.475 -2.325 -174.335 ;
        RECT -2.155 -175.500 -1.865 -174.335 ;
        RECT -1.695 -175.475 -1.415 -174.335 ;
        RECT -0.745 -175.475 -0.485 -174.335 ;
        RECT 6.385 -175.475 6.645 -174.335 ;
        RECT 7.315 -175.475 7.595 -174.335 ;
        RECT 7.765 -175.500 8.055 -174.335 ;
        RECT 8.225 -175.475 8.505 -174.335 ;
        RECT 9.175 -175.475 9.435 -174.335 ;
        RECT 16.305 -175.475 16.565 -174.335 ;
        RECT 17.235 -175.475 17.515 -174.335 ;
        RECT 17.685 -175.500 17.975 -174.335 ;
        RECT 18.145 -175.475 18.425 -174.335 ;
        RECT 19.095 -175.475 19.355 -174.335 ;
        RECT -286.255 -176.885 -285.995 -175.745 ;
        RECT -285.325 -176.885 -285.045 -175.745 ;
        RECT -284.875 -176.885 -284.585 -175.720 ;
        RECT -284.415 -176.885 -284.135 -175.745 ;
        RECT -283.465 -176.885 -283.205 -175.745 ;
        RECT -276.335 -176.885 -276.075 -175.745 ;
        RECT -275.405 -176.885 -275.125 -175.745 ;
        RECT -274.955 -176.885 -274.665 -175.720 ;
        RECT -274.495 -176.885 -274.215 -175.745 ;
        RECT -273.545 -176.885 -273.285 -175.745 ;
        RECT -266.415 -176.885 -266.155 -175.745 ;
        RECT -265.485 -176.885 -265.205 -175.745 ;
        RECT -265.035 -176.885 -264.745 -175.720 ;
        RECT -264.575 -176.885 -264.295 -175.745 ;
        RECT -263.625 -176.885 -263.365 -175.745 ;
        RECT -256.495 -176.885 -256.235 -175.745 ;
        RECT -255.565 -176.885 -255.285 -175.745 ;
        RECT -255.115 -176.885 -254.825 -175.720 ;
        RECT -254.655 -176.885 -254.375 -175.745 ;
        RECT -253.705 -176.885 -253.445 -175.745 ;
        RECT -246.575 -176.885 -246.315 -175.745 ;
        RECT -245.645 -176.885 -245.365 -175.745 ;
        RECT -245.195 -176.885 -244.905 -175.720 ;
        RECT -244.735 -176.885 -244.455 -175.745 ;
        RECT -243.785 -176.885 -243.525 -175.745 ;
        RECT -236.655 -176.885 -236.395 -175.745 ;
        RECT -235.725 -176.885 -235.445 -175.745 ;
        RECT -235.275 -176.885 -234.985 -175.720 ;
        RECT -234.815 -176.885 -234.535 -175.745 ;
        RECT -233.865 -176.885 -233.605 -175.745 ;
        RECT -226.735 -176.885 -226.475 -175.745 ;
        RECT -225.805 -176.885 -225.525 -175.745 ;
        RECT -225.355 -176.885 -225.065 -175.720 ;
        RECT -224.895 -176.885 -224.615 -175.745 ;
        RECT -223.945 -176.885 -223.685 -175.745 ;
        RECT -216.815 -176.885 -216.555 -175.745 ;
        RECT -215.885 -176.885 -215.605 -175.745 ;
        RECT -215.435 -176.885 -215.145 -175.720 ;
        RECT -214.975 -176.885 -214.695 -175.745 ;
        RECT -214.025 -176.885 -213.765 -175.745 ;
        RECT -206.895 -176.885 -206.635 -175.745 ;
        RECT -205.965 -176.885 -205.685 -175.745 ;
        RECT -205.515 -176.885 -205.225 -175.720 ;
        RECT -205.055 -176.885 -204.775 -175.745 ;
        RECT -204.105 -176.885 -203.845 -175.745 ;
        RECT -196.975 -176.885 -196.715 -175.745 ;
        RECT -196.045 -176.885 -195.765 -175.745 ;
        RECT -195.595 -176.885 -195.305 -175.720 ;
        RECT -195.135 -176.885 -194.855 -175.745 ;
        RECT -194.185 -176.885 -193.925 -175.745 ;
        RECT -187.055 -176.885 -186.795 -175.745 ;
        RECT -186.125 -176.885 -185.845 -175.745 ;
        RECT -185.675 -176.885 -185.385 -175.720 ;
        RECT -185.215 -176.885 -184.935 -175.745 ;
        RECT -184.265 -176.885 -184.005 -175.745 ;
        RECT -177.135 -176.885 -176.875 -175.745 ;
        RECT -176.205 -176.885 -175.925 -175.745 ;
        RECT -175.755 -176.885 -175.465 -175.720 ;
        RECT -175.295 -176.885 -175.015 -175.745 ;
        RECT -174.345 -176.885 -174.085 -175.745 ;
        RECT -167.215 -176.885 -166.955 -175.745 ;
        RECT -166.285 -176.885 -166.005 -175.745 ;
        RECT -165.835 -176.885 -165.545 -175.720 ;
        RECT -165.375 -176.885 -165.095 -175.745 ;
        RECT -164.425 -176.885 -164.165 -175.745 ;
        RECT -157.295 -176.885 -157.035 -175.745 ;
        RECT -156.365 -176.885 -156.085 -175.745 ;
        RECT -155.915 -176.885 -155.625 -175.720 ;
        RECT -155.455 -176.885 -155.175 -175.745 ;
        RECT -154.505 -176.885 -154.245 -175.745 ;
        RECT -147.375 -176.885 -147.115 -175.745 ;
        RECT -146.445 -176.885 -146.165 -175.745 ;
        RECT -145.995 -176.885 -145.705 -175.720 ;
        RECT -145.535 -176.885 -145.255 -175.745 ;
        RECT -144.585 -176.885 -144.325 -175.745 ;
        RECT -137.455 -176.885 -137.195 -175.745 ;
        RECT -136.525 -176.885 -136.245 -175.745 ;
        RECT -136.075 -176.885 -135.785 -175.720 ;
        RECT -135.615 -176.885 -135.335 -175.745 ;
        RECT -134.665 -176.885 -134.405 -175.745 ;
        RECT -127.535 -176.885 -127.275 -175.745 ;
        RECT -126.605 -176.885 -126.325 -175.745 ;
        RECT -126.155 -176.885 -125.865 -175.720 ;
        RECT -125.695 -176.885 -125.415 -175.745 ;
        RECT -124.745 -176.885 -124.485 -175.745 ;
        RECT -117.615 -176.885 -117.355 -175.745 ;
        RECT -116.685 -176.885 -116.405 -175.745 ;
        RECT -116.235 -176.885 -115.945 -175.720 ;
        RECT -115.775 -176.885 -115.495 -175.745 ;
        RECT -114.825 -176.885 -114.565 -175.745 ;
        RECT -107.695 -176.885 -107.435 -175.745 ;
        RECT -106.765 -176.885 -106.485 -175.745 ;
        RECT -106.315 -176.885 -106.025 -175.720 ;
        RECT -105.855 -176.885 -105.575 -175.745 ;
        RECT -104.905 -176.885 -104.645 -175.745 ;
        RECT -97.775 -176.885 -97.515 -175.745 ;
        RECT -96.845 -176.885 -96.565 -175.745 ;
        RECT -96.395 -176.885 -96.105 -175.720 ;
        RECT -95.935 -176.885 -95.655 -175.745 ;
        RECT -94.985 -176.885 -94.725 -175.745 ;
        RECT -87.855 -176.885 -87.595 -175.745 ;
        RECT -86.925 -176.885 -86.645 -175.745 ;
        RECT -86.475 -176.885 -86.185 -175.720 ;
        RECT -86.015 -176.885 -85.735 -175.745 ;
        RECT -85.065 -176.885 -84.805 -175.745 ;
        RECT -77.935 -176.885 -77.675 -175.745 ;
        RECT -77.005 -176.885 -76.725 -175.745 ;
        RECT -76.555 -176.885 -76.265 -175.720 ;
        RECT -76.095 -176.885 -75.815 -175.745 ;
        RECT -75.145 -176.885 -74.885 -175.745 ;
        RECT -68.015 -176.885 -67.755 -175.745 ;
        RECT -67.085 -176.885 -66.805 -175.745 ;
        RECT -66.635 -176.885 -66.345 -175.720 ;
        RECT -66.175 -176.885 -65.895 -175.745 ;
        RECT -65.225 -176.885 -64.965 -175.745 ;
        RECT -58.095 -176.885 -57.835 -175.745 ;
        RECT -57.165 -176.885 -56.885 -175.745 ;
        RECT -56.715 -176.885 -56.425 -175.720 ;
        RECT -56.255 -176.885 -55.975 -175.745 ;
        RECT -55.305 -176.885 -55.045 -175.745 ;
        RECT -48.175 -176.885 -47.915 -175.745 ;
        RECT -47.245 -176.885 -46.965 -175.745 ;
        RECT -46.795 -176.885 -46.505 -175.720 ;
        RECT -46.335 -176.885 -46.055 -175.745 ;
        RECT -45.385 -176.885 -45.125 -175.745 ;
        RECT -38.255 -176.885 -37.995 -175.745 ;
        RECT -37.325 -176.885 -37.045 -175.745 ;
        RECT -36.875 -176.885 -36.585 -175.720 ;
        RECT -36.415 -176.885 -36.135 -175.745 ;
        RECT -35.465 -176.885 -35.205 -175.745 ;
        RECT -28.335 -176.885 -28.075 -175.745 ;
        RECT -27.405 -176.885 -27.125 -175.745 ;
        RECT -26.955 -176.885 -26.665 -175.720 ;
        RECT -26.495 -176.885 -26.215 -175.745 ;
        RECT -25.545 -176.885 -25.285 -175.745 ;
        RECT -18.415 -176.885 -18.155 -175.745 ;
        RECT -17.485 -176.885 -17.205 -175.745 ;
        RECT -17.035 -176.885 -16.745 -175.720 ;
        RECT -16.575 -176.885 -16.295 -175.745 ;
        RECT -15.625 -176.885 -15.365 -175.745 ;
        RECT -8.495 -176.885 -8.235 -175.745 ;
        RECT -7.565 -176.885 -7.285 -175.745 ;
        RECT -7.115 -176.885 -6.825 -175.720 ;
        RECT -6.655 -176.885 -6.375 -175.745 ;
        RECT -5.705 -176.885 -5.445 -175.745 ;
        RECT 1.425 -176.885 1.685 -175.745 ;
        RECT 2.355 -176.885 2.635 -175.745 ;
        RECT 2.805 -176.885 3.095 -175.720 ;
        RECT 3.265 -176.885 3.545 -175.745 ;
        RECT 4.215 -176.885 4.475 -175.745 ;
        RECT 11.345 -176.885 11.605 -175.745 ;
        RECT 12.275 -176.885 12.555 -175.745 ;
        RECT 12.725 -176.885 13.015 -175.720 ;
        RECT 13.185 -176.885 13.465 -175.745 ;
        RECT 14.135 -176.885 14.395 -175.745 ;
        RECT 21.265 -176.885 21.525 -175.745 ;
        RECT 22.195 -176.885 22.475 -175.745 ;
        RECT 22.645 -176.885 22.935 -175.720 ;
        RECT -286.340 -177.055 -283.120 -176.885 ;
        RECT -276.420 -177.055 -273.200 -176.885 ;
        RECT -266.500 -177.055 -263.280 -176.885 ;
        RECT -256.580 -177.055 -253.360 -176.885 ;
        RECT -246.660 -177.055 -243.440 -176.885 ;
        RECT -236.740 -177.055 -233.520 -176.885 ;
        RECT -226.820 -177.055 -223.600 -176.885 ;
        RECT -216.900 -177.055 -213.680 -176.885 ;
        RECT -206.980 -177.055 -203.760 -176.885 ;
        RECT -197.060 -177.055 -193.840 -176.885 ;
        RECT -187.140 -177.055 -183.920 -176.885 ;
        RECT -177.220 -177.055 -174.000 -176.885 ;
        RECT -167.300 -177.055 -164.080 -176.885 ;
        RECT -157.380 -177.055 -154.160 -176.885 ;
        RECT -147.460 -177.055 -144.240 -176.885 ;
        RECT -137.540 -177.055 -134.320 -176.885 ;
        RECT -127.620 -177.055 -124.400 -176.885 ;
        RECT -117.700 -177.055 -114.480 -176.885 ;
        RECT -107.780 -177.055 -104.560 -176.885 ;
        RECT -97.860 -177.055 -94.640 -176.885 ;
        RECT -87.940 -177.055 -84.720 -176.885 ;
        RECT -78.020 -177.055 -74.800 -176.885 ;
        RECT -68.100 -177.055 -64.880 -176.885 ;
        RECT -58.180 -177.055 -54.960 -176.885 ;
        RECT -48.260 -177.055 -45.040 -176.885 ;
        RECT -38.340 -177.055 -35.120 -176.885 ;
        RECT -28.420 -177.055 -25.200 -176.885 ;
        RECT -18.500 -177.055 -15.280 -176.885 ;
        RECT -8.580 -177.055 -5.360 -176.885 ;
        RECT 1.340 -177.055 4.560 -176.885 ;
        RECT 11.260 -177.055 14.480 -176.885 ;
        RECT 21.180 -177.055 23.020 -176.885 ;
        RECT -290.245 -177.470 -290.075 -177.400 ;
        RECT -289.305 -177.470 -289.135 -177.400 ;
        RECT -290.245 -177.640 -289.135 -177.470 ;
        RECT -290.245 -177.925 -290.075 -177.640 ;
        RECT -291.005 -178.255 -290.075 -177.925 ;
        RECT -290.245 -178.780 -290.075 -178.255 ;
        RECT -289.835 -178.805 -289.545 -177.640 ;
        RECT -289.305 -177.925 -289.135 -177.640 ;
        RECT -280.325 -177.470 -280.155 -177.400 ;
        RECT -279.385 -177.470 -279.215 -177.400 ;
        RECT -280.325 -177.640 -279.215 -177.470 ;
        RECT -280.325 -177.925 -280.155 -177.640 ;
        RECT -289.305 -178.255 -288.375 -177.925 ;
        RECT -281.085 -178.255 -280.155 -177.925 ;
        RECT -289.305 -178.780 -289.135 -178.255 ;
        RECT -280.325 -178.780 -280.155 -178.255 ;
        RECT -279.915 -178.805 -279.625 -177.640 ;
        RECT -279.385 -177.925 -279.215 -177.640 ;
        RECT -270.405 -177.470 -270.235 -177.400 ;
        RECT -269.465 -177.470 -269.295 -177.400 ;
        RECT -270.405 -177.640 -269.295 -177.470 ;
        RECT -270.405 -177.925 -270.235 -177.640 ;
        RECT -279.385 -178.255 -278.455 -177.925 ;
        RECT -271.165 -178.255 -270.235 -177.925 ;
        RECT -279.385 -178.780 -279.215 -178.255 ;
        RECT -270.405 -178.780 -270.235 -178.255 ;
        RECT -269.995 -178.805 -269.705 -177.640 ;
        RECT -269.465 -177.925 -269.295 -177.640 ;
        RECT -260.485 -177.470 -260.315 -177.400 ;
        RECT -259.545 -177.470 -259.375 -177.400 ;
        RECT -260.485 -177.640 -259.375 -177.470 ;
        RECT -260.485 -177.925 -260.315 -177.640 ;
        RECT -269.465 -178.255 -268.535 -177.925 ;
        RECT -261.245 -178.255 -260.315 -177.925 ;
        RECT -269.465 -178.780 -269.295 -178.255 ;
        RECT -260.485 -178.780 -260.315 -178.255 ;
        RECT -260.075 -178.805 -259.785 -177.640 ;
        RECT -259.545 -177.925 -259.375 -177.640 ;
        RECT -250.565 -177.470 -250.395 -177.400 ;
        RECT -249.625 -177.470 -249.455 -177.400 ;
        RECT -250.565 -177.640 -249.455 -177.470 ;
        RECT -250.565 -177.925 -250.395 -177.640 ;
        RECT -259.545 -178.255 -258.615 -177.925 ;
        RECT -251.325 -178.255 -250.395 -177.925 ;
        RECT -259.545 -178.780 -259.375 -178.255 ;
        RECT -250.565 -178.780 -250.395 -178.255 ;
        RECT -250.155 -178.805 -249.865 -177.640 ;
        RECT -249.625 -177.925 -249.455 -177.640 ;
        RECT -240.645 -177.470 -240.475 -177.400 ;
        RECT -239.705 -177.470 -239.535 -177.400 ;
        RECT -240.645 -177.640 -239.535 -177.470 ;
        RECT -240.645 -177.925 -240.475 -177.640 ;
        RECT -249.625 -178.255 -248.695 -177.925 ;
        RECT -241.405 -178.255 -240.475 -177.925 ;
        RECT -249.625 -178.780 -249.455 -178.255 ;
        RECT -240.645 -178.780 -240.475 -178.255 ;
        RECT -240.235 -178.805 -239.945 -177.640 ;
        RECT -239.705 -177.925 -239.535 -177.640 ;
        RECT -230.725 -177.470 -230.555 -177.400 ;
        RECT -229.785 -177.470 -229.615 -177.400 ;
        RECT -230.725 -177.640 -229.615 -177.470 ;
        RECT -230.725 -177.925 -230.555 -177.640 ;
        RECT -239.705 -178.255 -238.775 -177.925 ;
        RECT -231.485 -178.255 -230.555 -177.925 ;
        RECT -239.705 -178.780 -239.535 -178.255 ;
        RECT -230.725 -178.780 -230.555 -178.255 ;
        RECT -230.315 -178.805 -230.025 -177.640 ;
        RECT -229.785 -177.925 -229.615 -177.640 ;
        RECT -220.805 -177.470 -220.635 -177.400 ;
        RECT -219.865 -177.470 -219.695 -177.400 ;
        RECT -220.805 -177.640 -219.695 -177.470 ;
        RECT -220.805 -177.925 -220.635 -177.640 ;
        RECT -229.785 -178.255 -228.855 -177.925 ;
        RECT -221.565 -178.255 -220.635 -177.925 ;
        RECT -229.785 -178.780 -229.615 -178.255 ;
        RECT -220.805 -178.780 -220.635 -178.255 ;
        RECT -220.395 -178.805 -220.105 -177.640 ;
        RECT -219.865 -177.925 -219.695 -177.640 ;
        RECT -210.885 -177.470 -210.715 -177.400 ;
        RECT -209.945 -177.470 -209.775 -177.400 ;
        RECT -210.885 -177.640 -209.775 -177.470 ;
        RECT -210.885 -177.925 -210.715 -177.640 ;
        RECT -219.865 -178.255 -218.935 -177.925 ;
        RECT -211.645 -178.255 -210.715 -177.925 ;
        RECT -219.865 -178.780 -219.695 -178.255 ;
        RECT -210.885 -178.780 -210.715 -178.255 ;
        RECT -210.475 -178.805 -210.185 -177.640 ;
        RECT -209.945 -177.925 -209.775 -177.640 ;
        RECT -200.965 -177.470 -200.795 -177.400 ;
        RECT -200.025 -177.470 -199.855 -177.400 ;
        RECT -200.965 -177.640 -199.855 -177.470 ;
        RECT -200.965 -177.925 -200.795 -177.640 ;
        RECT -209.945 -178.255 -209.015 -177.925 ;
        RECT -201.725 -178.255 -200.795 -177.925 ;
        RECT -209.945 -178.780 -209.775 -178.255 ;
        RECT -200.965 -178.780 -200.795 -178.255 ;
        RECT -200.555 -178.805 -200.265 -177.640 ;
        RECT -200.025 -177.925 -199.855 -177.640 ;
        RECT -191.045 -177.470 -190.875 -177.400 ;
        RECT -190.105 -177.470 -189.935 -177.400 ;
        RECT -191.045 -177.640 -189.935 -177.470 ;
        RECT -191.045 -177.925 -190.875 -177.640 ;
        RECT -200.025 -178.255 -199.095 -177.925 ;
        RECT -191.805 -178.255 -190.875 -177.925 ;
        RECT -200.025 -178.780 -199.855 -178.255 ;
        RECT -191.045 -178.780 -190.875 -178.255 ;
        RECT -190.635 -178.805 -190.345 -177.640 ;
        RECT -190.105 -177.925 -189.935 -177.640 ;
        RECT -181.125 -177.470 -180.955 -177.400 ;
        RECT -180.185 -177.470 -180.015 -177.400 ;
        RECT -181.125 -177.640 -180.015 -177.470 ;
        RECT -181.125 -177.925 -180.955 -177.640 ;
        RECT -190.105 -178.255 -189.175 -177.925 ;
        RECT -181.885 -178.255 -180.955 -177.925 ;
        RECT -190.105 -178.780 -189.935 -178.255 ;
        RECT -181.125 -178.780 -180.955 -178.255 ;
        RECT -180.715 -178.805 -180.425 -177.640 ;
        RECT -180.185 -177.925 -180.015 -177.640 ;
        RECT -171.205 -177.470 -171.035 -177.400 ;
        RECT -170.265 -177.470 -170.095 -177.400 ;
        RECT -171.205 -177.640 -170.095 -177.470 ;
        RECT -171.205 -177.925 -171.035 -177.640 ;
        RECT -180.185 -178.255 -179.255 -177.925 ;
        RECT -171.965 -178.255 -171.035 -177.925 ;
        RECT -180.185 -178.780 -180.015 -178.255 ;
        RECT -171.205 -178.780 -171.035 -178.255 ;
        RECT -170.795 -178.805 -170.505 -177.640 ;
        RECT -170.265 -177.925 -170.095 -177.640 ;
        RECT -161.285 -177.470 -161.115 -177.400 ;
        RECT -160.345 -177.470 -160.175 -177.400 ;
        RECT -161.285 -177.640 -160.175 -177.470 ;
        RECT -161.285 -177.925 -161.115 -177.640 ;
        RECT -170.265 -178.255 -169.335 -177.925 ;
        RECT -162.045 -178.255 -161.115 -177.925 ;
        RECT -170.265 -178.780 -170.095 -178.255 ;
        RECT -161.285 -178.780 -161.115 -178.255 ;
        RECT -160.875 -178.805 -160.585 -177.640 ;
        RECT -160.345 -177.925 -160.175 -177.640 ;
        RECT -151.365 -177.470 -151.195 -177.400 ;
        RECT -150.425 -177.470 -150.255 -177.400 ;
        RECT -151.365 -177.640 -150.255 -177.470 ;
        RECT -151.365 -177.925 -151.195 -177.640 ;
        RECT -160.345 -178.255 -159.415 -177.925 ;
        RECT -152.125 -178.255 -151.195 -177.925 ;
        RECT -160.345 -178.780 -160.175 -178.255 ;
        RECT -151.365 -178.780 -151.195 -178.255 ;
        RECT -150.955 -178.805 -150.665 -177.640 ;
        RECT -150.425 -177.925 -150.255 -177.640 ;
        RECT -141.445 -177.470 -141.275 -177.400 ;
        RECT -140.505 -177.470 -140.335 -177.400 ;
        RECT -141.445 -177.640 -140.335 -177.470 ;
        RECT -141.445 -177.925 -141.275 -177.640 ;
        RECT -150.425 -178.255 -149.495 -177.925 ;
        RECT -142.205 -178.255 -141.275 -177.925 ;
        RECT -150.425 -178.780 -150.255 -178.255 ;
        RECT -141.445 -178.780 -141.275 -178.255 ;
        RECT -141.035 -178.805 -140.745 -177.640 ;
        RECT -140.505 -177.925 -140.335 -177.640 ;
        RECT -131.525 -177.470 -131.355 -177.400 ;
        RECT -130.585 -177.470 -130.415 -177.400 ;
        RECT -131.525 -177.640 -130.415 -177.470 ;
        RECT -131.525 -177.925 -131.355 -177.640 ;
        RECT -140.505 -178.255 -139.575 -177.925 ;
        RECT -132.285 -178.255 -131.355 -177.925 ;
        RECT -140.505 -178.780 -140.335 -178.255 ;
        RECT -131.525 -178.780 -131.355 -178.255 ;
        RECT -131.115 -178.805 -130.825 -177.640 ;
        RECT -130.585 -177.925 -130.415 -177.640 ;
        RECT -121.605 -177.470 -121.435 -177.400 ;
        RECT -120.665 -177.470 -120.495 -177.400 ;
        RECT -121.605 -177.640 -120.495 -177.470 ;
        RECT -121.605 -177.925 -121.435 -177.640 ;
        RECT -130.585 -178.255 -129.655 -177.925 ;
        RECT -122.365 -178.255 -121.435 -177.925 ;
        RECT -130.585 -178.780 -130.415 -178.255 ;
        RECT -121.605 -178.780 -121.435 -178.255 ;
        RECT -121.195 -178.805 -120.905 -177.640 ;
        RECT -120.665 -177.925 -120.495 -177.640 ;
        RECT -111.685 -177.470 -111.515 -177.400 ;
        RECT -110.745 -177.470 -110.575 -177.400 ;
        RECT -111.685 -177.640 -110.575 -177.470 ;
        RECT -111.685 -177.925 -111.515 -177.640 ;
        RECT -120.665 -178.255 -119.735 -177.925 ;
        RECT -112.445 -178.255 -111.515 -177.925 ;
        RECT -120.665 -178.780 -120.495 -178.255 ;
        RECT -111.685 -178.780 -111.515 -178.255 ;
        RECT -111.275 -178.805 -110.985 -177.640 ;
        RECT -110.745 -177.925 -110.575 -177.640 ;
        RECT -101.765 -177.470 -101.595 -177.400 ;
        RECT -100.825 -177.470 -100.655 -177.400 ;
        RECT -101.765 -177.640 -100.655 -177.470 ;
        RECT -101.765 -177.925 -101.595 -177.640 ;
        RECT -110.745 -178.255 -109.815 -177.925 ;
        RECT -102.525 -178.255 -101.595 -177.925 ;
        RECT -110.745 -178.780 -110.575 -178.255 ;
        RECT -101.765 -178.780 -101.595 -178.255 ;
        RECT -101.355 -178.805 -101.065 -177.640 ;
        RECT -100.825 -177.925 -100.655 -177.640 ;
        RECT -91.845 -177.470 -91.675 -177.400 ;
        RECT -90.905 -177.470 -90.735 -177.400 ;
        RECT -91.845 -177.640 -90.735 -177.470 ;
        RECT -91.845 -177.925 -91.675 -177.640 ;
        RECT -100.825 -178.255 -99.895 -177.925 ;
        RECT -92.605 -178.255 -91.675 -177.925 ;
        RECT -100.825 -178.780 -100.655 -178.255 ;
        RECT -91.845 -178.780 -91.675 -178.255 ;
        RECT -91.435 -178.805 -91.145 -177.640 ;
        RECT -90.905 -177.925 -90.735 -177.640 ;
        RECT -81.925 -177.470 -81.755 -177.400 ;
        RECT -80.985 -177.470 -80.815 -177.400 ;
        RECT -81.925 -177.640 -80.815 -177.470 ;
        RECT -81.925 -177.925 -81.755 -177.640 ;
        RECT -90.905 -178.255 -89.975 -177.925 ;
        RECT -82.685 -178.255 -81.755 -177.925 ;
        RECT -90.905 -178.780 -90.735 -178.255 ;
        RECT -81.925 -178.780 -81.755 -178.255 ;
        RECT -81.515 -178.805 -81.225 -177.640 ;
        RECT -80.985 -177.925 -80.815 -177.640 ;
        RECT -72.005 -177.470 -71.835 -177.400 ;
        RECT -71.065 -177.470 -70.895 -177.400 ;
        RECT -72.005 -177.640 -70.895 -177.470 ;
        RECT -72.005 -177.925 -71.835 -177.640 ;
        RECT -80.985 -178.255 -80.055 -177.925 ;
        RECT -72.765 -178.255 -71.835 -177.925 ;
        RECT -80.985 -178.780 -80.815 -178.255 ;
        RECT -72.005 -178.780 -71.835 -178.255 ;
        RECT -71.595 -178.805 -71.305 -177.640 ;
        RECT -71.065 -177.925 -70.895 -177.640 ;
        RECT -62.085 -177.470 -61.915 -177.400 ;
        RECT -61.145 -177.470 -60.975 -177.400 ;
        RECT -62.085 -177.640 -60.975 -177.470 ;
        RECT -62.085 -177.925 -61.915 -177.640 ;
        RECT -71.065 -178.255 -70.135 -177.925 ;
        RECT -62.845 -178.255 -61.915 -177.925 ;
        RECT -71.065 -178.780 -70.895 -178.255 ;
        RECT -62.085 -178.780 -61.915 -178.255 ;
        RECT -61.675 -178.805 -61.385 -177.640 ;
        RECT -61.145 -177.925 -60.975 -177.640 ;
        RECT -52.165 -177.470 -51.995 -177.400 ;
        RECT -51.225 -177.470 -51.055 -177.400 ;
        RECT -52.165 -177.640 -51.055 -177.470 ;
        RECT -52.165 -177.925 -51.995 -177.640 ;
        RECT -61.145 -178.255 -60.215 -177.925 ;
        RECT -52.925 -178.255 -51.995 -177.925 ;
        RECT -61.145 -178.780 -60.975 -178.255 ;
        RECT -52.165 -178.780 -51.995 -178.255 ;
        RECT -51.755 -178.805 -51.465 -177.640 ;
        RECT -51.225 -177.925 -51.055 -177.640 ;
        RECT -42.245 -177.470 -42.075 -177.400 ;
        RECT -41.305 -177.470 -41.135 -177.400 ;
        RECT -42.245 -177.640 -41.135 -177.470 ;
        RECT -42.245 -177.925 -42.075 -177.640 ;
        RECT -51.225 -178.255 -50.295 -177.925 ;
        RECT -43.005 -178.255 -42.075 -177.925 ;
        RECT -51.225 -178.780 -51.055 -178.255 ;
        RECT -42.245 -178.780 -42.075 -178.255 ;
        RECT -41.835 -178.805 -41.545 -177.640 ;
        RECT -41.305 -177.925 -41.135 -177.640 ;
        RECT -32.325 -177.470 -32.155 -177.400 ;
        RECT -31.385 -177.470 -31.215 -177.400 ;
        RECT -32.325 -177.640 -31.215 -177.470 ;
        RECT -32.325 -177.925 -32.155 -177.640 ;
        RECT -41.305 -178.255 -40.375 -177.925 ;
        RECT -33.085 -178.255 -32.155 -177.925 ;
        RECT -41.305 -178.780 -41.135 -178.255 ;
        RECT -32.325 -178.780 -32.155 -178.255 ;
        RECT -31.915 -178.805 -31.625 -177.640 ;
        RECT -31.385 -177.925 -31.215 -177.640 ;
        RECT -22.405 -177.470 -22.235 -177.400 ;
        RECT -21.465 -177.470 -21.295 -177.400 ;
        RECT -22.405 -177.640 -21.295 -177.470 ;
        RECT -22.405 -177.925 -22.235 -177.640 ;
        RECT -31.385 -178.255 -30.455 -177.925 ;
        RECT -23.165 -178.255 -22.235 -177.925 ;
        RECT -31.385 -178.780 -31.215 -178.255 ;
        RECT -22.405 -178.780 -22.235 -178.255 ;
        RECT -21.995 -178.805 -21.705 -177.640 ;
        RECT -21.465 -177.925 -21.295 -177.640 ;
        RECT -12.485 -177.470 -12.315 -177.400 ;
        RECT -11.545 -177.470 -11.375 -177.400 ;
        RECT -12.485 -177.640 -11.375 -177.470 ;
        RECT -12.485 -177.925 -12.315 -177.640 ;
        RECT -21.465 -178.255 -20.535 -177.925 ;
        RECT -13.245 -178.255 -12.315 -177.925 ;
        RECT -21.465 -178.780 -21.295 -178.255 ;
        RECT -12.485 -178.780 -12.315 -178.255 ;
        RECT -12.075 -178.805 -11.785 -177.640 ;
        RECT -11.545 -177.925 -11.375 -177.640 ;
        RECT -2.565 -177.470 -2.395 -177.400 ;
        RECT -1.625 -177.470 -1.455 -177.400 ;
        RECT -2.565 -177.640 -1.455 -177.470 ;
        RECT -2.565 -177.925 -2.395 -177.640 ;
        RECT -11.545 -178.255 -10.615 -177.925 ;
        RECT -3.325 -178.255 -2.395 -177.925 ;
        RECT -11.545 -178.780 -11.375 -178.255 ;
        RECT -2.565 -178.780 -2.395 -178.255 ;
        RECT -2.155 -178.805 -1.865 -177.640 ;
        RECT -1.625 -177.925 -1.455 -177.640 ;
        RECT 7.355 -177.470 7.525 -177.400 ;
        RECT 8.295 -177.470 8.465 -177.400 ;
        RECT 7.355 -177.640 8.465 -177.470 ;
        RECT 7.355 -177.925 7.525 -177.640 ;
        RECT -1.625 -178.255 -0.695 -177.925 ;
        RECT 6.595 -178.255 7.525 -177.925 ;
        RECT -1.625 -178.780 -1.455 -178.255 ;
        RECT 7.355 -178.780 7.525 -178.255 ;
        RECT 7.765 -178.805 8.055 -177.640 ;
        RECT 8.295 -177.925 8.465 -177.640 ;
        RECT 17.275 -177.470 17.445 -177.400 ;
        RECT 18.215 -177.470 18.385 -177.400 ;
        RECT 17.275 -177.640 18.385 -177.470 ;
        RECT 17.275 -177.925 17.445 -177.640 ;
        RECT 8.295 -178.255 9.225 -177.925 ;
        RECT 16.515 -178.255 17.445 -177.925 ;
        RECT 8.295 -178.780 8.465 -178.255 ;
        RECT 17.275 -178.780 17.445 -178.255 ;
        RECT 17.685 -178.805 17.975 -177.640 ;
        RECT 18.215 -177.925 18.385 -177.640 ;
        RECT 18.215 -178.255 19.145 -177.925 ;
        RECT 18.215 -178.780 18.385 -178.255 ;
      LAYER mcon ;
        RECT -281.865 94.825 -281.695 94.995 ;
        RECT -281.395 94.820 -281.225 94.990 ;
        RECT -280.925 94.825 -280.755 94.995 ;
        RECT -281.865 94.365 -281.695 94.535 ;
        RECT -281.865 93.905 -281.695 94.075 ;
        RECT -271.945 94.825 -271.775 94.995 ;
        RECT -271.475 94.820 -271.305 94.990 ;
        RECT -271.005 94.825 -270.835 94.995 ;
        RECT -280.925 94.365 -280.755 94.535 ;
        RECT -271.945 94.365 -271.775 94.535 ;
        RECT -280.925 93.905 -280.755 94.075 ;
        RECT -271.945 93.905 -271.775 94.075 ;
        RECT -262.025 94.825 -261.855 94.995 ;
        RECT -261.555 94.820 -261.385 94.990 ;
        RECT -261.085 94.825 -260.915 94.995 ;
        RECT -271.005 94.365 -270.835 94.535 ;
        RECT -262.025 94.365 -261.855 94.535 ;
        RECT -271.005 93.905 -270.835 94.075 ;
        RECT -262.025 93.905 -261.855 94.075 ;
        RECT -252.105 94.825 -251.935 94.995 ;
        RECT -251.635 94.820 -251.465 94.990 ;
        RECT -251.165 94.825 -250.995 94.995 ;
        RECT -261.085 94.365 -260.915 94.535 ;
        RECT -252.105 94.365 -251.935 94.535 ;
        RECT -261.085 93.905 -260.915 94.075 ;
        RECT -252.105 93.905 -251.935 94.075 ;
        RECT -242.185 94.825 -242.015 94.995 ;
        RECT -241.715 94.820 -241.545 94.990 ;
        RECT -241.245 94.825 -241.075 94.995 ;
        RECT -251.165 94.365 -250.995 94.535 ;
        RECT -242.185 94.365 -242.015 94.535 ;
        RECT -251.165 93.905 -250.995 94.075 ;
        RECT -242.185 93.905 -242.015 94.075 ;
        RECT -232.265 94.825 -232.095 94.995 ;
        RECT -231.795 94.820 -231.625 94.990 ;
        RECT -231.325 94.825 -231.155 94.995 ;
        RECT -241.245 94.365 -241.075 94.535 ;
        RECT -232.265 94.365 -232.095 94.535 ;
        RECT -241.245 93.905 -241.075 94.075 ;
        RECT -232.265 93.905 -232.095 94.075 ;
        RECT -222.345 94.825 -222.175 94.995 ;
        RECT -221.875 94.820 -221.705 94.990 ;
        RECT -221.405 94.825 -221.235 94.995 ;
        RECT -231.325 94.365 -231.155 94.535 ;
        RECT -222.345 94.365 -222.175 94.535 ;
        RECT -231.325 93.905 -231.155 94.075 ;
        RECT -222.345 93.905 -222.175 94.075 ;
        RECT -212.425 94.825 -212.255 94.995 ;
        RECT -211.955 94.820 -211.785 94.990 ;
        RECT -211.485 94.825 -211.315 94.995 ;
        RECT -221.405 94.365 -221.235 94.535 ;
        RECT -212.425 94.365 -212.255 94.535 ;
        RECT -221.405 93.905 -221.235 94.075 ;
        RECT -212.425 93.905 -212.255 94.075 ;
        RECT -202.505 94.825 -202.335 94.995 ;
        RECT -202.035 94.820 -201.865 94.990 ;
        RECT -201.565 94.825 -201.395 94.995 ;
        RECT -211.485 94.365 -211.315 94.535 ;
        RECT -202.505 94.365 -202.335 94.535 ;
        RECT -211.485 93.905 -211.315 94.075 ;
        RECT -202.505 93.905 -202.335 94.075 ;
        RECT -192.585 94.825 -192.415 94.995 ;
        RECT -192.115 94.820 -191.945 94.990 ;
        RECT -191.645 94.825 -191.475 94.995 ;
        RECT -201.565 94.365 -201.395 94.535 ;
        RECT -192.585 94.365 -192.415 94.535 ;
        RECT -201.565 93.905 -201.395 94.075 ;
        RECT -192.585 93.905 -192.415 94.075 ;
        RECT -182.665 94.825 -182.495 94.995 ;
        RECT -182.195 94.820 -182.025 94.990 ;
        RECT -181.725 94.825 -181.555 94.995 ;
        RECT -191.645 94.365 -191.475 94.535 ;
        RECT -182.665 94.365 -182.495 94.535 ;
        RECT -191.645 93.905 -191.475 94.075 ;
        RECT -182.665 93.905 -182.495 94.075 ;
        RECT -172.745 94.825 -172.575 94.995 ;
        RECT -172.275 94.820 -172.105 94.990 ;
        RECT -171.805 94.825 -171.635 94.995 ;
        RECT -181.725 94.365 -181.555 94.535 ;
        RECT -172.745 94.365 -172.575 94.535 ;
        RECT -181.725 93.905 -181.555 94.075 ;
        RECT -172.745 93.905 -172.575 94.075 ;
        RECT -162.825 94.825 -162.655 94.995 ;
        RECT -162.355 94.820 -162.185 94.990 ;
        RECT -161.885 94.825 -161.715 94.995 ;
        RECT -171.805 94.365 -171.635 94.535 ;
        RECT -162.825 94.365 -162.655 94.535 ;
        RECT -171.805 93.905 -171.635 94.075 ;
        RECT -162.825 93.905 -162.655 94.075 ;
        RECT -152.905 94.825 -152.735 94.995 ;
        RECT -152.435 94.820 -152.265 94.990 ;
        RECT -151.965 94.825 -151.795 94.995 ;
        RECT -161.885 94.365 -161.715 94.535 ;
        RECT -152.905 94.365 -152.735 94.535 ;
        RECT -161.885 93.905 -161.715 94.075 ;
        RECT -152.905 93.905 -152.735 94.075 ;
        RECT -142.985 94.825 -142.815 94.995 ;
        RECT -142.515 94.820 -142.345 94.990 ;
        RECT -142.045 94.825 -141.875 94.995 ;
        RECT -151.965 94.365 -151.795 94.535 ;
        RECT -142.985 94.365 -142.815 94.535 ;
        RECT -151.965 93.905 -151.795 94.075 ;
        RECT -142.985 93.905 -142.815 94.075 ;
        RECT -133.065 94.825 -132.895 94.995 ;
        RECT -132.595 94.820 -132.425 94.990 ;
        RECT -132.125 94.825 -131.955 94.995 ;
        RECT -142.045 94.365 -141.875 94.535 ;
        RECT -133.065 94.365 -132.895 94.535 ;
        RECT -142.045 93.905 -141.875 94.075 ;
        RECT -133.065 93.905 -132.895 94.075 ;
        RECT -123.145 94.825 -122.975 94.995 ;
        RECT -122.675 94.820 -122.505 94.990 ;
        RECT -122.205 94.825 -122.035 94.995 ;
        RECT -132.125 94.365 -131.955 94.535 ;
        RECT -123.145 94.365 -122.975 94.535 ;
        RECT -132.125 93.905 -131.955 94.075 ;
        RECT -123.145 93.905 -122.975 94.075 ;
        RECT -113.225 94.825 -113.055 94.995 ;
        RECT -112.755 94.820 -112.585 94.990 ;
        RECT -112.285 94.825 -112.115 94.995 ;
        RECT -122.205 94.365 -122.035 94.535 ;
        RECT -113.225 94.365 -113.055 94.535 ;
        RECT -122.205 93.905 -122.035 94.075 ;
        RECT -113.225 93.905 -113.055 94.075 ;
        RECT -103.305 94.825 -103.135 94.995 ;
        RECT -102.835 94.820 -102.665 94.990 ;
        RECT -102.365 94.825 -102.195 94.995 ;
        RECT -112.285 94.365 -112.115 94.535 ;
        RECT -103.305 94.365 -103.135 94.535 ;
        RECT -112.285 93.905 -112.115 94.075 ;
        RECT -103.305 93.905 -103.135 94.075 ;
        RECT -93.385 94.825 -93.215 94.995 ;
        RECT -92.915 94.820 -92.745 94.990 ;
        RECT -92.445 94.825 -92.275 94.995 ;
        RECT -102.365 94.365 -102.195 94.535 ;
        RECT -93.385 94.365 -93.215 94.535 ;
        RECT -102.365 93.905 -102.195 94.075 ;
        RECT -93.385 93.905 -93.215 94.075 ;
        RECT -83.465 94.825 -83.295 94.995 ;
        RECT -82.995 94.820 -82.825 94.990 ;
        RECT -82.525 94.825 -82.355 94.995 ;
        RECT -92.445 94.365 -92.275 94.535 ;
        RECT -83.465 94.365 -83.295 94.535 ;
        RECT -92.445 93.905 -92.275 94.075 ;
        RECT -83.465 93.905 -83.295 94.075 ;
        RECT -73.545 94.825 -73.375 94.995 ;
        RECT -73.075 94.820 -72.905 94.990 ;
        RECT -72.605 94.825 -72.435 94.995 ;
        RECT -82.525 94.365 -82.355 94.535 ;
        RECT -73.545 94.365 -73.375 94.535 ;
        RECT -82.525 93.905 -82.355 94.075 ;
        RECT -73.545 93.905 -73.375 94.075 ;
        RECT -63.625 94.825 -63.455 94.995 ;
        RECT -63.155 94.820 -62.985 94.990 ;
        RECT -62.685 94.825 -62.515 94.995 ;
        RECT -72.605 94.365 -72.435 94.535 ;
        RECT -63.625 94.365 -63.455 94.535 ;
        RECT -72.605 93.905 -72.435 94.075 ;
        RECT -63.625 93.905 -63.455 94.075 ;
        RECT -53.705 94.825 -53.535 94.995 ;
        RECT -53.235 94.820 -53.065 94.990 ;
        RECT -52.765 94.825 -52.595 94.995 ;
        RECT -62.685 94.365 -62.515 94.535 ;
        RECT -53.705 94.365 -53.535 94.535 ;
        RECT -62.685 93.905 -62.515 94.075 ;
        RECT -53.705 93.905 -53.535 94.075 ;
        RECT -43.785 94.825 -43.615 94.995 ;
        RECT -43.315 94.820 -43.145 94.990 ;
        RECT -42.845 94.825 -42.675 94.995 ;
        RECT -52.765 94.365 -52.595 94.535 ;
        RECT -43.785 94.365 -43.615 94.535 ;
        RECT -52.765 93.905 -52.595 94.075 ;
        RECT -43.785 93.905 -43.615 94.075 ;
        RECT -33.865 94.825 -33.695 94.995 ;
        RECT -33.395 94.820 -33.225 94.990 ;
        RECT -32.925 94.825 -32.755 94.995 ;
        RECT -42.845 94.365 -42.675 94.535 ;
        RECT -33.865 94.365 -33.695 94.535 ;
        RECT -42.845 93.905 -42.675 94.075 ;
        RECT -33.865 93.905 -33.695 94.075 ;
        RECT -23.945 94.825 -23.775 94.995 ;
        RECT -23.475 94.820 -23.305 94.990 ;
        RECT -23.005 94.825 -22.835 94.995 ;
        RECT -32.925 94.365 -32.755 94.535 ;
        RECT -23.945 94.365 -23.775 94.535 ;
        RECT -32.925 93.905 -32.755 94.075 ;
        RECT -23.945 93.905 -23.775 94.075 ;
        RECT -14.025 94.825 -13.855 94.995 ;
        RECT -13.555 94.820 -13.385 94.990 ;
        RECT -13.085 94.825 -12.915 94.995 ;
        RECT -23.005 94.365 -22.835 94.535 ;
        RECT -14.025 94.365 -13.855 94.535 ;
        RECT -23.005 93.905 -22.835 94.075 ;
        RECT -14.025 93.905 -13.855 94.075 ;
        RECT -4.105 94.825 -3.935 94.995 ;
        RECT -3.635 94.820 -3.465 94.990 ;
        RECT -3.165 94.825 -2.995 94.995 ;
        RECT -13.085 94.365 -12.915 94.535 ;
        RECT -4.105 94.365 -3.935 94.535 ;
        RECT -13.085 93.905 -12.915 94.075 ;
        RECT -4.105 93.905 -3.935 94.075 ;
        RECT 5.815 94.825 5.985 94.995 ;
        RECT 6.285 94.820 6.455 94.990 ;
        RECT 6.755 94.825 6.925 94.995 ;
        RECT -3.165 94.365 -2.995 94.535 ;
        RECT 5.815 94.365 5.985 94.535 ;
        RECT -3.165 93.905 -2.995 94.075 ;
        RECT 5.815 93.905 5.985 94.075 ;
        RECT 15.735 94.825 15.905 94.995 ;
        RECT 16.205 94.820 16.375 94.990 ;
        RECT 16.675 94.825 16.845 94.995 ;
        RECT 6.755 94.365 6.925 94.535 ;
        RECT 15.735 94.365 15.905 94.535 ;
        RECT 6.755 93.905 6.925 94.075 ;
        RECT 15.735 93.905 15.905 94.075 ;
        RECT 25.655 94.825 25.825 94.995 ;
        RECT 26.125 94.820 26.295 94.990 ;
        RECT 16.675 94.365 16.845 94.535 ;
        RECT 25.655 94.365 25.825 94.535 ;
        RECT 16.675 93.905 16.845 94.075 ;
        RECT 25.655 93.905 25.825 94.075 ;
        RECT -287.735 93.245 -287.565 93.415 ;
        RECT -287.275 93.245 -287.105 93.415 ;
        RECT -286.815 93.245 -286.645 93.415 ;
        RECT -286.355 93.245 -286.185 93.415 ;
        RECT -285.895 93.245 -285.725 93.415 ;
        RECT -285.435 93.245 -285.265 93.415 ;
        RECT -284.975 93.245 -284.805 93.415 ;
        RECT -277.815 93.245 -277.645 93.415 ;
        RECT -277.355 93.245 -277.185 93.415 ;
        RECT -276.895 93.245 -276.725 93.415 ;
        RECT -276.435 93.245 -276.265 93.415 ;
        RECT -275.975 93.245 -275.805 93.415 ;
        RECT -275.515 93.245 -275.345 93.415 ;
        RECT -275.055 93.245 -274.885 93.415 ;
        RECT -267.895 93.245 -267.725 93.415 ;
        RECT -267.435 93.245 -267.265 93.415 ;
        RECT -266.975 93.245 -266.805 93.415 ;
        RECT -266.515 93.245 -266.345 93.415 ;
        RECT -266.055 93.245 -265.885 93.415 ;
        RECT -265.595 93.245 -265.425 93.415 ;
        RECT -265.135 93.245 -264.965 93.415 ;
        RECT -257.975 93.245 -257.805 93.415 ;
        RECT -257.515 93.245 -257.345 93.415 ;
        RECT -257.055 93.245 -256.885 93.415 ;
        RECT -256.595 93.245 -256.425 93.415 ;
        RECT -256.135 93.245 -255.965 93.415 ;
        RECT -255.675 93.245 -255.505 93.415 ;
        RECT -255.215 93.245 -255.045 93.415 ;
        RECT -248.055 93.245 -247.885 93.415 ;
        RECT -247.595 93.245 -247.425 93.415 ;
        RECT -247.135 93.245 -246.965 93.415 ;
        RECT -246.675 93.245 -246.505 93.415 ;
        RECT -246.215 93.245 -246.045 93.415 ;
        RECT -245.755 93.245 -245.585 93.415 ;
        RECT -245.295 93.245 -245.125 93.415 ;
        RECT -238.135 93.245 -237.965 93.415 ;
        RECT -237.675 93.245 -237.505 93.415 ;
        RECT -237.215 93.245 -237.045 93.415 ;
        RECT -236.755 93.245 -236.585 93.415 ;
        RECT -236.295 93.245 -236.125 93.415 ;
        RECT -235.835 93.245 -235.665 93.415 ;
        RECT -235.375 93.245 -235.205 93.415 ;
        RECT -228.215 93.245 -228.045 93.415 ;
        RECT -227.755 93.245 -227.585 93.415 ;
        RECT -227.295 93.245 -227.125 93.415 ;
        RECT -226.835 93.245 -226.665 93.415 ;
        RECT -226.375 93.245 -226.205 93.415 ;
        RECT -225.915 93.245 -225.745 93.415 ;
        RECT -225.455 93.245 -225.285 93.415 ;
        RECT -218.295 93.245 -218.125 93.415 ;
        RECT -217.835 93.245 -217.665 93.415 ;
        RECT -217.375 93.245 -217.205 93.415 ;
        RECT -216.915 93.245 -216.745 93.415 ;
        RECT -216.455 93.245 -216.285 93.415 ;
        RECT -215.995 93.245 -215.825 93.415 ;
        RECT -215.535 93.245 -215.365 93.415 ;
        RECT -208.375 93.245 -208.205 93.415 ;
        RECT -207.915 93.245 -207.745 93.415 ;
        RECT -207.455 93.245 -207.285 93.415 ;
        RECT -206.995 93.245 -206.825 93.415 ;
        RECT -206.535 93.245 -206.365 93.415 ;
        RECT -206.075 93.245 -205.905 93.415 ;
        RECT -205.615 93.245 -205.445 93.415 ;
        RECT -198.455 93.245 -198.285 93.415 ;
        RECT -197.995 93.245 -197.825 93.415 ;
        RECT -197.535 93.245 -197.365 93.415 ;
        RECT -197.075 93.245 -196.905 93.415 ;
        RECT -196.615 93.245 -196.445 93.415 ;
        RECT -196.155 93.245 -195.985 93.415 ;
        RECT -195.695 93.245 -195.525 93.415 ;
        RECT -188.535 93.245 -188.365 93.415 ;
        RECT -188.075 93.245 -187.905 93.415 ;
        RECT -187.615 93.245 -187.445 93.415 ;
        RECT -187.155 93.245 -186.985 93.415 ;
        RECT -186.695 93.245 -186.525 93.415 ;
        RECT -186.235 93.245 -186.065 93.415 ;
        RECT -185.775 93.245 -185.605 93.415 ;
        RECT -178.615 93.245 -178.445 93.415 ;
        RECT -178.155 93.245 -177.985 93.415 ;
        RECT -177.695 93.245 -177.525 93.415 ;
        RECT -177.235 93.245 -177.065 93.415 ;
        RECT -176.775 93.245 -176.605 93.415 ;
        RECT -176.315 93.245 -176.145 93.415 ;
        RECT -175.855 93.245 -175.685 93.415 ;
        RECT -168.695 93.245 -168.525 93.415 ;
        RECT -168.235 93.245 -168.065 93.415 ;
        RECT -167.775 93.245 -167.605 93.415 ;
        RECT -167.315 93.245 -167.145 93.415 ;
        RECT -166.855 93.245 -166.685 93.415 ;
        RECT -166.395 93.245 -166.225 93.415 ;
        RECT -165.935 93.245 -165.765 93.415 ;
        RECT -158.775 93.245 -158.605 93.415 ;
        RECT -158.315 93.245 -158.145 93.415 ;
        RECT -157.855 93.245 -157.685 93.415 ;
        RECT -157.395 93.245 -157.225 93.415 ;
        RECT -156.935 93.245 -156.765 93.415 ;
        RECT -156.475 93.245 -156.305 93.415 ;
        RECT -156.015 93.245 -155.845 93.415 ;
        RECT -148.855 93.245 -148.685 93.415 ;
        RECT -148.395 93.245 -148.225 93.415 ;
        RECT -147.935 93.245 -147.765 93.415 ;
        RECT -147.475 93.245 -147.305 93.415 ;
        RECT -147.015 93.245 -146.845 93.415 ;
        RECT -146.555 93.245 -146.385 93.415 ;
        RECT -146.095 93.245 -145.925 93.415 ;
        RECT -138.935 93.245 -138.765 93.415 ;
        RECT -138.475 93.245 -138.305 93.415 ;
        RECT -138.015 93.245 -137.845 93.415 ;
        RECT -137.555 93.245 -137.385 93.415 ;
        RECT -137.095 93.245 -136.925 93.415 ;
        RECT -136.635 93.245 -136.465 93.415 ;
        RECT -136.175 93.245 -136.005 93.415 ;
        RECT -129.015 93.245 -128.845 93.415 ;
        RECT -128.555 93.245 -128.385 93.415 ;
        RECT -128.095 93.245 -127.925 93.415 ;
        RECT -127.635 93.245 -127.465 93.415 ;
        RECT -127.175 93.245 -127.005 93.415 ;
        RECT -126.715 93.245 -126.545 93.415 ;
        RECT -126.255 93.245 -126.085 93.415 ;
        RECT -119.095 93.245 -118.925 93.415 ;
        RECT -118.635 93.245 -118.465 93.415 ;
        RECT -118.175 93.245 -118.005 93.415 ;
        RECT -117.715 93.245 -117.545 93.415 ;
        RECT -117.255 93.245 -117.085 93.415 ;
        RECT -116.795 93.245 -116.625 93.415 ;
        RECT -116.335 93.245 -116.165 93.415 ;
        RECT -109.175 93.245 -109.005 93.415 ;
        RECT -108.715 93.245 -108.545 93.415 ;
        RECT -108.255 93.245 -108.085 93.415 ;
        RECT -107.795 93.245 -107.625 93.415 ;
        RECT -107.335 93.245 -107.165 93.415 ;
        RECT -106.875 93.245 -106.705 93.415 ;
        RECT -106.415 93.245 -106.245 93.415 ;
        RECT -99.255 93.245 -99.085 93.415 ;
        RECT -98.795 93.245 -98.625 93.415 ;
        RECT -98.335 93.245 -98.165 93.415 ;
        RECT -97.875 93.245 -97.705 93.415 ;
        RECT -97.415 93.245 -97.245 93.415 ;
        RECT -96.955 93.245 -96.785 93.415 ;
        RECT -96.495 93.245 -96.325 93.415 ;
        RECT -89.335 93.245 -89.165 93.415 ;
        RECT -88.875 93.245 -88.705 93.415 ;
        RECT -88.415 93.245 -88.245 93.415 ;
        RECT -87.955 93.245 -87.785 93.415 ;
        RECT -87.495 93.245 -87.325 93.415 ;
        RECT -87.035 93.245 -86.865 93.415 ;
        RECT -86.575 93.245 -86.405 93.415 ;
        RECT -79.415 93.245 -79.245 93.415 ;
        RECT -78.955 93.245 -78.785 93.415 ;
        RECT -78.495 93.245 -78.325 93.415 ;
        RECT -78.035 93.245 -77.865 93.415 ;
        RECT -77.575 93.245 -77.405 93.415 ;
        RECT -77.115 93.245 -76.945 93.415 ;
        RECT -76.655 93.245 -76.485 93.415 ;
        RECT -69.495 93.245 -69.325 93.415 ;
        RECT -69.035 93.245 -68.865 93.415 ;
        RECT -68.575 93.245 -68.405 93.415 ;
        RECT -68.115 93.245 -67.945 93.415 ;
        RECT -67.655 93.245 -67.485 93.415 ;
        RECT -67.195 93.245 -67.025 93.415 ;
        RECT -66.735 93.245 -66.565 93.415 ;
        RECT -59.575 93.245 -59.405 93.415 ;
        RECT -59.115 93.245 -58.945 93.415 ;
        RECT -58.655 93.245 -58.485 93.415 ;
        RECT -58.195 93.245 -58.025 93.415 ;
        RECT -57.735 93.245 -57.565 93.415 ;
        RECT -57.275 93.245 -57.105 93.415 ;
        RECT -56.815 93.245 -56.645 93.415 ;
        RECT -49.655 93.245 -49.485 93.415 ;
        RECT -49.195 93.245 -49.025 93.415 ;
        RECT -48.735 93.245 -48.565 93.415 ;
        RECT -48.275 93.245 -48.105 93.415 ;
        RECT -47.815 93.245 -47.645 93.415 ;
        RECT -47.355 93.245 -47.185 93.415 ;
        RECT -46.895 93.245 -46.725 93.415 ;
        RECT -39.735 93.245 -39.565 93.415 ;
        RECT -39.275 93.245 -39.105 93.415 ;
        RECT -38.815 93.245 -38.645 93.415 ;
        RECT -38.355 93.245 -38.185 93.415 ;
        RECT -37.895 93.245 -37.725 93.415 ;
        RECT -37.435 93.245 -37.265 93.415 ;
        RECT -36.975 93.245 -36.805 93.415 ;
        RECT -29.815 93.245 -29.645 93.415 ;
        RECT -29.355 93.245 -29.185 93.415 ;
        RECT -28.895 93.245 -28.725 93.415 ;
        RECT -28.435 93.245 -28.265 93.415 ;
        RECT -27.975 93.245 -27.805 93.415 ;
        RECT -27.515 93.245 -27.345 93.415 ;
        RECT -27.055 93.245 -26.885 93.415 ;
        RECT -19.895 93.245 -19.725 93.415 ;
        RECT -19.435 93.245 -19.265 93.415 ;
        RECT -18.975 93.245 -18.805 93.415 ;
        RECT -18.515 93.245 -18.345 93.415 ;
        RECT -18.055 93.245 -17.885 93.415 ;
        RECT -17.595 93.245 -17.425 93.415 ;
        RECT -17.135 93.245 -16.965 93.415 ;
        RECT -9.975 93.245 -9.805 93.415 ;
        RECT -9.515 93.245 -9.345 93.415 ;
        RECT -9.055 93.245 -8.885 93.415 ;
        RECT -8.595 93.245 -8.425 93.415 ;
        RECT -8.135 93.245 -7.965 93.415 ;
        RECT -7.675 93.245 -7.505 93.415 ;
        RECT -7.215 93.245 -7.045 93.415 ;
        RECT -0.055 93.245 0.115 93.415 ;
        RECT 0.405 93.245 0.575 93.415 ;
        RECT 0.865 93.245 1.035 93.415 ;
        RECT 1.325 93.245 1.495 93.415 ;
        RECT 1.785 93.245 1.955 93.415 ;
        RECT 2.245 93.245 2.415 93.415 ;
        RECT 2.705 93.245 2.875 93.415 ;
        RECT 9.865 93.245 10.035 93.415 ;
        RECT 10.325 93.245 10.495 93.415 ;
        RECT 10.785 93.245 10.955 93.415 ;
        RECT 11.245 93.245 11.415 93.415 ;
        RECT 11.705 93.245 11.875 93.415 ;
        RECT 12.165 93.245 12.335 93.415 ;
        RECT 12.625 93.245 12.795 93.415 ;
        RECT 19.785 93.245 19.955 93.415 ;
        RECT 20.245 93.245 20.415 93.415 ;
        RECT 20.705 93.245 20.875 93.415 ;
        RECT 21.165 93.245 21.335 93.415 ;
        RECT 21.625 93.245 21.795 93.415 ;
        RECT 22.085 93.245 22.255 93.415 ;
        RECT 22.545 93.245 22.715 93.415 ;
        RECT -282.775 90.525 -282.605 90.695 ;
        RECT -282.315 90.525 -282.145 90.695 ;
        RECT -281.855 90.525 -281.685 90.695 ;
        RECT -281.395 90.525 -281.225 90.695 ;
        RECT -280.935 90.525 -280.765 90.695 ;
        RECT -280.475 90.525 -280.305 90.695 ;
        RECT -280.015 90.525 -279.845 90.695 ;
        RECT -272.855 90.525 -272.685 90.695 ;
        RECT -272.395 90.525 -272.225 90.695 ;
        RECT -271.935 90.525 -271.765 90.695 ;
        RECT -271.475 90.525 -271.305 90.695 ;
        RECT -271.015 90.525 -270.845 90.695 ;
        RECT -270.555 90.525 -270.385 90.695 ;
        RECT -270.095 90.525 -269.925 90.695 ;
        RECT -262.935 90.525 -262.765 90.695 ;
        RECT -262.475 90.525 -262.305 90.695 ;
        RECT -262.015 90.525 -261.845 90.695 ;
        RECT -261.555 90.525 -261.385 90.695 ;
        RECT -261.095 90.525 -260.925 90.695 ;
        RECT -260.635 90.525 -260.465 90.695 ;
        RECT -260.175 90.525 -260.005 90.695 ;
        RECT -253.015 90.525 -252.845 90.695 ;
        RECT -252.555 90.525 -252.385 90.695 ;
        RECT -252.095 90.525 -251.925 90.695 ;
        RECT -251.635 90.525 -251.465 90.695 ;
        RECT -251.175 90.525 -251.005 90.695 ;
        RECT -250.715 90.525 -250.545 90.695 ;
        RECT -250.255 90.525 -250.085 90.695 ;
        RECT -243.095 90.525 -242.925 90.695 ;
        RECT -242.635 90.525 -242.465 90.695 ;
        RECT -242.175 90.525 -242.005 90.695 ;
        RECT -241.715 90.525 -241.545 90.695 ;
        RECT -241.255 90.525 -241.085 90.695 ;
        RECT -240.795 90.525 -240.625 90.695 ;
        RECT -240.335 90.525 -240.165 90.695 ;
        RECT -233.175 90.525 -233.005 90.695 ;
        RECT -232.715 90.525 -232.545 90.695 ;
        RECT -232.255 90.525 -232.085 90.695 ;
        RECT -231.795 90.525 -231.625 90.695 ;
        RECT -231.335 90.525 -231.165 90.695 ;
        RECT -230.875 90.525 -230.705 90.695 ;
        RECT -230.415 90.525 -230.245 90.695 ;
        RECT -223.255 90.525 -223.085 90.695 ;
        RECT -222.795 90.525 -222.625 90.695 ;
        RECT -222.335 90.525 -222.165 90.695 ;
        RECT -221.875 90.525 -221.705 90.695 ;
        RECT -221.415 90.525 -221.245 90.695 ;
        RECT -220.955 90.525 -220.785 90.695 ;
        RECT -220.495 90.525 -220.325 90.695 ;
        RECT -213.335 90.525 -213.165 90.695 ;
        RECT -212.875 90.525 -212.705 90.695 ;
        RECT -212.415 90.525 -212.245 90.695 ;
        RECT -211.955 90.525 -211.785 90.695 ;
        RECT -211.495 90.525 -211.325 90.695 ;
        RECT -211.035 90.525 -210.865 90.695 ;
        RECT -210.575 90.525 -210.405 90.695 ;
        RECT -203.415 90.525 -203.245 90.695 ;
        RECT -202.955 90.525 -202.785 90.695 ;
        RECT -202.495 90.525 -202.325 90.695 ;
        RECT -202.035 90.525 -201.865 90.695 ;
        RECT -201.575 90.525 -201.405 90.695 ;
        RECT -201.115 90.525 -200.945 90.695 ;
        RECT -200.655 90.525 -200.485 90.695 ;
        RECT -193.495 90.525 -193.325 90.695 ;
        RECT -193.035 90.525 -192.865 90.695 ;
        RECT -192.575 90.525 -192.405 90.695 ;
        RECT -192.115 90.525 -191.945 90.695 ;
        RECT -191.655 90.525 -191.485 90.695 ;
        RECT -191.195 90.525 -191.025 90.695 ;
        RECT -190.735 90.525 -190.565 90.695 ;
        RECT -183.575 90.525 -183.405 90.695 ;
        RECT -183.115 90.525 -182.945 90.695 ;
        RECT -182.655 90.525 -182.485 90.695 ;
        RECT -182.195 90.525 -182.025 90.695 ;
        RECT -181.735 90.525 -181.565 90.695 ;
        RECT -181.275 90.525 -181.105 90.695 ;
        RECT -180.815 90.525 -180.645 90.695 ;
        RECT -173.655 90.525 -173.485 90.695 ;
        RECT -173.195 90.525 -173.025 90.695 ;
        RECT -172.735 90.525 -172.565 90.695 ;
        RECT -172.275 90.525 -172.105 90.695 ;
        RECT -171.815 90.525 -171.645 90.695 ;
        RECT -171.355 90.525 -171.185 90.695 ;
        RECT -170.895 90.525 -170.725 90.695 ;
        RECT -163.735 90.525 -163.565 90.695 ;
        RECT -163.275 90.525 -163.105 90.695 ;
        RECT -162.815 90.525 -162.645 90.695 ;
        RECT -162.355 90.525 -162.185 90.695 ;
        RECT -161.895 90.525 -161.725 90.695 ;
        RECT -161.435 90.525 -161.265 90.695 ;
        RECT -160.975 90.525 -160.805 90.695 ;
        RECT -153.815 90.525 -153.645 90.695 ;
        RECT -153.355 90.525 -153.185 90.695 ;
        RECT -152.895 90.525 -152.725 90.695 ;
        RECT -152.435 90.525 -152.265 90.695 ;
        RECT -151.975 90.525 -151.805 90.695 ;
        RECT -151.515 90.525 -151.345 90.695 ;
        RECT -151.055 90.525 -150.885 90.695 ;
        RECT -143.895 90.525 -143.725 90.695 ;
        RECT -143.435 90.525 -143.265 90.695 ;
        RECT -142.975 90.525 -142.805 90.695 ;
        RECT -142.515 90.525 -142.345 90.695 ;
        RECT -142.055 90.525 -141.885 90.695 ;
        RECT -141.595 90.525 -141.425 90.695 ;
        RECT -141.135 90.525 -140.965 90.695 ;
        RECT -133.975 90.525 -133.805 90.695 ;
        RECT -133.515 90.525 -133.345 90.695 ;
        RECT -133.055 90.525 -132.885 90.695 ;
        RECT -132.595 90.525 -132.425 90.695 ;
        RECT -132.135 90.525 -131.965 90.695 ;
        RECT -131.675 90.525 -131.505 90.695 ;
        RECT -131.215 90.525 -131.045 90.695 ;
        RECT -124.055 90.525 -123.885 90.695 ;
        RECT -123.595 90.525 -123.425 90.695 ;
        RECT -123.135 90.525 -122.965 90.695 ;
        RECT -122.675 90.525 -122.505 90.695 ;
        RECT -122.215 90.525 -122.045 90.695 ;
        RECT -121.755 90.525 -121.585 90.695 ;
        RECT -121.295 90.525 -121.125 90.695 ;
        RECT -114.135 90.525 -113.965 90.695 ;
        RECT -113.675 90.525 -113.505 90.695 ;
        RECT -113.215 90.525 -113.045 90.695 ;
        RECT -112.755 90.525 -112.585 90.695 ;
        RECT -112.295 90.525 -112.125 90.695 ;
        RECT -111.835 90.525 -111.665 90.695 ;
        RECT -111.375 90.525 -111.205 90.695 ;
        RECT -104.215 90.525 -104.045 90.695 ;
        RECT -103.755 90.525 -103.585 90.695 ;
        RECT -103.295 90.525 -103.125 90.695 ;
        RECT -102.835 90.525 -102.665 90.695 ;
        RECT -102.375 90.525 -102.205 90.695 ;
        RECT -101.915 90.525 -101.745 90.695 ;
        RECT -101.455 90.525 -101.285 90.695 ;
        RECT -94.295 90.525 -94.125 90.695 ;
        RECT -93.835 90.525 -93.665 90.695 ;
        RECT -93.375 90.525 -93.205 90.695 ;
        RECT -92.915 90.525 -92.745 90.695 ;
        RECT -92.455 90.525 -92.285 90.695 ;
        RECT -91.995 90.525 -91.825 90.695 ;
        RECT -91.535 90.525 -91.365 90.695 ;
        RECT -84.375 90.525 -84.205 90.695 ;
        RECT -83.915 90.525 -83.745 90.695 ;
        RECT -83.455 90.525 -83.285 90.695 ;
        RECT -82.995 90.525 -82.825 90.695 ;
        RECT -82.535 90.525 -82.365 90.695 ;
        RECT -82.075 90.525 -81.905 90.695 ;
        RECT -81.615 90.525 -81.445 90.695 ;
        RECT -74.455 90.525 -74.285 90.695 ;
        RECT -73.995 90.525 -73.825 90.695 ;
        RECT -73.535 90.525 -73.365 90.695 ;
        RECT -73.075 90.525 -72.905 90.695 ;
        RECT -72.615 90.525 -72.445 90.695 ;
        RECT -72.155 90.525 -71.985 90.695 ;
        RECT -71.695 90.525 -71.525 90.695 ;
        RECT -64.535 90.525 -64.365 90.695 ;
        RECT -64.075 90.525 -63.905 90.695 ;
        RECT -63.615 90.525 -63.445 90.695 ;
        RECT -63.155 90.525 -62.985 90.695 ;
        RECT -62.695 90.525 -62.525 90.695 ;
        RECT -62.235 90.525 -62.065 90.695 ;
        RECT -61.775 90.525 -61.605 90.695 ;
        RECT -54.615 90.525 -54.445 90.695 ;
        RECT -54.155 90.525 -53.985 90.695 ;
        RECT -53.695 90.525 -53.525 90.695 ;
        RECT -53.235 90.525 -53.065 90.695 ;
        RECT -52.775 90.525 -52.605 90.695 ;
        RECT -52.315 90.525 -52.145 90.695 ;
        RECT -51.855 90.525 -51.685 90.695 ;
        RECT -44.695 90.525 -44.525 90.695 ;
        RECT -44.235 90.525 -44.065 90.695 ;
        RECT -43.775 90.525 -43.605 90.695 ;
        RECT -43.315 90.525 -43.145 90.695 ;
        RECT -42.855 90.525 -42.685 90.695 ;
        RECT -42.395 90.525 -42.225 90.695 ;
        RECT -41.935 90.525 -41.765 90.695 ;
        RECT -34.775 90.525 -34.605 90.695 ;
        RECT -34.315 90.525 -34.145 90.695 ;
        RECT -33.855 90.525 -33.685 90.695 ;
        RECT -33.395 90.525 -33.225 90.695 ;
        RECT -32.935 90.525 -32.765 90.695 ;
        RECT -32.475 90.525 -32.305 90.695 ;
        RECT -32.015 90.525 -31.845 90.695 ;
        RECT -24.855 90.525 -24.685 90.695 ;
        RECT -24.395 90.525 -24.225 90.695 ;
        RECT -23.935 90.525 -23.765 90.695 ;
        RECT -23.475 90.525 -23.305 90.695 ;
        RECT -23.015 90.525 -22.845 90.695 ;
        RECT -22.555 90.525 -22.385 90.695 ;
        RECT -22.095 90.525 -21.925 90.695 ;
        RECT -14.935 90.525 -14.765 90.695 ;
        RECT -14.475 90.525 -14.305 90.695 ;
        RECT -14.015 90.525 -13.845 90.695 ;
        RECT -13.555 90.525 -13.385 90.695 ;
        RECT -13.095 90.525 -12.925 90.695 ;
        RECT -12.635 90.525 -12.465 90.695 ;
        RECT -12.175 90.525 -12.005 90.695 ;
        RECT -5.015 90.525 -4.845 90.695 ;
        RECT -4.555 90.525 -4.385 90.695 ;
        RECT -4.095 90.525 -3.925 90.695 ;
        RECT -3.635 90.525 -3.465 90.695 ;
        RECT -3.175 90.525 -3.005 90.695 ;
        RECT -2.715 90.525 -2.545 90.695 ;
        RECT -2.255 90.525 -2.085 90.695 ;
        RECT 4.905 90.525 5.075 90.695 ;
        RECT 5.365 90.525 5.535 90.695 ;
        RECT 5.825 90.525 5.995 90.695 ;
        RECT 6.285 90.525 6.455 90.695 ;
        RECT 6.745 90.525 6.915 90.695 ;
        RECT 7.205 90.525 7.375 90.695 ;
        RECT 7.665 90.525 7.835 90.695 ;
        RECT 14.825 90.525 14.995 90.695 ;
        RECT 15.285 90.525 15.455 90.695 ;
        RECT 15.745 90.525 15.915 90.695 ;
        RECT 16.205 90.525 16.375 90.695 ;
        RECT 16.665 90.525 16.835 90.695 ;
        RECT 17.125 90.525 17.295 90.695 ;
        RECT 17.585 90.525 17.755 90.695 ;
        RECT 24.745 90.525 24.915 90.695 ;
        RECT 25.205 90.525 25.375 90.695 ;
        RECT 25.665 90.525 25.835 90.695 ;
        RECT 26.125 90.525 26.295 90.695 ;
        RECT -286.825 89.865 -286.655 90.035 ;
        RECT -286.355 89.940 -286.185 90.110 ;
        RECT -286.825 89.405 -286.655 89.575 ;
        RECT -286.825 88.945 -286.655 89.115 ;
        RECT -285.885 89.865 -285.715 90.035 ;
        RECT -276.905 89.865 -276.735 90.035 ;
        RECT -276.435 89.940 -276.265 90.110 ;
        RECT -285.885 89.405 -285.715 89.575 ;
        RECT -276.905 89.405 -276.735 89.575 ;
        RECT -285.885 88.945 -285.715 89.115 ;
        RECT -276.905 88.945 -276.735 89.115 ;
        RECT -275.965 89.865 -275.795 90.035 ;
        RECT -266.985 89.865 -266.815 90.035 ;
        RECT -266.515 89.940 -266.345 90.110 ;
        RECT -275.965 89.405 -275.795 89.575 ;
        RECT -266.985 89.405 -266.815 89.575 ;
        RECT -275.965 88.945 -275.795 89.115 ;
        RECT -266.985 88.945 -266.815 89.115 ;
        RECT -266.045 89.865 -265.875 90.035 ;
        RECT -257.065 89.865 -256.895 90.035 ;
        RECT -256.595 89.940 -256.425 90.110 ;
        RECT -266.045 89.405 -265.875 89.575 ;
        RECT -257.065 89.405 -256.895 89.575 ;
        RECT -266.045 88.945 -265.875 89.115 ;
        RECT -257.065 88.945 -256.895 89.115 ;
        RECT -256.125 89.865 -255.955 90.035 ;
        RECT -247.145 89.865 -246.975 90.035 ;
        RECT -246.675 89.940 -246.505 90.110 ;
        RECT -256.125 89.405 -255.955 89.575 ;
        RECT -247.145 89.405 -246.975 89.575 ;
        RECT -256.125 88.945 -255.955 89.115 ;
        RECT -247.145 88.945 -246.975 89.115 ;
        RECT -246.205 89.865 -246.035 90.035 ;
        RECT -237.225 89.865 -237.055 90.035 ;
        RECT -236.755 89.940 -236.585 90.110 ;
        RECT -246.205 89.405 -246.035 89.575 ;
        RECT -237.225 89.405 -237.055 89.575 ;
        RECT -246.205 88.945 -246.035 89.115 ;
        RECT -237.225 88.945 -237.055 89.115 ;
        RECT -236.285 89.865 -236.115 90.035 ;
        RECT -227.305 89.865 -227.135 90.035 ;
        RECT -226.835 89.940 -226.665 90.110 ;
        RECT -236.285 89.405 -236.115 89.575 ;
        RECT -227.305 89.405 -227.135 89.575 ;
        RECT -236.285 88.945 -236.115 89.115 ;
        RECT -227.305 88.945 -227.135 89.115 ;
        RECT -226.365 89.865 -226.195 90.035 ;
        RECT -217.385 89.865 -217.215 90.035 ;
        RECT -216.915 89.940 -216.745 90.110 ;
        RECT -226.365 89.405 -226.195 89.575 ;
        RECT -217.385 89.405 -217.215 89.575 ;
        RECT -226.365 88.945 -226.195 89.115 ;
        RECT -217.385 88.945 -217.215 89.115 ;
        RECT -216.445 89.865 -216.275 90.035 ;
        RECT -207.465 89.865 -207.295 90.035 ;
        RECT -206.995 89.940 -206.825 90.110 ;
        RECT -216.445 89.405 -216.275 89.575 ;
        RECT -207.465 89.405 -207.295 89.575 ;
        RECT -216.445 88.945 -216.275 89.115 ;
        RECT -207.465 88.945 -207.295 89.115 ;
        RECT -206.525 89.865 -206.355 90.035 ;
        RECT -197.545 89.865 -197.375 90.035 ;
        RECT -197.075 89.940 -196.905 90.110 ;
        RECT -206.525 89.405 -206.355 89.575 ;
        RECT -197.545 89.405 -197.375 89.575 ;
        RECT -206.525 88.945 -206.355 89.115 ;
        RECT -197.545 88.945 -197.375 89.115 ;
        RECT -196.605 89.865 -196.435 90.035 ;
        RECT -187.625 89.865 -187.455 90.035 ;
        RECT -187.155 89.940 -186.985 90.110 ;
        RECT -196.605 89.405 -196.435 89.575 ;
        RECT -187.625 89.405 -187.455 89.575 ;
        RECT -196.605 88.945 -196.435 89.115 ;
        RECT -187.625 88.945 -187.455 89.115 ;
        RECT -186.685 89.865 -186.515 90.035 ;
        RECT -177.705 89.865 -177.535 90.035 ;
        RECT -177.235 89.940 -177.065 90.110 ;
        RECT -186.685 89.405 -186.515 89.575 ;
        RECT -177.705 89.405 -177.535 89.575 ;
        RECT -186.685 88.945 -186.515 89.115 ;
        RECT -177.705 88.945 -177.535 89.115 ;
        RECT -176.765 89.865 -176.595 90.035 ;
        RECT -167.785 89.865 -167.615 90.035 ;
        RECT -167.315 89.940 -167.145 90.110 ;
        RECT -176.765 89.405 -176.595 89.575 ;
        RECT -167.785 89.405 -167.615 89.575 ;
        RECT -176.765 88.945 -176.595 89.115 ;
        RECT -167.785 88.945 -167.615 89.115 ;
        RECT -166.845 89.865 -166.675 90.035 ;
        RECT -157.865 89.865 -157.695 90.035 ;
        RECT -157.395 89.940 -157.225 90.110 ;
        RECT -166.845 89.405 -166.675 89.575 ;
        RECT -157.865 89.405 -157.695 89.575 ;
        RECT -166.845 88.945 -166.675 89.115 ;
        RECT -157.865 88.945 -157.695 89.115 ;
        RECT -156.925 89.865 -156.755 90.035 ;
        RECT -147.945 89.865 -147.775 90.035 ;
        RECT -147.475 89.940 -147.305 90.110 ;
        RECT -156.925 89.405 -156.755 89.575 ;
        RECT -147.945 89.405 -147.775 89.575 ;
        RECT -156.925 88.945 -156.755 89.115 ;
        RECT -147.945 88.945 -147.775 89.115 ;
        RECT -147.005 89.865 -146.835 90.035 ;
        RECT -138.025 89.865 -137.855 90.035 ;
        RECT -137.555 89.940 -137.385 90.110 ;
        RECT -147.005 89.405 -146.835 89.575 ;
        RECT -138.025 89.405 -137.855 89.575 ;
        RECT -147.005 88.945 -146.835 89.115 ;
        RECT -138.025 88.945 -137.855 89.115 ;
        RECT -137.085 89.865 -136.915 90.035 ;
        RECT -128.105 89.865 -127.935 90.035 ;
        RECT -127.635 89.940 -127.465 90.110 ;
        RECT -137.085 89.405 -136.915 89.575 ;
        RECT -128.105 89.405 -127.935 89.575 ;
        RECT -137.085 88.945 -136.915 89.115 ;
        RECT -128.105 88.945 -127.935 89.115 ;
        RECT -127.165 89.865 -126.995 90.035 ;
        RECT -118.185 89.865 -118.015 90.035 ;
        RECT -117.715 89.940 -117.545 90.110 ;
        RECT -127.165 89.405 -126.995 89.575 ;
        RECT -118.185 89.405 -118.015 89.575 ;
        RECT -127.165 88.945 -126.995 89.115 ;
        RECT -118.185 88.945 -118.015 89.115 ;
        RECT -117.245 89.865 -117.075 90.035 ;
        RECT -108.265 89.865 -108.095 90.035 ;
        RECT -107.795 89.940 -107.625 90.110 ;
        RECT -117.245 89.405 -117.075 89.575 ;
        RECT -108.265 89.405 -108.095 89.575 ;
        RECT -117.245 88.945 -117.075 89.115 ;
        RECT -108.265 88.945 -108.095 89.115 ;
        RECT -107.325 89.865 -107.155 90.035 ;
        RECT -98.345 89.865 -98.175 90.035 ;
        RECT -97.875 89.940 -97.705 90.110 ;
        RECT -107.325 89.405 -107.155 89.575 ;
        RECT -98.345 89.405 -98.175 89.575 ;
        RECT -107.325 88.945 -107.155 89.115 ;
        RECT -98.345 88.945 -98.175 89.115 ;
        RECT -97.405 89.865 -97.235 90.035 ;
        RECT -88.425 89.865 -88.255 90.035 ;
        RECT -87.955 89.940 -87.785 90.110 ;
        RECT -97.405 89.405 -97.235 89.575 ;
        RECT -88.425 89.405 -88.255 89.575 ;
        RECT -97.405 88.945 -97.235 89.115 ;
        RECT -88.425 88.945 -88.255 89.115 ;
        RECT -87.485 89.865 -87.315 90.035 ;
        RECT -78.505 89.865 -78.335 90.035 ;
        RECT -78.035 89.940 -77.865 90.110 ;
        RECT -87.485 89.405 -87.315 89.575 ;
        RECT -78.505 89.405 -78.335 89.575 ;
        RECT -87.485 88.945 -87.315 89.115 ;
        RECT -78.505 88.945 -78.335 89.115 ;
        RECT -77.565 89.865 -77.395 90.035 ;
        RECT -68.585 89.865 -68.415 90.035 ;
        RECT -68.115 89.940 -67.945 90.110 ;
        RECT -77.565 89.405 -77.395 89.575 ;
        RECT -68.585 89.405 -68.415 89.575 ;
        RECT -77.565 88.945 -77.395 89.115 ;
        RECT -68.585 88.945 -68.415 89.115 ;
        RECT -67.645 89.865 -67.475 90.035 ;
        RECT -58.665 89.865 -58.495 90.035 ;
        RECT -58.195 89.940 -58.025 90.110 ;
        RECT -67.645 89.405 -67.475 89.575 ;
        RECT -58.665 89.405 -58.495 89.575 ;
        RECT -67.645 88.945 -67.475 89.115 ;
        RECT -58.665 88.945 -58.495 89.115 ;
        RECT -57.725 89.865 -57.555 90.035 ;
        RECT -48.745 89.865 -48.575 90.035 ;
        RECT -48.275 89.940 -48.105 90.110 ;
        RECT -57.725 89.405 -57.555 89.575 ;
        RECT -48.745 89.405 -48.575 89.575 ;
        RECT -57.725 88.945 -57.555 89.115 ;
        RECT -48.745 88.945 -48.575 89.115 ;
        RECT -47.805 89.865 -47.635 90.035 ;
        RECT -38.825 89.865 -38.655 90.035 ;
        RECT -38.355 89.940 -38.185 90.110 ;
        RECT -47.805 89.405 -47.635 89.575 ;
        RECT -38.825 89.405 -38.655 89.575 ;
        RECT -47.805 88.945 -47.635 89.115 ;
        RECT -38.825 88.945 -38.655 89.115 ;
        RECT -37.885 89.865 -37.715 90.035 ;
        RECT -28.905 89.865 -28.735 90.035 ;
        RECT -28.435 89.940 -28.265 90.110 ;
        RECT -37.885 89.405 -37.715 89.575 ;
        RECT -28.905 89.405 -28.735 89.575 ;
        RECT -37.885 88.945 -37.715 89.115 ;
        RECT -28.905 88.945 -28.735 89.115 ;
        RECT -27.965 89.865 -27.795 90.035 ;
        RECT -18.985 89.865 -18.815 90.035 ;
        RECT -18.515 89.940 -18.345 90.110 ;
        RECT -27.965 89.405 -27.795 89.575 ;
        RECT -18.985 89.405 -18.815 89.575 ;
        RECT -27.965 88.945 -27.795 89.115 ;
        RECT -18.985 88.945 -18.815 89.115 ;
        RECT -18.045 89.865 -17.875 90.035 ;
        RECT -9.065 89.865 -8.895 90.035 ;
        RECT -8.595 89.940 -8.425 90.110 ;
        RECT -18.045 89.405 -17.875 89.575 ;
        RECT -9.065 89.405 -8.895 89.575 ;
        RECT -18.045 88.945 -17.875 89.115 ;
        RECT -9.065 88.945 -8.895 89.115 ;
        RECT -8.125 89.865 -7.955 90.035 ;
        RECT 0.855 89.865 1.025 90.035 ;
        RECT 1.325 89.940 1.495 90.110 ;
        RECT -8.125 89.405 -7.955 89.575 ;
        RECT 0.855 89.405 1.025 89.575 ;
        RECT -8.125 88.945 -7.955 89.115 ;
        RECT 0.855 88.945 1.025 89.115 ;
        RECT 1.795 89.865 1.965 90.035 ;
        RECT 10.775 89.865 10.945 90.035 ;
        RECT 11.245 89.940 11.415 90.110 ;
        RECT 1.795 89.405 1.965 89.575 ;
        RECT 10.775 89.405 10.945 89.575 ;
        RECT 1.795 88.945 1.965 89.115 ;
        RECT 10.775 88.945 10.945 89.115 ;
        RECT 11.715 89.865 11.885 90.035 ;
        RECT 20.695 89.865 20.865 90.035 ;
        RECT 21.165 89.940 21.335 90.110 ;
        RECT 11.715 89.405 11.885 89.575 ;
        RECT 20.695 89.405 20.865 89.575 ;
        RECT 11.715 88.945 11.885 89.115 ;
        RECT 20.695 88.945 20.865 89.115 ;
        RECT 21.635 89.865 21.805 90.035 ;
        RECT 21.635 89.405 21.805 89.575 ;
        RECT 21.635 88.945 21.805 89.115 ;
        RECT -283.885 10.775 -283.715 10.945 ;
        RECT -283.415 10.770 -283.245 10.940 ;
        RECT -282.945 10.775 -282.775 10.945 ;
        RECT -283.885 10.315 -283.715 10.485 ;
        RECT -283.885 9.855 -283.715 10.025 ;
        RECT -273.965 10.775 -273.795 10.945 ;
        RECT -273.495 10.770 -273.325 10.940 ;
        RECT -273.025 10.775 -272.855 10.945 ;
        RECT -282.945 10.315 -282.775 10.485 ;
        RECT -273.965 10.315 -273.795 10.485 ;
        RECT -282.945 9.855 -282.775 10.025 ;
        RECT -273.965 9.855 -273.795 10.025 ;
        RECT -264.045 10.775 -263.875 10.945 ;
        RECT -263.575 10.770 -263.405 10.940 ;
        RECT -263.105 10.775 -262.935 10.945 ;
        RECT -273.025 10.315 -272.855 10.485 ;
        RECT -264.045 10.315 -263.875 10.485 ;
        RECT -273.025 9.855 -272.855 10.025 ;
        RECT -264.045 9.855 -263.875 10.025 ;
        RECT -254.125 10.775 -253.955 10.945 ;
        RECT -253.655 10.770 -253.485 10.940 ;
        RECT -253.185 10.775 -253.015 10.945 ;
        RECT -263.105 10.315 -262.935 10.485 ;
        RECT -254.125 10.315 -253.955 10.485 ;
        RECT -263.105 9.855 -262.935 10.025 ;
        RECT -254.125 9.855 -253.955 10.025 ;
        RECT -244.205 10.775 -244.035 10.945 ;
        RECT -243.735 10.770 -243.565 10.940 ;
        RECT -243.265 10.775 -243.095 10.945 ;
        RECT -253.185 10.315 -253.015 10.485 ;
        RECT -244.205 10.315 -244.035 10.485 ;
        RECT -253.185 9.855 -253.015 10.025 ;
        RECT -244.205 9.855 -244.035 10.025 ;
        RECT -234.285 10.775 -234.115 10.945 ;
        RECT -233.815 10.770 -233.645 10.940 ;
        RECT -233.345 10.775 -233.175 10.945 ;
        RECT -243.265 10.315 -243.095 10.485 ;
        RECT -234.285 10.315 -234.115 10.485 ;
        RECT -243.265 9.855 -243.095 10.025 ;
        RECT -234.285 9.855 -234.115 10.025 ;
        RECT -224.365 10.775 -224.195 10.945 ;
        RECT -223.895 10.770 -223.725 10.940 ;
        RECT -223.425 10.775 -223.255 10.945 ;
        RECT -233.345 10.315 -233.175 10.485 ;
        RECT -224.365 10.315 -224.195 10.485 ;
        RECT -233.345 9.855 -233.175 10.025 ;
        RECT -224.365 9.855 -224.195 10.025 ;
        RECT -214.445 10.775 -214.275 10.945 ;
        RECT -213.975 10.770 -213.805 10.940 ;
        RECT -213.505 10.775 -213.335 10.945 ;
        RECT -223.425 10.315 -223.255 10.485 ;
        RECT -214.445 10.315 -214.275 10.485 ;
        RECT -223.425 9.855 -223.255 10.025 ;
        RECT -214.445 9.855 -214.275 10.025 ;
        RECT -204.525 10.775 -204.355 10.945 ;
        RECT -204.055 10.770 -203.885 10.940 ;
        RECT -203.585 10.775 -203.415 10.945 ;
        RECT -213.505 10.315 -213.335 10.485 ;
        RECT -204.525 10.315 -204.355 10.485 ;
        RECT -213.505 9.855 -213.335 10.025 ;
        RECT -204.525 9.855 -204.355 10.025 ;
        RECT -194.605 10.775 -194.435 10.945 ;
        RECT -194.135 10.770 -193.965 10.940 ;
        RECT -193.665 10.775 -193.495 10.945 ;
        RECT -203.585 10.315 -203.415 10.485 ;
        RECT -194.605 10.315 -194.435 10.485 ;
        RECT -203.585 9.855 -203.415 10.025 ;
        RECT -194.605 9.855 -194.435 10.025 ;
        RECT -184.685 10.775 -184.515 10.945 ;
        RECT -184.215 10.770 -184.045 10.940 ;
        RECT -183.745 10.775 -183.575 10.945 ;
        RECT -193.665 10.315 -193.495 10.485 ;
        RECT -184.685 10.315 -184.515 10.485 ;
        RECT -193.665 9.855 -193.495 10.025 ;
        RECT -184.685 9.855 -184.515 10.025 ;
        RECT -174.765 10.775 -174.595 10.945 ;
        RECT -174.295 10.770 -174.125 10.940 ;
        RECT -173.825 10.775 -173.655 10.945 ;
        RECT -183.745 10.315 -183.575 10.485 ;
        RECT -174.765 10.315 -174.595 10.485 ;
        RECT -183.745 9.855 -183.575 10.025 ;
        RECT -174.765 9.855 -174.595 10.025 ;
        RECT -164.845 10.775 -164.675 10.945 ;
        RECT -164.375 10.770 -164.205 10.940 ;
        RECT -163.905 10.775 -163.735 10.945 ;
        RECT -173.825 10.315 -173.655 10.485 ;
        RECT -164.845 10.315 -164.675 10.485 ;
        RECT -173.825 9.855 -173.655 10.025 ;
        RECT -164.845 9.855 -164.675 10.025 ;
        RECT -154.925 10.775 -154.755 10.945 ;
        RECT -154.455 10.770 -154.285 10.940 ;
        RECT -153.985 10.775 -153.815 10.945 ;
        RECT -163.905 10.315 -163.735 10.485 ;
        RECT -154.925 10.315 -154.755 10.485 ;
        RECT -163.905 9.855 -163.735 10.025 ;
        RECT -154.925 9.855 -154.755 10.025 ;
        RECT -145.005 10.775 -144.835 10.945 ;
        RECT -144.535 10.770 -144.365 10.940 ;
        RECT -144.065 10.775 -143.895 10.945 ;
        RECT -153.985 10.315 -153.815 10.485 ;
        RECT -145.005 10.315 -144.835 10.485 ;
        RECT -153.985 9.855 -153.815 10.025 ;
        RECT -145.005 9.855 -144.835 10.025 ;
        RECT -135.085 10.775 -134.915 10.945 ;
        RECT -134.615 10.770 -134.445 10.940 ;
        RECT -134.145 10.775 -133.975 10.945 ;
        RECT -144.065 10.315 -143.895 10.485 ;
        RECT -135.085 10.315 -134.915 10.485 ;
        RECT -144.065 9.855 -143.895 10.025 ;
        RECT -135.085 9.855 -134.915 10.025 ;
        RECT -125.165 10.775 -124.995 10.945 ;
        RECT -124.695 10.770 -124.525 10.940 ;
        RECT -124.225 10.775 -124.055 10.945 ;
        RECT -134.145 10.315 -133.975 10.485 ;
        RECT -125.165 10.315 -124.995 10.485 ;
        RECT -134.145 9.855 -133.975 10.025 ;
        RECT -125.165 9.855 -124.995 10.025 ;
        RECT -115.245 10.775 -115.075 10.945 ;
        RECT -114.775 10.770 -114.605 10.940 ;
        RECT -114.305 10.775 -114.135 10.945 ;
        RECT -124.225 10.315 -124.055 10.485 ;
        RECT -115.245 10.315 -115.075 10.485 ;
        RECT -124.225 9.855 -124.055 10.025 ;
        RECT -115.245 9.855 -115.075 10.025 ;
        RECT -105.325 10.775 -105.155 10.945 ;
        RECT -104.855 10.770 -104.685 10.940 ;
        RECT -104.385 10.775 -104.215 10.945 ;
        RECT -114.305 10.315 -114.135 10.485 ;
        RECT -105.325 10.315 -105.155 10.485 ;
        RECT -114.305 9.855 -114.135 10.025 ;
        RECT -105.325 9.855 -105.155 10.025 ;
        RECT -95.405 10.775 -95.235 10.945 ;
        RECT -94.935 10.770 -94.765 10.940 ;
        RECT -94.465 10.775 -94.295 10.945 ;
        RECT -104.385 10.315 -104.215 10.485 ;
        RECT -95.405 10.315 -95.235 10.485 ;
        RECT -104.385 9.855 -104.215 10.025 ;
        RECT -95.405 9.855 -95.235 10.025 ;
        RECT -85.485 10.775 -85.315 10.945 ;
        RECT -85.015 10.770 -84.845 10.940 ;
        RECT -84.545 10.775 -84.375 10.945 ;
        RECT -94.465 10.315 -94.295 10.485 ;
        RECT -85.485 10.315 -85.315 10.485 ;
        RECT -94.465 9.855 -94.295 10.025 ;
        RECT -85.485 9.855 -85.315 10.025 ;
        RECT -75.565 10.775 -75.395 10.945 ;
        RECT -75.095 10.770 -74.925 10.940 ;
        RECT -74.625 10.775 -74.455 10.945 ;
        RECT -84.545 10.315 -84.375 10.485 ;
        RECT -75.565 10.315 -75.395 10.485 ;
        RECT -84.545 9.855 -84.375 10.025 ;
        RECT -75.565 9.855 -75.395 10.025 ;
        RECT -65.645 10.775 -65.475 10.945 ;
        RECT -65.175 10.770 -65.005 10.940 ;
        RECT -64.705 10.775 -64.535 10.945 ;
        RECT -74.625 10.315 -74.455 10.485 ;
        RECT -65.645 10.315 -65.475 10.485 ;
        RECT -74.625 9.855 -74.455 10.025 ;
        RECT -65.645 9.855 -65.475 10.025 ;
        RECT -55.725 10.775 -55.555 10.945 ;
        RECT -55.255 10.770 -55.085 10.940 ;
        RECT -54.785 10.775 -54.615 10.945 ;
        RECT -64.705 10.315 -64.535 10.485 ;
        RECT -55.725 10.315 -55.555 10.485 ;
        RECT -64.705 9.855 -64.535 10.025 ;
        RECT -55.725 9.855 -55.555 10.025 ;
        RECT -45.805 10.775 -45.635 10.945 ;
        RECT -45.335 10.770 -45.165 10.940 ;
        RECT -44.865 10.775 -44.695 10.945 ;
        RECT -54.785 10.315 -54.615 10.485 ;
        RECT -45.805 10.315 -45.635 10.485 ;
        RECT -54.785 9.855 -54.615 10.025 ;
        RECT -45.805 9.855 -45.635 10.025 ;
        RECT -35.885 10.775 -35.715 10.945 ;
        RECT -35.415 10.770 -35.245 10.940 ;
        RECT -34.945 10.775 -34.775 10.945 ;
        RECT -44.865 10.315 -44.695 10.485 ;
        RECT -35.885 10.315 -35.715 10.485 ;
        RECT -44.865 9.855 -44.695 10.025 ;
        RECT -35.885 9.855 -35.715 10.025 ;
        RECT -25.965 10.775 -25.795 10.945 ;
        RECT -25.495 10.770 -25.325 10.940 ;
        RECT -25.025 10.775 -24.855 10.945 ;
        RECT -34.945 10.315 -34.775 10.485 ;
        RECT -25.965 10.315 -25.795 10.485 ;
        RECT -34.945 9.855 -34.775 10.025 ;
        RECT -25.965 9.855 -25.795 10.025 ;
        RECT -16.045 10.775 -15.875 10.945 ;
        RECT -15.575 10.770 -15.405 10.940 ;
        RECT -15.105 10.775 -14.935 10.945 ;
        RECT -25.025 10.315 -24.855 10.485 ;
        RECT -16.045 10.315 -15.875 10.485 ;
        RECT -25.025 9.855 -24.855 10.025 ;
        RECT -16.045 9.855 -15.875 10.025 ;
        RECT -6.125 10.775 -5.955 10.945 ;
        RECT -5.655 10.770 -5.485 10.940 ;
        RECT -5.185 10.775 -5.015 10.945 ;
        RECT -15.105 10.315 -14.935 10.485 ;
        RECT -6.125 10.315 -5.955 10.485 ;
        RECT -15.105 9.855 -14.935 10.025 ;
        RECT -6.125 9.855 -5.955 10.025 ;
        RECT 3.795 10.775 3.965 10.945 ;
        RECT 4.265 10.770 4.435 10.940 ;
        RECT 4.735 10.775 4.905 10.945 ;
        RECT -5.185 10.315 -5.015 10.485 ;
        RECT 3.795 10.315 3.965 10.485 ;
        RECT -5.185 9.855 -5.015 10.025 ;
        RECT 3.795 9.855 3.965 10.025 ;
        RECT 13.715 10.775 13.885 10.945 ;
        RECT 14.185 10.770 14.355 10.940 ;
        RECT 14.655 10.775 14.825 10.945 ;
        RECT 4.735 10.315 4.905 10.485 ;
        RECT 13.715 10.315 13.885 10.485 ;
        RECT 4.735 9.855 4.905 10.025 ;
        RECT 13.715 9.855 13.885 10.025 ;
        RECT 23.635 10.775 23.805 10.945 ;
        RECT 24.105 10.770 24.275 10.940 ;
        RECT 14.655 10.315 14.825 10.485 ;
        RECT 23.635 10.315 23.805 10.485 ;
        RECT 14.655 9.855 14.825 10.025 ;
        RECT 23.635 9.855 23.805 10.025 ;
        RECT -289.755 9.195 -289.585 9.365 ;
        RECT -289.295 9.195 -289.125 9.365 ;
        RECT -288.835 9.195 -288.665 9.365 ;
        RECT -288.375 9.195 -288.205 9.365 ;
        RECT -287.915 9.195 -287.745 9.365 ;
        RECT -287.455 9.195 -287.285 9.365 ;
        RECT -286.995 9.195 -286.825 9.365 ;
        RECT -279.835 9.195 -279.665 9.365 ;
        RECT -279.375 9.195 -279.205 9.365 ;
        RECT -278.915 9.195 -278.745 9.365 ;
        RECT -278.455 9.195 -278.285 9.365 ;
        RECT -277.995 9.195 -277.825 9.365 ;
        RECT -277.535 9.195 -277.365 9.365 ;
        RECT -277.075 9.195 -276.905 9.365 ;
        RECT -269.915 9.195 -269.745 9.365 ;
        RECT -269.455 9.195 -269.285 9.365 ;
        RECT -268.995 9.195 -268.825 9.365 ;
        RECT -268.535 9.195 -268.365 9.365 ;
        RECT -268.075 9.195 -267.905 9.365 ;
        RECT -267.615 9.195 -267.445 9.365 ;
        RECT -267.155 9.195 -266.985 9.365 ;
        RECT -259.995 9.195 -259.825 9.365 ;
        RECT -259.535 9.195 -259.365 9.365 ;
        RECT -259.075 9.195 -258.905 9.365 ;
        RECT -258.615 9.195 -258.445 9.365 ;
        RECT -258.155 9.195 -257.985 9.365 ;
        RECT -257.695 9.195 -257.525 9.365 ;
        RECT -257.235 9.195 -257.065 9.365 ;
        RECT -250.075 9.195 -249.905 9.365 ;
        RECT -249.615 9.195 -249.445 9.365 ;
        RECT -249.155 9.195 -248.985 9.365 ;
        RECT -248.695 9.195 -248.525 9.365 ;
        RECT -248.235 9.195 -248.065 9.365 ;
        RECT -247.775 9.195 -247.605 9.365 ;
        RECT -247.315 9.195 -247.145 9.365 ;
        RECT -240.155 9.195 -239.985 9.365 ;
        RECT -239.695 9.195 -239.525 9.365 ;
        RECT -239.235 9.195 -239.065 9.365 ;
        RECT -238.775 9.195 -238.605 9.365 ;
        RECT -238.315 9.195 -238.145 9.365 ;
        RECT -237.855 9.195 -237.685 9.365 ;
        RECT -237.395 9.195 -237.225 9.365 ;
        RECT -230.235 9.195 -230.065 9.365 ;
        RECT -229.775 9.195 -229.605 9.365 ;
        RECT -229.315 9.195 -229.145 9.365 ;
        RECT -228.855 9.195 -228.685 9.365 ;
        RECT -228.395 9.195 -228.225 9.365 ;
        RECT -227.935 9.195 -227.765 9.365 ;
        RECT -227.475 9.195 -227.305 9.365 ;
        RECT -220.315 9.195 -220.145 9.365 ;
        RECT -219.855 9.195 -219.685 9.365 ;
        RECT -219.395 9.195 -219.225 9.365 ;
        RECT -218.935 9.195 -218.765 9.365 ;
        RECT -218.475 9.195 -218.305 9.365 ;
        RECT -218.015 9.195 -217.845 9.365 ;
        RECT -217.555 9.195 -217.385 9.365 ;
        RECT -210.395 9.195 -210.225 9.365 ;
        RECT -209.935 9.195 -209.765 9.365 ;
        RECT -209.475 9.195 -209.305 9.365 ;
        RECT -209.015 9.195 -208.845 9.365 ;
        RECT -208.555 9.195 -208.385 9.365 ;
        RECT -208.095 9.195 -207.925 9.365 ;
        RECT -207.635 9.195 -207.465 9.365 ;
        RECT -200.475 9.195 -200.305 9.365 ;
        RECT -200.015 9.195 -199.845 9.365 ;
        RECT -199.555 9.195 -199.385 9.365 ;
        RECT -199.095 9.195 -198.925 9.365 ;
        RECT -198.635 9.195 -198.465 9.365 ;
        RECT -198.175 9.195 -198.005 9.365 ;
        RECT -197.715 9.195 -197.545 9.365 ;
        RECT -190.555 9.195 -190.385 9.365 ;
        RECT -190.095 9.195 -189.925 9.365 ;
        RECT -189.635 9.195 -189.465 9.365 ;
        RECT -189.175 9.195 -189.005 9.365 ;
        RECT -188.715 9.195 -188.545 9.365 ;
        RECT -188.255 9.195 -188.085 9.365 ;
        RECT -187.795 9.195 -187.625 9.365 ;
        RECT -180.635 9.195 -180.465 9.365 ;
        RECT -180.175 9.195 -180.005 9.365 ;
        RECT -179.715 9.195 -179.545 9.365 ;
        RECT -179.255 9.195 -179.085 9.365 ;
        RECT -178.795 9.195 -178.625 9.365 ;
        RECT -178.335 9.195 -178.165 9.365 ;
        RECT -177.875 9.195 -177.705 9.365 ;
        RECT -170.715 9.195 -170.545 9.365 ;
        RECT -170.255 9.195 -170.085 9.365 ;
        RECT -169.795 9.195 -169.625 9.365 ;
        RECT -169.335 9.195 -169.165 9.365 ;
        RECT -168.875 9.195 -168.705 9.365 ;
        RECT -168.415 9.195 -168.245 9.365 ;
        RECT -167.955 9.195 -167.785 9.365 ;
        RECT -160.795 9.195 -160.625 9.365 ;
        RECT -160.335 9.195 -160.165 9.365 ;
        RECT -159.875 9.195 -159.705 9.365 ;
        RECT -159.415 9.195 -159.245 9.365 ;
        RECT -158.955 9.195 -158.785 9.365 ;
        RECT -158.495 9.195 -158.325 9.365 ;
        RECT -158.035 9.195 -157.865 9.365 ;
        RECT -150.875 9.195 -150.705 9.365 ;
        RECT -150.415 9.195 -150.245 9.365 ;
        RECT -149.955 9.195 -149.785 9.365 ;
        RECT -149.495 9.195 -149.325 9.365 ;
        RECT -149.035 9.195 -148.865 9.365 ;
        RECT -148.575 9.195 -148.405 9.365 ;
        RECT -148.115 9.195 -147.945 9.365 ;
        RECT -140.955 9.195 -140.785 9.365 ;
        RECT -140.495 9.195 -140.325 9.365 ;
        RECT -140.035 9.195 -139.865 9.365 ;
        RECT -139.575 9.195 -139.405 9.365 ;
        RECT -139.115 9.195 -138.945 9.365 ;
        RECT -138.655 9.195 -138.485 9.365 ;
        RECT -138.195 9.195 -138.025 9.365 ;
        RECT -131.035 9.195 -130.865 9.365 ;
        RECT -130.575 9.195 -130.405 9.365 ;
        RECT -130.115 9.195 -129.945 9.365 ;
        RECT -129.655 9.195 -129.485 9.365 ;
        RECT -129.195 9.195 -129.025 9.365 ;
        RECT -128.735 9.195 -128.565 9.365 ;
        RECT -128.275 9.195 -128.105 9.365 ;
        RECT -121.115 9.195 -120.945 9.365 ;
        RECT -120.655 9.195 -120.485 9.365 ;
        RECT -120.195 9.195 -120.025 9.365 ;
        RECT -119.735 9.195 -119.565 9.365 ;
        RECT -119.275 9.195 -119.105 9.365 ;
        RECT -118.815 9.195 -118.645 9.365 ;
        RECT -118.355 9.195 -118.185 9.365 ;
        RECT -111.195 9.195 -111.025 9.365 ;
        RECT -110.735 9.195 -110.565 9.365 ;
        RECT -110.275 9.195 -110.105 9.365 ;
        RECT -109.815 9.195 -109.645 9.365 ;
        RECT -109.355 9.195 -109.185 9.365 ;
        RECT -108.895 9.195 -108.725 9.365 ;
        RECT -108.435 9.195 -108.265 9.365 ;
        RECT -101.275 9.195 -101.105 9.365 ;
        RECT -100.815 9.195 -100.645 9.365 ;
        RECT -100.355 9.195 -100.185 9.365 ;
        RECT -99.895 9.195 -99.725 9.365 ;
        RECT -99.435 9.195 -99.265 9.365 ;
        RECT -98.975 9.195 -98.805 9.365 ;
        RECT -98.515 9.195 -98.345 9.365 ;
        RECT -91.355 9.195 -91.185 9.365 ;
        RECT -90.895 9.195 -90.725 9.365 ;
        RECT -90.435 9.195 -90.265 9.365 ;
        RECT -89.975 9.195 -89.805 9.365 ;
        RECT -89.515 9.195 -89.345 9.365 ;
        RECT -89.055 9.195 -88.885 9.365 ;
        RECT -88.595 9.195 -88.425 9.365 ;
        RECT -81.435 9.195 -81.265 9.365 ;
        RECT -80.975 9.195 -80.805 9.365 ;
        RECT -80.515 9.195 -80.345 9.365 ;
        RECT -80.055 9.195 -79.885 9.365 ;
        RECT -79.595 9.195 -79.425 9.365 ;
        RECT -79.135 9.195 -78.965 9.365 ;
        RECT -78.675 9.195 -78.505 9.365 ;
        RECT -71.515 9.195 -71.345 9.365 ;
        RECT -71.055 9.195 -70.885 9.365 ;
        RECT -70.595 9.195 -70.425 9.365 ;
        RECT -70.135 9.195 -69.965 9.365 ;
        RECT -69.675 9.195 -69.505 9.365 ;
        RECT -69.215 9.195 -69.045 9.365 ;
        RECT -68.755 9.195 -68.585 9.365 ;
        RECT -61.595 9.195 -61.425 9.365 ;
        RECT -61.135 9.195 -60.965 9.365 ;
        RECT -60.675 9.195 -60.505 9.365 ;
        RECT -60.215 9.195 -60.045 9.365 ;
        RECT -59.755 9.195 -59.585 9.365 ;
        RECT -59.295 9.195 -59.125 9.365 ;
        RECT -58.835 9.195 -58.665 9.365 ;
        RECT -51.675 9.195 -51.505 9.365 ;
        RECT -51.215 9.195 -51.045 9.365 ;
        RECT -50.755 9.195 -50.585 9.365 ;
        RECT -50.295 9.195 -50.125 9.365 ;
        RECT -49.835 9.195 -49.665 9.365 ;
        RECT -49.375 9.195 -49.205 9.365 ;
        RECT -48.915 9.195 -48.745 9.365 ;
        RECT -41.755 9.195 -41.585 9.365 ;
        RECT -41.295 9.195 -41.125 9.365 ;
        RECT -40.835 9.195 -40.665 9.365 ;
        RECT -40.375 9.195 -40.205 9.365 ;
        RECT -39.915 9.195 -39.745 9.365 ;
        RECT -39.455 9.195 -39.285 9.365 ;
        RECT -38.995 9.195 -38.825 9.365 ;
        RECT -31.835 9.195 -31.665 9.365 ;
        RECT -31.375 9.195 -31.205 9.365 ;
        RECT -30.915 9.195 -30.745 9.365 ;
        RECT -30.455 9.195 -30.285 9.365 ;
        RECT -29.995 9.195 -29.825 9.365 ;
        RECT -29.535 9.195 -29.365 9.365 ;
        RECT -29.075 9.195 -28.905 9.365 ;
        RECT -21.915 9.195 -21.745 9.365 ;
        RECT -21.455 9.195 -21.285 9.365 ;
        RECT -20.995 9.195 -20.825 9.365 ;
        RECT -20.535 9.195 -20.365 9.365 ;
        RECT -20.075 9.195 -19.905 9.365 ;
        RECT -19.615 9.195 -19.445 9.365 ;
        RECT -19.155 9.195 -18.985 9.365 ;
        RECT -11.995 9.195 -11.825 9.365 ;
        RECT -11.535 9.195 -11.365 9.365 ;
        RECT -11.075 9.195 -10.905 9.365 ;
        RECT -10.615 9.195 -10.445 9.365 ;
        RECT -10.155 9.195 -9.985 9.365 ;
        RECT -9.695 9.195 -9.525 9.365 ;
        RECT -9.235 9.195 -9.065 9.365 ;
        RECT -2.075 9.195 -1.905 9.365 ;
        RECT -1.615 9.195 -1.445 9.365 ;
        RECT -1.155 9.195 -0.985 9.365 ;
        RECT -0.695 9.195 -0.525 9.365 ;
        RECT -0.235 9.195 -0.065 9.365 ;
        RECT 0.225 9.195 0.395 9.365 ;
        RECT 0.685 9.195 0.855 9.365 ;
        RECT 7.845 9.195 8.015 9.365 ;
        RECT 8.305 9.195 8.475 9.365 ;
        RECT 8.765 9.195 8.935 9.365 ;
        RECT 9.225 9.195 9.395 9.365 ;
        RECT 9.685 9.195 9.855 9.365 ;
        RECT 10.145 9.195 10.315 9.365 ;
        RECT 10.605 9.195 10.775 9.365 ;
        RECT 17.765 9.195 17.935 9.365 ;
        RECT 18.225 9.195 18.395 9.365 ;
        RECT 18.685 9.195 18.855 9.365 ;
        RECT 19.145 9.195 19.315 9.365 ;
        RECT 19.605 9.195 19.775 9.365 ;
        RECT 20.065 9.195 20.235 9.365 ;
        RECT 20.525 9.195 20.695 9.365 ;
        RECT -284.795 6.475 -284.625 6.645 ;
        RECT -284.335 6.475 -284.165 6.645 ;
        RECT -283.875 6.475 -283.705 6.645 ;
        RECT -283.415 6.475 -283.245 6.645 ;
        RECT -282.955 6.475 -282.785 6.645 ;
        RECT -282.495 6.475 -282.325 6.645 ;
        RECT -282.035 6.475 -281.865 6.645 ;
        RECT -274.875 6.475 -274.705 6.645 ;
        RECT -274.415 6.475 -274.245 6.645 ;
        RECT -273.955 6.475 -273.785 6.645 ;
        RECT -273.495 6.475 -273.325 6.645 ;
        RECT -273.035 6.475 -272.865 6.645 ;
        RECT -272.575 6.475 -272.405 6.645 ;
        RECT -272.115 6.475 -271.945 6.645 ;
        RECT -264.955 6.475 -264.785 6.645 ;
        RECT -264.495 6.475 -264.325 6.645 ;
        RECT -264.035 6.475 -263.865 6.645 ;
        RECT -263.575 6.475 -263.405 6.645 ;
        RECT -263.115 6.475 -262.945 6.645 ;
        RECT -262.655 6.475 -262.485 6.645 ;
        RECT -262.195 6.475 -262.025 6.645 ;
        RECT -255.035 6.475 -254.865 6.645 ;
        RECT -254.575 6.475 -254.405 6.645 ;
        RECT -254.115 6.475 -253.945 6.645 ;
        RECT -253.655 6.475 -253.485 6.645 ;
        RECT -253.195 6.475 -253.025 6.645 ;
        RECT -252.735 6.475 -252.565 6.645 ;
        RECT -252.275 6.475 -252.105 6.645 ;
        RECT -245.115 6.475 -244.945 6.645 ;
        RECT -244.655 6.475 -244.485 6.645 ;
        RECT -244.195 6.475 -244.025 6.645 ;
        RECT -243.735 6.475 -243.565 6.645 ;
        RECT -243.275 6.475 -243.105 6.645 ;
        RECT -242.815 6.475 -242.645 6.645 ;
        RECT -242.355 6.475 -242.185 6.645 ;
        RECT -235.195 6.475 -235.025 6.645 ;
        RECT -234.735 6.475 -234.565 6.645 ;
        RECT -234.275 6.475 -234.105 6.645 ;
        RECT -233.815 6.475 -233.645 6.645 ;
        RECT -233.355 6.475 -233.185 6.645 ;
        RECT -232.895 6.475 -232.725 6.645 ;
        RECT -232.435 6.475 -232.265 6.645 ;
        RECT -225.275 6.475 -225.105 6.645 ;
        RECT -224.815 6.475 -224.645 6.645 ;
        RECT -224.355 6.475 -224.185 6.645 ;
        RECT -223.895 6.475 -223.725 6.645 ;
        RECT -223.435 6.475 -223.265 6.645 ;
        RECT -222.975 6.475 -222.805 6.645 ;
        RECT -222.515 6.475 -222.345 6.645 ;
        RECT -215.355 6.475 -215.185 6.645 ;
        RECT -214.895 6.475 -214.725 6.645 ;
        RECT -214.435 6.475 -214.265 6.645 ;
        RECT -213.975 6.475 -213.805 6.645 ;
        RECT -213.515 6.475 -213.345 6.645 ;
        RECT -213.055 6.475 -212.885 6.645 ;
        RECT -212.595 6.475 -212.425 6.645 ;
        RECT -205.435 6.475 -205.265 6.645 ;
        RECT -204.975 6.475 -204.805 6.645 ;
        RECT -204.515 6.475 -204.345 6.645 ;
        RECT -204.055 6.475 -203.885 6.645 ;
        RECT -203.595 6.475 -203.425 6.645 ;
        RECT -203.135 6.475 -202.965 6.645 ;
        RECT -202.675 6.475 -202.505 6.645 ;
        RECT -195.515 6.475 -195.345 6.645 ;
        RECT -195.055 6.475 -194.885 6.645 ;
        RECT -194.595 6.475 -194.425 6.645 ;
        RECT -194.135 6.475 -193.965 6.645 ;
        RECT -193.675 6.475 -193.505 6.645 ;
        RECT -193.215 6.475 -193.045 6.645 ;
        RECT -192.755 6.475 -192.585 6.645 ;
        RECT -185.595 6.475 -185.425 6.645 ;
        RECT -185.135 6.475 -184.965 6.645 ;
        RECT -184.675 6.475 -184.505 6.645 ;
        RECT -184.215 6.475 -184.045 6.645 ;
        RECT -183.755 6.475 -183.585 6.645 ;
        RECT -183.295 6.475 -183.125 6.645 ;
        RECT -182.835 6.475 -182.665 6.645 ;
        RECT -175.675 6.475 -175.505 6.645 ;
        RECT -175.215 6.475 -175.045 6.645 ;
        RECT -174.755 6.475 -174.585 6.645 ;
        RECT -174.295 6.475 -174.125 6.645 ;
        RECT -173.835 6.475 -173.665 6.645 ;
        RECT -173.375 6.475 -173.205 6.645 ;
        RECT -172.915 6.475 -172.745 6.645 ;
        RECT -165.755 6.475 -165.585 6.645 ;
        RECT -165.295 6.475 -165.125 6.645 ;
        RECT -164.835 6.475 -164.665 6.645 ;
        RECT -164.375 6.475 -164.205 6.645 ;
        RECT -163.915 6.475 -163.745 6.645 ;
        RECT -163.455 6.475 -163.285 6.645 ;
        RECT -162.995 6.475 -162.825 6.645 ;
        RECT -155.835 6.475 -155.665 6.645 ;
        RECT -155.375 6.475 -155.205 6.645 ;
        RECT -154.915 6.475 -154.745 6.645 ;
        RECT -154.455 6.475 -154.285 6.645 ;
        RECT -153.995 6.475 -153.825 6.645 ;
        RECT -153.535 6.475 -153.365 6.645 ;
        RECT -153.075 6.475 -152.905 6.645 ;
        RECT -145.915 6.475 -145.745 6.645 ;
        RECT -145.455 6.475 -145.285 6.645 ;
        RECT -144.995 6.475 -144.825 6.645 ;
        RECT -144.535 6.475 -144.365 6.645 ;
        RECT -144.075 6.475 -143.905 6.645 ;
        RECT -143.615 6.475 -143.445 6.645 ;
        RECT -143.155 6.475 -142.985 6.645 ;
        RECT -135.995 6.475 -135.825 6.645 ;
        RECT -135.535 6.475 -135.365 6.645 ;
        RECT -135.075 6.475 -134.905 6.645 ;
        RECT -134.615 6.475 -134.445 6.645 ;
        RECT -134.155 6.475 -133.985 6.645 ;
        RECT -133.695 6.475 -133.525 6.645 ;
        RECT -133.235 6.475 -133.065 6.645 ;
        RECT -126.075 6.475 -125.905 6.645 ;
        RECT -125.615 6.475 -125.445 6.645 ;
        RECT -125.155 6.475 -124.985 6.645 ;
        RECT -124.695 6.475 -124.525 6.645 ;
        RECT -124.235 6.475 -124.065 6.645 ;
        RECT -123.775 6.475 -123.605 6.645 ;
        RECT -123.315 6.475 -123.145 6.645 ;
        RECT -116.155 6.475 -115.985 6.645 ;
        RECT -115.695 6.475 -115.525 6.645 ;
        RECT -115.235 6.475 -115.065 6.645 ;
        RECT -114.775 6.475 -114.605 6.645 ;
        RECT -114.315 6.475 -114.145 6.645 ;
        RECT -113.855 6.475 -113.685 6.645 ;
        RECT -113.395 6.475 -113.225 6.645 ;
        RECT -106.235 6.475 -106.065 6.645 ;
        RECT -105.775 6.475 -105.605 6.645 ;
        RECT -105.315 6.475 -105.145 6.645 ;
        RECT -104.855 6.475 -104.685 6.645 ;
        RECT -104.395 6.475 -104.225 6.645 ;
        RECT -103.935 6.475 -103.765 6.645 ;
        RECT -103.475 6.475 -103.305 6.645 ;
        RECT -96.315 6.475 -96.145 6.645 ;
        RECT -95.855 6.475 -95.685 6.645 ;
        RECT -95.395 6.475 -95.225 6.645 ;
        RECT -94.935 6.475 -94.765 6.645 ;
        RECT -94.475 6.475 -94.305 6.645 ;
        RECT -94.015 6.475 -93.845 6.645 ;
        RECT -93.555 6.475 -93.385 6.645 ;
        RECT -86.395 6.475 -86.225 6.645 ;
        RECT -85.935 6.475 -85.765 6.645 ;
        RECT -85.475 6.475 -85.305 6.645 ;
        RECT -85.015 6.475 -84.845 6.645 ;
        RECT -84.555 6.475 -84.385 6.645 ;
        RECT -84.095 6.475 -83.925 6.645 ;
        RECT -83.635 6.475 -83.465 6.645 ;
        RECT -76.475 6.475 -76.305 6.645 ;
        RECT -76.015 6.475 -75.845 6.645 ;
        RECT -75.555 6.475 -75.385 6.645 ;
        RECT -75.095 6.475 -74.925 6.645 ;
        RECT -74.635 6.475 -74.465 6.645 ;
        RECT -74.175 6.475 -74.005 6.645 ;
        RECT -73.715 6.475 -73.545 6.645 ;
        RECT -66.555 6.475 -66.385 6.645 ;
        RECT -66.095 6.475 -65.925 6.645 ;
        RECT -65.635 6.475 -65.465 6.645 ;
        RECT -65.175 6.475 -65.005 6.645 ;
        RECT -64.715 6.475 -64.545 6.645 ;
        RECT -64.255 6.475 -64.085 6.645 ;
        RECT -63.795 6.475 -63.625 6.645 ;
        RECT -56.635 6.475 -56.465 6.645 ;
        RECT -56.175 6.475 -56.005 6.645 ;
        RECT -55.715 6.475 -55.545 6.645 ;
        RECT -55.255 6.475 -55.085 6.645 ;
        RECT -54.795 6.475 -54.625 6.645 ;
        RECT -54.335 6.475 -54.165 6.645 ;
        RECT -53.875 6.475 -53.705 6.645 ;
        RECT -46.715 6.475 -46.545 6.645 ;
        RECT -46.255 6.475 -46.085 6.645 ;
        RECT -45.795 6.475 -45.625 6.645 ;
        RECT -45.335 6.475 -45.165 6.645 ;
        RECT -44.875 6.475 -44.705 6.645 ;
        RECT -44.415 6.475 -44.245 6.645 ;
        RECT -43.955 6.475 -43.785 6.645 ;
        RECT -36.795 6.475 -36.625 6.645 ;
        RECT -36.335 6.475 -36.165 6.645 ;
        RECT -35.875 6.475 -35.705 6.645 ;
        RECT -35.415 6.475 -35.245 6.645 ;
        RECT -34.955 6.475 -34.785 6.645 ;
        RECT -34.495 6.475 -34.325 6.645 ;
        RECT -34.035 6.475 -33.865 6.645 ;
        RECT -26.875 6.475 -26.705 6.645 ;
        RECT -26.415 6.475 -26.245 6.645 ;
        RECT -25.955 6.475 -25.785 6.645 ;
        RECT -25.495 6.475 -25.325 6.645 ;
        RECT -25.035 6.475 -24.865 6.645 ;
        RECT -24.575 6.475 -24.405 6.645 ;
        RECT -24.115 6.475 -23.945 6.645 ;
        RECT -16.955 6.475 -16.785 6.645 ;
        RECT -16.495 6.475 -16.325 6.645 ;
        RECT -16.035 6.475 -15.865 6.645 ;
        RECT -15.575 6.475 -15.405 6.645 ;
        RECT -15.115 6.475 -14.945 6.645 ;
        RECT -14.655 6.475 -14.485 6.645 ;
        RECT -14.195 6.475 -14.025 6.645 ;
        RECT -7.035 6.475 -6.865 6.645 ;
        RECT -6.575 6.475 -6.405 6.645 ;
        RECT -6.115 6.475 -5.945 6.645 ;
        RECT -5.655 6.475 -5.485 6.645 ;
        RECT -5.195 6.475 -5.025 6.645 ;
        RECT -4.735 6.475 -4.565 6.645 ;
        RECT -4.275 6.475 -4.105 6.645 ;
        RECT 2.885 6.475 3.055 6.645 ;
        RECT 3.345 6.475 3.515 6.645 ;
        RECT 3.805 6.475 3.975 6.645 ;
        RECT 4.265 6.475 4.435 6.645 ;
        RECT 4.725 6.475 4.895 6.645 ;
        RECT 5.185 6.475 5.355 6.645 ;
        RECT 5.645 6.475 5.815 6.645 ;
        RECT 12.805 6.475 12.975 6.645 ;
        RECT 13.265 6.475 13.435 6.645 ;
        RECT 13.725 6.475 13.895 6.645 ;
        RECT 14.185 6.475 14.355 6.645 ;
        RECT 14.645 6.475 14.815 6.645 ;
        RECT 15.105 6.475 15.275 6.645 ;
        RECT 15.565 6.475 15.735 6.645 ;
        RECT 22.725 6.475 22.895 6.645 ;
        RECT 23.185 6.475 23.355 6.645 ;
        RECT 23.645 6.475 23.815 6.645 ;
        RECT 24.105 6.475 24.275 6.645 ;
        RECT -288.845 5.815 -288.675 5.985 ;
        RECT -288.375 5.890 -288.205 6.060 ;
        RECT -288.845 5.355 -288.675 5.525 ;
        RECT -288.845 4.895 -288.675 5.065 ;
        RECT -287.905 5.815 -287.735 5.985 ;
        RECT -278.925 5.815 -278.755 5.985 ;
        RECT -278.455 5.890 -278.285 6.060 ;
        RECT -287.905 5.355 -287.735 5.525 ;
        RECT -278.925 5.355 -278.755 5.525 ;
        RECT -287.905 4.895 -287.735 5.065 ;
        RECT -278.925 4.895 -278.755 5.065 ;
        RECT -277.985 5.815 -277.815 5.985 ;
        RECT -269.005 5.815 -268.835 5.985 ;
        RECT -268.535 5.890 -268.365 6.060 ;
        RECT -277.985 5.355 -277.815 5.525 ;
        RECT -269.005 5.355 -268.835 5.525 ;
        RECT -277.985 4.895 -277.815 5.065 ;
        RECT -269.005 4.895 -268.835 5.065 ;
        RECT -268.065 5.815 -267.895 5.985 ;
        RECT -259.085 5.815 -258.915 5.985 ;
        RECT -258.615 5.890 -258.445 6.060 ;
        RECT -268.065 5.355 -267.895 5.525 ;
        RECT -259.085 5.355 -258.915 5.525 ;
        RECT -268.065 4.895 -267.895 5.065 ;
        RECT -259.085 4.895 -258.915 5.065 ;
        RECT -258.145 5.815 -257.975 5.985 ;
        RECT -249.165 5.815 -248.995 5.985 ;
        RECT -248.695 5.890 -248.525 6.060 ;
        RECT -258.145 5.355 -257.975 5.525 ;
        RECT -249.165 5.355 -248.995 5.525 ;
        RECT -258.145 4.895 -257.975 5.065 ;
        RECT -249.165 4.895 -248.995 5.065 ;
        RECT -248.225 5.815 -248.055 5.985 ;
        RECT -239.245 5.815 -239.075 5.985 ;
        RECT -238.775 5.890 -238.605 6.060 ;
        RECT -248.225 5.355 -248.055 5.525 ;
        RECT -239.245 5.355 -239.075 5.525 ;
        RECT -248.225 4.895 -248.055 5.065 ;
        RECT -239.245 4.895 -239.075 5.065 ;
        RECT -238.305 5.815 -238.135 5.985 ;
        RECT -229.325 5.815 -229.155 5.985 ;
        RECT -228.855 5.890 -228.685 6.060 ;
        RECT -238.305 5.355 -238.135 5.525 ;
        RECT -229.325 5.355 -229.155 5.525 ;
        RECT -238.305 4.895 -238.135 5.065 ;
        RECT -229.325 4.895 -229.155 5.065 ;
        RECT -228.385 5.815 -228.215 5.985 ;
        RECT -219.405 5.815 -219.235 5.985 ;
        RECT -218.935 5.890 -218.765 6.060 ;
        RECT -228.385 5.355 -228.215 5.525 ;
        RECT -219.405 5.355 -219.235 5.525 ;
        RECT -228.385 4.895 -228.215 5.065 ;
        RECT -219.405 4.895 -219.235 5.065 ;
        RECT -218.465 5.815 -218.295 5.985 ;
        RECT -209.485 5.815 -209.315 5.985 ;
        RECT -209.015 5.890 -208.845 6.060 ;
        RECT -218.465 5.355 -218.295 5.525 ;
        RECT -209.485 5.355 -209.315 5.525 ;
        RECT -218.465 4.895 -218.295 5.065 ;
        RECT -209.485 4.895 -209.315 5.065 ;
        RECT -208.545 5.815 -208.375 5.985 ;
        RECT -199.565 5.815 -199.395 5.985 ;
        RECT -199.095 5.890 -198.925 6.060 ;
        RECT -208.545 5.355 -208.375 5.525 ;
        RECT -199.565 5.355 -199.395 5.525 ;
        RECT -208.545 4.895 -208.375 5.065 ;
        RECT -199.565 4.895 -199.395 5.065 ;
        RECT -198.625 5.815 -198.455 5.985 ;
        RECT -189.645 5.815 -189.475 5.985 ;
        RECT -189.175 5.890 -189.005 6.060 ;
        RECT -198.625 5.355 -198.455 5.525 ;
        RECT -189.645 5.355 -189.475 5.525 ;
        RECT -198.625 4.895 -198.455 5.065 ;
        RECT -189.645 4.895 -189.475 5.065 ;
        RECT -188.705 5.815 -188.535 5.985 ;
        RECT -179.725 5.815 -179.555 5.985 ;
        RECT -179.255 5.890 -179.085 6.060 ;
        RECT -188.705 5.355 -188.535 5.525 ;
        RECT -179.725 5.355 -179.555 5.525 ;
        RECT -188.705 4.895 -188.535 5.065 ;
        RECT -179.725 4.895 -179.555 5.065 ;
        RECT -178.785 5.815 -178.615 5.985 ;
        RECT -169.805 5.815 -169.635 5.985 ;
        RECT -169.335 5.890 -169.165 6.060 ;
        RECT -178.785 5.355 -178.615 5.525 ;
        RECT -169.805 5.355 -169.635 5.525 ;
        RECT -178.785 4.895 -178.615 5.065 ;
        RECT -169.805 4.895 -169.635 5.065 ;
        RECT -168.865 5.815 -168.695 5.985 ;
        RECT -159.885 5.815 -159.715 5.985 ;
        RECT -159.415 5.890 -159.245 6.060 ;
        RECT -168.865 5.355 -168.695 5.525 ;
        RECT -159.885 5.355 -159.715 5.525 ;
        RECT -168.865 4.895 -168.695 5.065 ;
        RECT -159.885 4.895 -159.715 5.065 ;
        RECT -158.945 5.815 -158.775 5.985 ;
        RECT -149.965 5.815 -149.795 5.985 ;
        RECT -149.495 5.890 -149.325 6.060 ;
        RECT -158.945 5.355 -158.775 5.525 ;
        RECT -149.965 5.355 -149.795 5.525 ;
        RECT -158.945 4.895 -158.775 5.065 ;
        RECT -149.965 4.895 -149.795 5.065 ;
        RECT -149.025 5.815 -148.855 5.985 ;
        RECT -140.045 5.815 -139.875 5.985 ;
        RECT -139.575 5.890 -139.405 6.060 ;
        RECT -149.025 5.355 -148.855 5.525 ;
        RECT -140.045 5.355 -139.875 5.525 ;
        RECT -149.025 4.895 -148.855 5.065 ;
        RECT -140.045 4.895 -139.875 5.065 ;
        RECT -139.105 5.815 -138.935 5.985 ;
        RECT -130.125 5.815 -129.955 5.985 ;
        RECT -129.655 5.890 -129.485 6.060 ;
        RECT -139.105 5.355 -138.935 5.525 ;
        RECT -130.125 5.355 -129.955 5.525 ;
        RECT -139.105 4.895 -138.935 5.065 ;
        RECT -130.125 4.895 -129.955 5.065 ;
        RECT -129.185 5.815 -129.015 5.985 ;
        RECT -120.205 5.815 -120.035 5.985 ;
        RECT -119.735 5.890 -119.565 6.060 ;
        RECT -129.185 5.355 -129.015 5.525 ;
        RECT -120.205 5.355 -120.035 5.525 ;
        RECT -129.185 4.895 -129.015 5.065 ;
        RECT -120.205 4.895 -120.035 5.065 ;
        RECT -119.265 5.815 -119.095 5.985 ;
        RECT -110.285 5.815 -110.115 5.985 ;
        RECT -109.815 5.890 -109.645 6.060 ;
        RECT -119.265 5.355 -119.095 5.525 ;
        RECT -110.285 5.355 -110.115 5.525 ;
        RECT -119.265 4.895 -119.095 5.065 ;
        RECT -110.285 4.895 -110.115 5.065 ;
        RECT -109.345 5.815 -109.175 5.985 ;
        RECT -100.365 5.815 -100.195 5.985 ;
        RECT -99.895 5.890 -99.725 6.060 ;
        RECT -109.345 5.355 -109.175 5.525 ;
        RECT -100.365 5.355 -100.195 5.525 ;
        RECT -109.345 4.895 -109.175 5.065 ;
        RECT -100.365 4.895 -100.195 5.065 ;
        RECT -99.425 5.815 -99.255 5.985 ;
        RECT -90.445 5.815 -90.275 5.985 ;
        RECT -89.975 5.890 -89.805 6.060 ;
        RECT -99.425 5.355 -99.255 5.525 ;
        RECT -90.445 5.355 -90.275 5.525 ;
        RECT -99.425 4.895 -99.255 5.065 ;
        RECT -90.445 4.895 -90.275 5.065 ;
        RECT -89.505 5.815 -89.335 5.985 ;
        RECT -80.525 5.815 -80.355 5.985 ;
        RECT -80.055 5.890 -79.885 6.060 ;
        RECT -89.505 5.355 -89.335 5.525 ;
        RECT -80.525 5.355 -80.355 5.525 ;
        RECT -89.505 4.895 -89.335 5.065 ;
        RECT -80.525 4.895 -80.355 5.065 ;
        RECT -79.585 5.815 -79.415 5.985 ;
        RECT -70.605 5.815 -70.435 5.985 ;
        RECT -70.135 5.890 -69.965 6.060 ;
        RECT -79.585 5.355 -79.415 5.525 ;
        RECT -70.605 5.355 -70.435 5.525 ;
        RECT -79.585 4.895 -79.415 5.065 ;
        RECT -70.605 4.895 -70.435 5.065 ;
        RECT -69.665 5.815 -69.495 5.985 ;
        RECT -60.685 5.815 -60.515 5.985 ;
        RECT -60.215 5.890 -60.045 6.060 ;
        RECT -69.665 5.355 -69.495 5.525 ;
        RECT -60.685 5.355 -60.515 5.525 ;
        RECT -69.665 4.895 -69.495 5.065 ;
        RECT -60.685 4.895 -60.515 5.065 ;
        RECT -59.745 5.815 -59.575 5.985 ;
        RECT -50.765 5.815 -50.595 5.985 ;
        RECT -50.295 5.890 -50.125 6.060 ;
        RECT -59.745 5.355 -59.575 5.525 ;
        RECT -50.765 5.355 -50.595 5.525 ;
        RECT -59.745 4.895 -59.575 5.065 ;
        RECT -50.765 4.895 -50.595 5.065 ;
        RECT -49.825 5.815 -49.655 5.985 ;
        RECT -40.845 5.815 -40.675 5.985 ;
        RECT -40.375 5.890 -40.205 6.060 ;
        RECT -49.825 5.355 -49.655 5.525 ;
        RECT -40.845 5.355 -40.675 5.525 ;
        RECT -49.825 4.895 -49.655 5.065 ;
        RECT -40.845 4.895 -40.675 5.065 ;
        RECT -39.905 5.815 -39.735 5.985 ;
        RECT -30.925 5.815 -30.755 5.985 ;
        RECT -30.455 5.890 -30.285 6.060 ;
        RECT -39.905 5.355 -39.735 5.525 ;
        RECT -30.925 5.355 -30.755 5.525 ;
        RECT -39.905 4.895 -39.735 5.065 ;
        RECT -30.925 4.895 -30.755 5.065 ;
        RECT -29.985 5.815 -29.815 5.985 ;
        RECT -21.005 5.815 -20.835 5.985 ;
        RECT -20.535 5.890 -20.365 6.060 ;
        RECT -29.985 5.355 -29.815 5.525 ;
        RECT -21.005 5.355 -20.835 5.525 ;
        RECT -29.985 4.895 -29.815 5.065 ;
        RECT -21.005 4.895 -20.835 5.065 ;
        RECT -20.065 5.815 -19.895 5.985 ;
        RECT -11.085 5.815 -10.915 5.985 ;
        RECT -10.615 5.890 -10.445 6.060 ;
        RECT -20.065 5.355 -19.895 5.525 ;
        RECT -11.085 5.355 -10.915 5.525 ;
        RECT -20.065 4.895 -19.895 5.065 ;
        RECT -11.085 4.895 -10.915 5.065 ;
        RECT -10.145 5.815 -9.975 5.985 ;
        RECT -1.165 5.815 -0.995 5.985 ;
        RECT -0.695 5.890 -0.525 6.060 ;
        RECT -10.145 5.355 -9.975 5.525 ;
        RECT -1.165 5.355 -0.995 5.525 ;
        RECT -10.145 4.895 -9.975 5.065 ;
        RECT -1.165 4.895 -0.995 5.065 ;
        RECT -0.225 5.815 -0.055 5.985 ;
        RECT 8.755 5.815 8.925 5.985 ;
        RECT 9.225 5.890 9.395 6.060 ;
        RECT -0.225 5.355 -0.055 5.525 ;
        RECT 8.755 5.355 8.925 5.525 ;
        RECT -0.225 4.895 -0.055 5.065 ;
        RECT 8.755 4.895 8.925 5.065 ;
        RECT 9.695 5.815 9.865 5.985 ;
        RECT 18.675 5.815 18.845 5.985 ;
        RECT 19.145 5.890 19.315 6.060 ;
        RECT 9.695 5.355 9.865 5.525 ;
        RECT 18.675 5.355 18.845 5.525 ;
        RECT 9.695 4.895 9.865 5.065 ;
        RECT 18.675 4.895 18.845 5.065 ;
        RECT 19.615 5.815 19.785 5.985 ;
        RECT 19.615 5.355 19.785 5.525 ;
        RECT 19.615 4.895 19.785 5.065 ;
        RECT -283.525 -78.175 -283.355 -78.005 ;
        RECT -283.055 -78.180 -282.885 -78.010 ;
        RECT -282.585 -78.175 -282.415 -78.005 ;
        RECT -283.525 -78.635 -283.355 -78.465 ;
        RECT -283.525 -79.095 -283.355 -78.925 ;
        RECT -273.605 -78.175 -273.435 -78.005 ;
        RECT -273.135 -78.180 -272.965 -78.010 ;
        RECT -272.665 -78.175 -272.495 -78.005 ;
        RECT -282.585 -78.635 -282.415 -78.465 ;
        RECT -273.605 -78.635 -273.435 -78.465 ;
        RECT -282.585 -79.095 -282.415 -78.925 ;
        RECT -273.605 -79.095 -273.435 -78.925 ;
        RECT -263.685 -78.175 -263.515 -78.005 ;
        RECT -263.215 -78.180 -263.045 -78.010 ;
        RECT -262.745 -78.175 -262.575 -78.005 ;
        RECT -272.665 -78.635 -272.495 -78.465 ;
        RECT -263.685 -78.635 -263.515 -78.465 ;
        RECT -272.665 -79.095 -272.495 -78.925 ;
        RECT -263.685 -79.095 -263.515 -78.925 ;
        RECT -253.765 -78.175 -253.595 -78.005 ;
        RECT -253.295 -78.180 -253.125 -78.010 ;
        RECT -252.825 -78.175 -252.655 -78.005 ;
        RECT -262.745 -78.635 -262.575 -78.465 ;
        RECT -253.765 -78.635 -253.595 -78.465 ;
        RECT -262.745 -79.095 -262.575 -78.925 ;
        RECT -253.765 -79.095 -253.595 -78.925 ;
        RECT -243.845 -78.175 -243.675 -78.005 ;
        RECT -243.375 -78.180 -243.205 -78.010 ;
        RECT -242.905 -78.175 -242.735 -78.005 ;
        RECT -252.825 -78.635 -252.655 -78.465 ;
        RECT -243.845 -78.635 -243.675 -78.465 ;
        RECT -252.825 -79.095 -252.655 -78.925 ;
        RECT -243.845 -79.095 -243.675 -78.925 ;
        RECT -233.925 -78.175 -233.755 -78.005 ;
        RECT -233.455 -78.180 -233.285 -78.010 ;
        RECT -232.985 -78.175 -232.815 -78.005 ;
        RECT -242.905 -78.635 -242.735 -78.465 ;
        RECT -233.925 -78.635 -233.755 -78.465 ;
        RECT -242.905 -79.095 -242.735 -78.925 ;
        RECT -233.925 -79.095 -233.755 -78.925 ;
        RECT -224.005 -78.175 -223.835 -78.005 ;
        RECT -223.535 -78.180 -223.365 -78.010 ;
        RECT -223.065 -78.175 -222.895 -78.005 ;
        RECT -232.985 -78.635 -232.815 -78.465 ;
        RECT -224.005 -78.635 -223.835 -78.465 ;
        RECT -232.985 -79.095 -232.815 -78.925 ;
        RECT -224.005 -79.095 -223.835 -78.925 ;
        RECT -214.085 -78.175 -213.915 -78.005 ;
        RECT -213.615 -78.180 -213.445 -78.010 ;
        RECT -213.145 -78.175 -212.975 -78.005 ;
        RECT -223.065 -78.635 -222.895 -78.465 ;
        RECT -214.085 -78.635 -213.915 -78.465 ;
        RECT -223.065 -79.095 -222.895 -78.925 ;
        RECT -214.085 -79.095 -213.915 -78.925 ;
        RECT -204.165 -78.175 -203.995 -78.005 ;
        RECT -203.695 -78.180 -203.525 -78.010 ;
        RECT -203.225 -78.175 -203.055 -78.005 ;
        RECT -213.145 -78.635 -212.975 -78.465 ;
        RECT -204.165 -78.635 -203.995 -78.465 ;
        RECT -213.145 -79.095 -212.975 -78.925 ;
        RECT -204.165 -79.095 -203.995 -78.925 ;
        RECT -194.245 -78.175 -194.075 -78.005 ;
        RECT -193.775 -78.180 -193.605 -78.010 ;
        RECT -193.305 -78.175 -193.135 -78.005 ;
        RECT -203.225 -78.635 -203.055 -78.465 ;
        RECT -194.245 -78.635 -194.075 -78.465 ;
        RECT -203.225 -79.095 -203.055 -78.925 ;
        RECT -194.245 -79.095 -194.075 -78.925 ;
        RECT -184.325 -78.175 -184.155 -78.005 ;
        RECT -183.855 -78.180 -183.685 -78.010 ;
        RECT -183.385 -78.175 -183.215 -78.005 ;
        RECT -193.305 -78.635 -193.135 -78.465 ;
        RECT -184.325 -78.635 -184.155 -78.465 ;
        RECT -193.305 -79.095 -193.135 -78.925 ;
        RECT -184.325 -79.095 -184.155 -78.925 ;
        RECT -174.405 -78.175 -174.235 -78.005 ;
        RECT -173.935 -78.180 -173.765 -78.010 ;
        RECT -173.465 -78.175 -173.295 -78.005 ;
        RECT -183.385 -78.635 -183.215 -78.465 ;
        RECT -174.405 -78.635 -174.235 -78.465 ;
        RECT -183.385 -79.095 -183.215 -78.925 ;
        RECT -174.405 -79.095 -174.235 -78.925 ;
        RECT -164.485 -78.175 -164.315 -78.005 ;
        RECT -164.015 -78.180 -163.845 -78.010 ;
        RECT -163.545 -78.175 -163.375 -78.005 ;
        RECT -173.465 -78.635 -173.295 -78.465 ;
        RECT -164.485 -78.635 -164.315 -78.465 ;
        RECT -173.465 -79.095 -173.295 -78.925 ;
        RECT -164.485 -79.095 -164.315 -78.925 ;
        RECT -154.565 -78.175 -154.395 -78.005 ;
        RECT -154.095 -78.180 -153.925 -78.010 ;
        RECT -153.625 -78.175 -153.455 -78.005 ;
        RECT -163.545 -78.635 -163.375 -78.465 ;
        RECT -154.565 -78.635 -154.395 -78.465 ;
        RECT -163.545 -79.095 -163.375 -78.925 ;
        RECT -154.565 -79.095 -154.395 -78.925 ;
        RECT -144.645 -78.175 -144.475 -78.005 ;
        RECT -144.175 -78.180 -144.005 -78.010 ;
        RECT -143.705 -78.175 -143.535 -78.005 ;
        RECT -153.625 -78.635 -153.455 -78.465 ;
        RECT -144.645 -78.635 -144.475 -78.465 ;
        RECT -153.625 -79.095 -153.455 -78.925 ;
        RECT -144.645 -79.095 -144.475 -78.925 ;
        RECT -134.725 -78.175 -134.555 -78.005 ;
        RECT -134.255 -78.180 -134.085 -78.010 ;
        RECT -133.785 -78.175 -133.615 -78.005 ;
        RECT -143.705 -78.635 -143.535 -78.465 ;
        RECT -134.725 -78.635 -134.555 -78.465 ;
        RECT -143.705 -79.095 -143.535 -78.925 ;
        RECT -134.725 -79.095 -134.555 -78.925 ;
        RECT -124.805 -78.175 -124.635 -78.005 ;
        RECT -124.335 -78.180 -124.165 -78.010 ;
        RECT -123.865 -78.175 -123.695 -78.005 ;
        RECT -133.785 -78.635 -133.615 -78.465 ;
        RECT -124.805 -78.635 -124.635 -78.465 ;
        RECT -133.785 -79.095 -133.615 -78.925 ;
        RECT -124.805 -79.095 -124.635 -78.925 ;
        RECT -114.885 -78.175 -114.715 -78.005 ;
        RECT -114.415 -78.180 -114.245 -78.010 ;
        RECT -113.945 -78.175 -113.775 -78.005 ;
        RECT -123.865 -78.635 -123.695 -78.465 ;
        RECT -114.885 -78.635 -114.715 -78.465 ;
        RECT -123.865 -79.095 -123.695 -78.925 ;
        RECT -114.885 -79.095 -114.715 -78.925 ;
        RECT -104.965 -78.175 -104.795 -78.005 ;
        RECT -104.495 -78.180 -104.325 -78.010 ;
        RECT -104.025 -78.175 -103.855 -78.005 ;
        RECT -113.945 -78.635 -113.775 -78.465 ;
        RECT -104.965 -78.635 -104.795 -78.465 ;
        RECT -113.945 -79.095 -113.775 -78.925 ;
        RECT -104.965 -79.095 -104.795 -78.925 ;
        RECT -95.045 -78.175 -94.875 -78.005 ;
        RECT -94.575 -78.180 -94.405 -78.010 ;
        RECT -94.105 -78.175 -93.935 -78.005 ;
        RECT -104.025 -78.635 -103.855 -78.465 ;
        RECT -95.045 -78.635 -94.875 -78.465 ;
        RECT -104.025 -79.095 -103.855 -78.925 ;
        RECT -95.045 -79.095 -94.875 -78.925 ;
        RECT -85.125 -78.175 -84.955 -78.005 ;
        RECT -84.655 -78.180 -84.485 -78.010 ;
        RECT -84.185 -78.175 -84.015 -78.005 ;
        RECT -94.105 -78.635 -93.935 -78.465 ;
        RECT -85.125 -78.635 -84.955 -78.465 ;
        RECT -94.105 -79.095 -93.935 -78.925 ;
        RECT -85.125 -79.095 -84.955 -78.925 ;
        RECT -75.205 -78.175 -75.035 -78.005 ;
        RECT -74.735 -78.180 -74.565 -78.010 ;
        RECT -74.265 -78.175 -74.095 -78.005 ;
        RECT -84.185 -78.635 -84.015 -78.465 ;
        RECT -75.205 -78.635 -75.035 -78.465 ;
        RECT -84.185 -79.095 -84.015 -78.925 ;
        RECT -75.205 -79.095 -75.035 -78.925 ;
        RECT -65.285 -78.175 -65.115 -78.005 ;
        RECT -64.815 -78.180 -64.645 -78.010 ;
        RECT -64.345 -78.175 -64.175 -78.005 ;
        RECT -74.265 -78.635 -74.095 -78.465 ;
        RECT -65.285 -78.635 -65.115 -78.465 ;
        RECT -74.265 -79.095 -74.095 -78.925 ;
        RECT -65.285 -79.095 -65.115 -78.925 ;
        RECT -55.365 -78.175 -55.195 -78.005 ;
        RECT -54.895 -78.180 -54.725 -78.010 ;
        RECT -54.425 -78.175 -54.255 -78.005 ;
        RECT -64.345 -78.635 -64.175 -78.465 ;
        RECT -55.365 -78.635 -55.195 -78.465 ;
        RECT -64.345 -79.095 -64.175 -78.925 ;
        RECT -55.365 -79.095 -55.195 -78.925 ;
        RECT -45.445 -78.175 -45.275 -78.005 ;
        RECT -44.975 -78.180 -44.805 -78.010 ;
        RECT -44.505 -78.175 -44.335 -78.005 ;
        RECT -54.425 -78.635 -54.255 -78.465 ;
        RECT -45.445 -78.635 -45.275 -78.465 ;
        RECT -54.425 -79.095 -54.255 -78.925 ;
        RECT -45.445 -79.095 -45.275 -78.925 ;
        RECT -35.525 -78.175 -35.355 -78.005 ;
        RECT -35.055 -78.180 -34.885 -78.010 ;
        RECT -34.585 -78.175 -34.415 -78.005 ;
        RECT -44.505 -78.635 -44.335 -78.465 ;
        RECT -35.525 -78.635 -35.355 -78.465 ;
        RECT -44.505 -79.095 -44.335 -78.925 ;
        RECT -35.525 -79.095 -35.355 -78.925 ;
        RECT -25.605 -78.175 -25.435 -78.005 ;
        RECT -25.135 -78.180 -24.965 -78.010 ;
        RECT -24.665 -78.175 -24.495 -78.005 ;
        RECT -34.585 -78.635 -34.415 -78.465 ;
        RECT -25.605 -78.635 -25.435 -78.465 ;
        RECT -34.585 -79.095 -34.415 -78.925 ;
        RECT -25.605 -79.095 -25.435 -78.925 ;
        RECT -15.685 -78.175 -15.515 -78.005 ;
        RECT -15.215 -78.180 -15.045 -78.010 ;
        RECT -14.745 -78.175 -14.575 -78.005 ;
        RECT -24.665 -78.635 -24.495 -78.465 ;
        RECT -15.685 -78.635 -15.515 -78.465 ;
        RECT -24.665 -79.095 -24.495 -78.925 ;
        RECT -15.685 -79.095 -15.515 -78.925 ;
        RECT -5.765 -78.175 -5.595 -78.005 ;
        RECT -5.295 -78.180 -5.125 -78.010 ;
        RECT -4.825 -78.175 -4.655 -78.005 ;
        RECT -14.745 -78.635 -14.575 -78.465 ;
        RECT -5.765 -78.635 -5.595 -78.465 ;
        RECT -14.745 -79.095 -14.575 -78.925 ;
        RECT -5.765 -79.095 -5.595 -78.925 ;
        RECT 4.155 -78.175 4.325 -78.005 ;
        RECT 4.625 -78.180 4.795 -78.010 ;
        RECT 5.095 -78.175 5.265 -78.005 ;
        RECT -4.825 -78.635 -4.655 -78.465 ;
        RECT 4.155 -78.635 4.325 -78.465 ;
        RECT -4.825 -79.095 -4.655 -78.925 ;
        RECT 4.155 -79.095 4.325 -78.925 ;
        RECT 14.075 -78.175 14.245 -78.005 ;
        RECT 14.545 -78.180 14.715 -78.010 ;
        RECT 15.015 -78.175 15.185 -78.005 ;
        RECT 5.095 -78.635 5.265 -78.465 ;
        RECT 14.075 -78.635 14.245 -78.465 ;
        RECT 5.095 -79.095 5.265 -78.925 ;
        RECT 14.075 -79.095 14.245 -78.925 ;
        RECT 23.995 -78.175 24.165 -78.005 ;
        RECT 24.465 -78.180 24.635 -78.010 ;
        RECT 15.015 -78.635 15.185 -78.465 ;
        RECT 23.995 -78.635 24.165 -78.465 ;
        RECT 15.015 -79.095 15.185 -78.925 ;
        RECT 23.995 -79.095 24.165 -78.925 ;
        RECT -289.395 -79.755 -289.225 -79.585 ;
        RECT -288.935 -79.755 -288.765 -79.585 ;
        RECT -288.475 -79.755 -288.305 -79.585 ;
        RECT -288.015 -79.755 -287.845 -79.585 ;
        RECT -287.555 -79.755 -287.385 -79.585 ;
        RECT -287.095 -79.755 -286.925 -79.585 ;
        RECT -286.635 -79.755 -286.465 -79.585 ;
        RECT -279.475 -79.755 -279.305 -79.585 ;
        RECT -279.015 -79.755 -278.845 -79.585 ;
        RECT -278.555 -79.755 -278.385 -79.585 ;
        RECT -278.095 -79.755 -277.925 -79.585 ;
        RECT -277.635 -79.755 -277.465 -79.585 ;
        RECT -277.175 -79.755 -277.005 -79.585 ;
        RECT -276.715 -79.755 -276.545 -79.585 ;
        RECT -269.555 -79.755 -269.385 -79.585 ;
        RECT -269.095 -79.755 -268.925 -79.585 ;
        RECT -268.635 -79.755 -268.465 -79.585 ;
        RECT -268.175 -79.755 -268.005 -79.585 ;
        RECT -267.715 -79.755 -267.545 -79.585 ;
        RECT -267.255 -79.755 -267.085 -79.585 ;
        RECT -266.795 -79.755 -266.625 -79.585 ;
        RECT -259.635 -79.755 -259.465 -79.585 ;
        RECT -259.175 -79.755 -259.005 -79.585 ;
        RECT -258.715 -79.755 -258.545 -79.585 ;
        RECT -258.255 -79.755 -258.085 -79.585 ;
        RECT -257.795 -79.755 -257.625 -79.585 ;
        RECT -257.335 -79.755 -257.165 -79.585 ;
        RECT -256.875 -79.755 -256.705 -79.585 ;
        RECT -249.715 -79.755 -249.545 -79.585 ;
        RECT -249.255 -79.755 -249.085 -79.585 ;
        RECT -248.795 -79.755 -248.625 -79.585 ;
        RECT -248.335 -79.755 -248.165 -79.585 ;
        RECT -247.875 -79.755 -247.705 -79.585 ;
        RECT -247.415 -79.755 -247.245 -79.585 ;
        RECT -246.955 -79.755 -246.785 -79.585 ;
        RECT -239.795 -79.755 -239.625 -79.585 ;
        RECT -239.335 -79.755 -239.165 -79.585 ;
        RECT -238.875 -79.755 -238.705 -79.585 ;
        RECT -238.415 -79.755 -238.245 -79.585 ;
        RECT -237.955 -79.755 -237.785 -79.585 ;
        RECT -237.495 -79.755 -237.325 -79.585 ;
        RECT -237.035 -79.755 -236.865 -79.585 ;
        RECT -229.875 -79.755 -229.705 -79.585 ;
        RECT -229.415 -79.755 -229.245 -79.585 ;
        RECT -228.955 -79.755 -228.785 -79.585 ;
        RECT -228.495 -79.755 -228.325 -79.585 ;
        RECT -228.035 -79.755 -227.865 -79.585 ;
        RECT -227.575 -79.755 -227.405 -79.585 ;
        RECT -227.115 -79.755 -226.945 -79.585 ;
        RECT -219.955 -79.755 -219.785 -79.585 ;
        RECT -219.495 -79.755 -219.325 -79.585 ;
        RECT -219.035 -79.755 -218.865 -79.585 ;
        RECT -218.575 -79.755 -218.405 -79.585 ;
        RECT -218.115 -79.755 -217.945 -79.585 ;
        RECT -217.655 -79.755 -217.485 -79.585 ;
        RECT -217.195 -79.755 -217.025 -79.585 ;
        RECT -210.035 -79.755 -209.865 -79.585 ;
        RECT -209.575 -79.755 -209.405 -79.585 ;
        RECT -209.115 -79.755 -208.945 -79.585 ;
        RECT -208.655 -79.755 -208.485 -79.585 ;
        RECT -208.195 -79.755 -208.025 -79.585 ;
        RECT -207.735 -79.755 -207.565 -79.585 ;
        RECT -207.275 -79.755 -207.105 -79.585 ;
        RECT -200.115 -79.755 -199.945 -79.585 ;
        RECT -199.655 -79.755 -199.485 -79.585 ;
        RECT -199.195 -79.755 -199.025 -79.585 ;
        RECT -198.735 -79.755 -198.565 -79.585 ;
        RECT -198.275 -79.755 -198.105 -79.585 ;
        RECT -197.815 -79.755 -197.645 -79.585 ;
        RECT -197.355 -79.755 -197.185 -79.585 ;
        RECT -190.195 -79.755 -190.025 -79.585 ;
        RECT -189.735 -79.755 -189.565 -79.585 ;
        RECT -189.275 -79.755 -189.105 -79.585 ;
        RECT -188.815 -79.755 -188.645 -79.585 ;
        RECT -188.355 -79.755 -188.185 -79.585 ;
        RECT -187.895 -79.755 -187.725 -79.585 ;
        RECT -187.435 -79.755 -187.265 -79.585 ;
        RECT -180.275 -79.755 -180.105 -79.585 ;
        RECT -179.815 -79.755 -179.645 -79.585 ;
        RECT -179.355 -79.755 -179.185 -79.585 ;
        RECT -178.895 -79.755 -178.725 -79.585 ;
        RECT -178.435 -79.755 -178.265 -79.585 ;
        RECT -177.975 -79.755 -177.805 -79.585 ;
        RECT -177.515 -79.755 -177.345 -79.585 ;
        RECT -170.355 -79.755 -170.185 -79.585 ;
        RECT -169.895 -79.755 -169.725 -79.585 ;
        RECT -169.435 -79.755 -169.265 -79.585 ;
        RECT -168.975 -79.755 -168.805 -79.585 ;
        RECT -168.515 -79.755 -168.345 -79.585 ;
        RECT -168.055 -79.755 -167.885 -79.585 ;
        RECT -167.595 -79.755 -167.425 -79.585 ;
        RECT -160.435 -79.755 -160.265 -79.585 ;
        RECT -159.975 -79.755 -159.805 -79.585 ;
        RECT -159.515 -79.755 -159.345 -79.585 ;
        RECT -159.055 -79.755 -158.885 -79.585 ;
        RECT -158.595 -79.755 -158.425 -79.585 ;
        RECT -158.135 -79.755 -157.965 -79.585 ;
        RECT -157.675 -79.755 -157.505 -79.585 ;
        RECT -150.515 -79.755 -150.345 -79.585 ;
        RECT -150.055 -79.755 -149.885 -79.585 ;
        RECT -149.595 -79.755 -149.425 -79.585 ;
        RECT -149.135 -79.755 -148.965 -79.585 ;
        RECT -148.675 -79.755 -148.505 -79.585 ;
        RECT -148.215 -79.755 -148.045 -79.585 ;
        RECT -147.755 -79.755 -147.585 -79.585 ;
        RECT -140.595 -79.755 -140.425 -79.585 ;
        RECT -140.135 -79.755 -139.965 -79.585 ;
        RECT -139.675 -79.755 -139.505 -79.585 ;
        RECT -139.215 -79.755 -139.045 -79.585 ;
        RECT -138.755 -79.755 -138.585 -79.585 ;
        RECT -138.295 -79.755 -138.125 -79.585 ;
        RECT -137.835 -79.755 -137.665 -79.585 ;
        RECT -130.675 -79.755 -130.505 -79.585 ;
        RECT -130.215 -79.755 -130.045 -79.585 ;
        RECT -129.755 -79.755 -129.585 -79.585 ;
        RECT -129.295 -79.755 -129.125 -79.585 ;
        RECT -128.835 -79.755 -128.665 -79.585 ;
        RECT -128.375 -79.755 -128.205 -79.585 ;
        RECT -127.915 -79.755 -127.745 -79.585 ;
        RECT -120.755 -79.755 -120.585 -79.585 ;
        RECT -120.295 -79.755 -120.125 -79.585 ;
        RECT -119.835 -79.755 -119.665 -79.585 ;
        RECT -119.375 -79.755 -119.205 -79.585 ;
        RECT -118.915 -79.755 -118.745 -79.585 ;
        RECT -118.455 -79.755 -118.285 -79.585 ;
        RECT -117.995 -79.755 -117.825 -79.585 ;
        RECT -110.835 -79.755 -110.665 -79.585 ;
        RECT -110.375 -79.755 -110.205 -79.585 ;
        RECT -109.915 -79.755 -109.745 -79.585 ;
        RECT -109.455 -79.755 -109.285 -79.585 ;
        RECT -108.995 -79.755 -108.825 -79.585 ;
        RECT -108.535 -79.755 -108.365 -79.585 ;
        RECT -108.075 -79.755 -107.905 -79.585 ;
        RECT -100.915 -79.755 -100.745 -79.585 ;
        RECT -100.455 -79.755 -100.285 -79.585 ;
        RECT -99.995 -79.755 -99.825 -79.585 ;
        RECT -99.535 -79.755 -99.365 -79.585 ;
        RECT -99.075 -79.755 -98.905 -79.585 ;
        RECT -98.615 -79.755 -98.445 -79.585 ;
        RECT -98.155 -79.755 -97.985 -79.585 ;
        RECT -90.995 -79.755 -90.825 -79.585 ;
        RECT -90.535 -79.755 -90.365 -79.585 ;
        RECT -90.075 -79.755 -89.905 -79.585 ;
        RECT -89.615 -79.755 -89.445 -79.585 ;
        RECT -89.155 -79.755 -88.985 -79.585 ;
        RECT -88.695 -79.755 -88.525 -79.585 ;
        RECT -88.235 -79.755 -88.065 -79.585 ;
        RECT -81.075 -79.755 -80.905 -79.585 ;
        RECT -80.615 -79.755 -80.445 -79.585 ;
        RECT -80.155 -79.755 -79.985 -79.585 ;
        RECT -79.695 -79.755 -79.525 -79.585 ;
        RECT -79.235 -79.755 -79.065 -79.585 ;
        RECT -78.775 -79.755 -78.605 -79.585 ;
        RECT -78.315 -79.755 -78.145 -79.585 ;
        RECT -71.155 -79.755 -70.985 -79.585 ;
        RECT -70.695 -79.755 -70.525 -79.585 ;
        RECT -70.235 -79.755 -70.065 -79.585 ;
        RECT -69.775 -79.755 -69.605 -79.585 ;
        RECT -69.315 -79.755 -69.145 -79.585 ;
        RECT -68.855 -79.755 -68.685 -79.585 ;
        RECT -68.395 -79.755 -68.225 -79.585 ;
        RECT -61.235 -79.755 -61.065 -79.585 ;
        RECT -60.775 -79.755 -60.605 -79.585 ;
        RECT -60.315 -79.755 -60.145 -79.585 ;
        RECT -59.855 -79.755 -59.685 -79.585 ;
        RECT -59.395 -79.755 -59.225 -79.585 ;
        RECT -58.935 -79.755 -58.765 -79.585 ;
        RECT -58.475 -79.755 -58.305 -79.585 ;
        RECT -51.315 -79.755 -51.145 -79.585 ;
        RECT -50.855 -79.755 -50.685 -79.585 ;
        RECT -50.395 -79.755 -50.225 -79.585 ;
        RECT -49.935 -79.755 -49.765 -79.585 ;
        RECT -49.475 -79.755 -49.305 -79.585 ;
        RECT -49.015 -79.755 -48.845 -79.585 ;
        RECT -48.555 -79.755 -48.385 -79.585 ;
        RECT -41.395 -79.755 -41.225 -79.585 ;
        RECT -40.935 -79.755 -40.765 -79.585 ;
        RECT -40.475 -79.755 -40.305 -79.585 ;
        RECT -40.015 -79.755 -39.845 -79.585 ;
        RECT -39.555 -79.755 -39.385 -79.585 ;
        RECT -39.095 -79.755 -38.925 -79.585 ;
        RECT -38.635 -79.755 -38.465 -79.585 ;
        RECT -31.475 -79.755 -31.305 -79.585 ;
        RECT -31.015 -79.755 -30.845 -79.585 ;
        RECT -30.555 -79.755 -30.385 -79.585 ;
        RECT -30.095 -79.755 -29.925 -79.585 ;
        RECT -29.635 -79.755 -29.465 -79.585 ;
        RECT -29.175 -79.755 -29.005 -79.585 ;
        RECT -28.715 -79.755 -28.545 -79.585 ;
        RECT -21.555 -79.755 -21.385 -79.585 ;
        RECT -21.095 -79.755 -20.925 -79.585 ;
        RECT -20.635 -79.755 -20.465 -79.585 ;
        RECT -20.175 -79.755 -20.005 -79.585 ;
        RECT -19.715 -79.755 -19.545 -79.585 ;
        RECT -19.255 -79.755 -19.085 -79.585 ;
        RECT -18.795 -79.755 -18.625 -79.585 ;
        RECT -11.635 -79.755 -11.465 -79.585 ;
        RECT -11.175 -79.755 -11.005 -79.585 ;
        RECT -10.715 -79.755 -10.545 -79.585 ;
        RECT -10.255 -79.755 -10.085 -79.585 ;
        RECT -9.795 -79.755 -9.625 -79.585 ;
        RECT -9.335 -79.755 -9.165 -79.585 ;
        RECT -8.875 -79.755 -8.705 -79.585 ;
        RECT -1.715 -79.755 -1.545 -79.585 ;
        RECT -1.255 -79.755 -1.085 -79.585 ;
        RECT -0.795 -79.755 -0.625 -79.585 ;
        RECT -0.335 -79.755 -0.165 -79.585 ;
        RECT 0.125 -79.755 0.295 -79.585 ;
        RECT 0.585 -79.755 0.755 -79.585 ;
        RECT 1.045 -79.755 1.215 -79.585 ;
        RECT 8.205 -79.755 8.375 -79.585 ;
        RECT 8.665 -79.755 8.835 -79.585 ;
        RECT 9.125 -79.755 9.295 -79.585 ;
        RECT 9.585 -79.755 9.755 -79.585 ;
        RECT 10.045 -79.755 10.215 -79.585 ;
        RECT 10.505 -79.755 10.675 -79.585 ;
        RECT 10.965 -79.755 11.135 -79.585 ;
        RECT 18.125 -79.755 18.295 -79.585 ;
        RECT 18.585 -79.755 18.755 -79.585 ;
        RECT 19.045 -79.755 19.215 -79.585 ;
        RECT 19.505 -79.755 19.675 -79.585 ;
        RECT 19.965 -79.755 20.135 -79.585 ;
        RECT 20.425 -79.755 20.595 -79.585 ;
        RECT 20.885 -79.755 21.055 -79.585 ;
        RECT -284.435 -82.475 -284.265 -82.305 ;
        RECT -283.975 -82.475 -283.805 -82.305 ;
        RECT -283.515 -82.475 -283.345 -82.305 ;
        RECT -283.055 -82.475 -282.885 -82.305 ;
        RECT -282.595 -82.475 -282.425 -82.305 ;
        RECT -282.135 -82.475 -281.965 -82.305 ;
        RECT -281.675 -82.475 -281.505 -82.305 ;
        RECT -274.515 -82.475 -274.345 -82.305 ;
        RECT -274.055 -82.475 -273.885 -82.305 ;
        RECT -273.595 -82.475 -273.425 -82.305 ;
        RECT -273.135 -82.475 -272.965 -82.305 ;
        RECT -272.675 -82.475 -272.505 -82.305 ;
        RECT -272.215 -82.475 -272.045 -82.305 ;
        RECT -271.755 -82.475 -271.585 -82.305 ;
        RECT -264.595 -82.475 -264.425 -82.305 ;
        RECT -264.135 -82.475 -263.965 -82.305 ;
        RECT -263.675 -82.475 -263.505 -82.305 ;
        RECT -263.215 -82.475 -263.045 -82.305 ;
        RECT -262.755 -82.475 -262.585 -82.305 ;
        RECT -262.295 -82.475 -262.125 -82.305 ;
        RECT -261.835 -82.475 -261.665 -82.305 ;
        RECT -254.675 -82.475 -254.505 -82.305 ;
        RECT -254.215 -82.475 -254.045 -82.305 ;
        RECT -253.755 -82.475 -253.585 -82.305 ;
        RECT -253.295 -82.475 -253.125 -82.305 ;
        RECT -252.835 -82.475 -252.665 -82.305 ;
        RECT -252.375 -82.475 -252.205 -82.305 ;
        RECT -251.915 -82.475 -251.745 -82.305 ;
        RECT -244.755 -82.475 -244.585 -82.305 ;
        RECT -244.295 -82.475 -244.125 -82.305 ;
        RECT -243.835 -82.475 -243.665 -82.305 ;
        RECT -243.375 -82.475 -243.205 -82.305 ;
        RECT -242.915 -82.475 -242.745 -82.305 ;
        RECT -242.455 -82.475 -242.285 -82.305 ;
        RECT -241.995 -82.475 -241.825 -82.305 ;
        RECT -234.835 -82.475 -234.665 -82.305 ;
        RECT -234.375 -82.475 -234.205 -82.305 ;
        RECT -233.915 -82.475 -233.745 -82.305 ;
        RECT -233.455 -82.475 -233.285 -82.305 ;
        RECT -232.995 -82.475 -232.825 -82.305 ;
        RECT -232.535 -82.475 -232.365 -82.305 ;
        RECT -232.075 -82.475 -231.905 -82.305 ;
        RECT -224.915 -82.475 -224.745 -82.305 ;
        RECT -224.455 -82.475 -224.285 -82.305 ;
        RECT -223.995 -82.475 -223.825 -82.305 ;
        RECT -223.535 -82.475 -223.365 -82.305 ;
        RECT -223.075 -82.475 -222.905 -82.305 ;
        RECT -222.615 -82.475 -222.445 -82.305 ;
        RECT -222.155 -82.475 -221.985 -82.305 ;
        RECT -214.995 -82.475 -214.825 -82.305 ;
        RECT -214.535 -82.475 -214.365 -82.305 ;
        RECT -214.075 -82.475 -213.905 -82.305 ;
        RECT -213.615 -82.475 -213.445 -82.305 ;
        RECT -213.155 -82.475 -212.985 -82.305 ;
        RECT -212.695 -82.475 -212.525 -82.305 ;
        RECT -212.235 -82.475 -212.065 -82.305 ;
        RECT -205.075 -82.475 -204.905 -82.305 ;
        RECT -204.615 -82.475 -204.445 -82.305 ;
        RECT -204.155 -82.475 -203.985 -82.305 ;
        RECT -203.695 -82.475 -203.525 -82.305 ;
        RECT -203.235 -82.475 -203.065 -82.305 ;
        RECT -202.775 -82.475 -202.605 -82.305 ;
        RECT -202.315 -82.475 -202.145 -82.305 ;
        RECT -195.155 -82.475 -194.985 -82.305 ;
        RECT -194.695 -82.475 -194.525 -82.305 ;
        RECT -194.235 -82.475 -194.065 -82.305 ;
        RECT -193.775 -82.475 -193.605 -82.305 ;
        RECT -193.315 -82.475 -193.145 -82.305 ;
        RECT -192.855 -82.475 -192.685 -82.305 ;
        RECT -192.395 -82.475 -192.225 -82.305 ;
        RECT -185.235 -82.475 -185.065 -82.305 ;
        RECT -184.775 -82.475 -184.605 -82.305 ;
        RECT -184.315 -82.475 -184.145 -82.305 ;
        RECT -183.855 -82.475 -183.685 -82.305 ;
        RECT -183.395 -82.475 -183.225 -82.305 ;
        RECT -182.935 -82.475 -182.765 -82.305 ;
        RECT -182.475 -82.475 -182.305 -82.305 ;
        RECT -175.315 -82.475 -175.145 -82.305 ;
        RECT -174.855 -82.475 -174.685 -82.305 ;
        RECT -174.395 -82.475 -174.225 -82.305 ;
        RECT -173.935 -82.475 -173.765 -82.305 ;
        RECT -173.475 -82.475 -173.305 -82.305 ;
        RECT -173.015 -82.475 -172.845 -82.305 ;
        RECT -172.555 -82.475 -172.385 -82.305 ;
        RECT -165.395 -82.475 -165.225 -82.305 ;
        RECT -164.935 -82.475 -164.765 -82.305 ;
        RECT -164.475 -82.475 -164.305 -82.305 ;
        RECT -164.015 -82.475 -163.845 -82.305 ;
        RECT -163.555 -82.475 -163.385 -82.305 ;
        RECT -163.095 -82.475 -162.925 -82.305 ;
        RECT -162.635 -82.475 -162.465 -82.305 ;
        RECT -155.475 -82.475 -155.305 -82.305 ;
        RECT -155.015 -82.475 -154.845 -82.305 ;
        RECT -154.555 -82.475 -154.385 -82.305 ;
        RECT -154.095 -82.475 -153.925 -82.305 ;
        RECT -153.635 -82.475 -153.465 -82.305 ;
        RECT -153.175 -82.475 -153.005 -82.305 ;
        RECT -152.715 -82.475 -152.545 -82.305 ;
        RECT -145.555 -82.475 -145.385 -82.305 ;
        RECT -145.095 -82.475 -144.925 -82.305 ;
        RECT -144.635 -82.475 -144.465 -82.305 ;
        RECT -144.175 -82.475 -144.005 -82.305 ;
        RECT -143.715 -82.475 -143.545 -82.305 ;
        RECT -143.255 -82.475 -143.085 -82.305 ;
        RECT -142.795 -82.475 -142.625 -82.305 ;
        RECT -135.635 -82.475 -135.465 -82.305 ;
        RECT -135.175 -82.475 -135.005 -82.305 ;
        RECT -134.715 -82.475 -134.545 -82.305 ;
        RECT -134.255 -82.475 -134.085 -82.305 ;
        RECT -133.795 -82.475 -133.625 -82.305 ;
        RECT -133.335 -82.475 -133.165 -82.305 ;
        RECT -132.875 -82.475 -132.705 -82.305 ;
        RECT -125.715 -82.475 -125.545 -82.305 ;
        RECT -125.255 -82.475 -125.085 -82.305 ;
        RECT -124.795 -82.475 -124.625 -82.305 ;
        RECT -124.335 -82.475 -124.165 -82.305 ;
        RECT -123.875 -82.475 -123.705 -82.305 ;
        RECT -123.415 -82.475 -123.245 -82.305 ;
        RECT -122.955 -82.475 -122.785 -82.305 ;
        RECT -115.795 -82.475 -115.625 -82.305 ;
        RECT -115.335 -82.475 -115.165 -82.305 ;
        RECT -114.875 -82.475 -114.705 -82.305 ;
        RECT -114.415 -82.475 -114.245 -82.305 ;
        RECT -113.955 -82.475 -113.785 -82.305 ;
        RECT -113.495 -82.475 -113.325 -82.305 ;
        RECT -113.035 -82.475 -112.865 -82.305 ;
        RECT -105.875 -82.475 -105.705 -82.305 ;
        RECT -105.415 -82.475 -105.245 -82.305 ;
        RECT -104.955 -82.475 -104.785 -82.305 ;
        RECT -104.495 -82.475 -104.325 -82.305 ;
        RECT -104.035 -82.475 -103.865 -82.305 ;
        RECT -103.575 -82.475 -103.405 -82.305 ;
        RECT -103.115 -82.475 -102.945 -82.305 ;
        RECT -95.955 -82.475 -95.785 -82.305 ;
        RECT -95.495 -82.475 -95.325 -82.305 ;
        RECT -95.035 -82.475 -94.865 -82.305 ;
        RECT -94.575 -82.475 -94.405 -82.305 ;
        RECT -94.115 -82.475 -93.945 -82.305 ;
        RECT -93.655 -82.475 -93.485 -82.305 ;
        RECT -93.195 -82.475 -93.025 -82.305 ;
        RECT -86.035 -82.475 -85.865 -82.305 ;
        RECT -85.575 -82.475 -85.405 -82.305 ;
        RECT -85.115 -82.475 -84.945 -82.305 ;
        RECT -84.655 -82.475 -84.485 -82.305 ;
        RECT -84.195 -82.475 -84.025 -82.305 ;
        RECT -83.735 -82.475 -83.565 -82.305 ;
        RECT -83.275 -82.475 -83.105 -82.305 ;
        RECT -76.115 -82.475 -75.945 -82.305 ;
        RECT -75.655 -82.475 -75.485 -82.305 ;
        RECT -75.195 -82.475 -75.025 -82.305 ;
        RECT -74.735 -82.475 -74.565 -82.305 ;
        RECT -74.275 -82.475 -74.105 -82.305 ;
        RECT -73.815 -82.475 -73.645 -82.305 ;
        RECT -73.355 -82.475 -73.185 -82.305 ;
        RECT -66.195 -82.475 -66.025 -82.305 ;
        RECT -65.735 -82.475 -65.565 -82.305 ;
        RECT -65.275 -82.475 -65.105 -82.305 ;
        RECT -64.815 -82.475 -64.645 -82.305 ;
        RECT -64.355 -82.475 -64.185 -82.305 ;
        RECT -63.895 -82.475 -63.725 -82.305 ;
        RECT -63.435 -82.475 -63.265 -82.305 ;
        RECT -56.275 -82.475 -56.105 -82.305 ;
        RECT -55.815 -82.475 -55.645 -82.305 ;
        RECT -55.355 -82.475 -55.185 -82.305 ;
        RECT -54.895 -82.475 -54.725 -82.305 ;
        RECT -54.435 -82.475 -54.265 -82.305 ;
        RECT -53.975 -82.475 -53.805 -82.305 ;
        RECT -53.515 -82.475 -53.345 -82.305 ;
        RECT -46.355 -82.475 -46.185 -82.305 ;
        RECT -45.895 -82.475 -45.725 -82.305 ;
        RECT -45.435 -82.475 -45.265 -82.305 ;
        RECT -44.975 -82.475 -44.805 -82.305 ;
        RECT -44.515 -82.475 -44.345 -82.305 ;
        RECT -44.055 -82.475 -43.885 -82.305 ;
        RECT -43.595 -82.475 -43.425 -82.305 ;
        RECT -36.435 -82.475 -36.265 -82.305 ;
        RECT -35.975 -82.475 -35.805 -82.305 ;
        RECT -35.515 -82.475 -35.345 -82.305 ;
        RECT -35.055 -82.475 -34.885 -82.305 ;
        RECT -34.595 -82.475 -34.425 -82.305 ;
        RECT -34.135 -82.475 -33.965 -82.305 ;
        RECT -33.675 -82.475 -33.505 -82.305 ;
        RECT -26.515 -82.475 -26.345 -82.305 ;
        RECT -26.055 -82.475 -25.885 -82.305 ;
        RECT -25.595 -82.475 -25.425 -82.305 ;
        RECT -25.135 -82.475 -24.965 -82.305 ;
        RECT -24.675 -82.475 -24.505 -82.305 ;
        RECT -24.215 -82.475 -24.045 -82.305 ;
        RECT -23.755 -82.475 -23.585 -82.305 ;
        RECT -16.595 -82.475 -16.425 -82.305 ;
        RECT -16.135 -82.475 -15.965 -82.305 ;
        RECT -15.675 -82.475 -15.505 -82.305 ;
        RECT -15.215 -82.475 -15.045 -82.305 ;
        RECT -14.755 -82.475 -14.585 -82.305 ;
        RECT -14.295 -82.475 -14.125 -82.305 ;
        RECT -13.835 -82.475 -13.665 -82.305 ;
        RECT -6.675 -82.475 -6.505 -82.305 ;
        RECT -6.215 -82.475 -6.045 -82.305 ;
        RECT -5.755 -82.475 -5.585 -82.305 ;
        RECT -5.295 -82.475 -5.125 -82.305 ;
        RECT -4.835 -82.475 -4.665 -82.305 ;
        RECT -4.375 -82.475 -4.205 -82.305 ;
        RECT -3.915 -82.475 -3.745 -82.305 ;
        RECT 3.245 -82.475 3.415 -82.305 ;
        RECT 3.705 -82.475 3.875 -82.305 ;
        RECT 4.165 -82.475 4.335 -82.305 ;
        RECT 4.625 -82.475 4.795 -82.305 ;
        RECT 5.085 -82.475 5.255 -82.305 ;
        RECT 5.545 -82.475 5.715 -82.305 ;
        RECT 6.005 -82.475 6.175 -82.305 ;
        RECT 13.165 -82.475 13.335 -82.305 ;
        RECT 13.625 -82.475 13.795 -82.305 ;
        RECT 14.085 -82.475 14.255 -82.305 ;
        RECT 14.545 -82.475 14.715 -82.305 ;
        RECT 15.005 -82.475 15.175 -82.305 ;
        RECT 15.465 -82.475 15.635 -82.305 ;
        RECT 15.925 -82.475 16.095 -82.305 ;
        RECT 23.085 -82.475 23.255 -82.305 ;
        RECT 23.545 -82.475 23.715 -82.305 ;
        RECT 24.005 -82.475 24.175 -82.305 ;
        RECT 24.465 -82.475 24.635 -82.305 ;
        RECT -288.485 -83.135 -288.315 -82.965 ;
        RECT -288.015 -83.060 -287.845 -82.890 ;
        RECT -288.485 -83.595 -288.315 -83.425 ;
        RECT -288.485 -84.055 -288.315 -83.885 ;
        RECT -287.545 -83.135 -287.375 -82.965 ;
        RECT -278.565 -83.135 -278.395 -82.965 ;
        RECT -278.095 -83.060 -277.925 -82.890 ;
        RECT -287.545 -83.595 -287.375 -83.425 ;
        RECT -278.565 -83.595 -278.395 -83.425 ;
        RECT -287.545 -84.055 -287.375 -83.885 ;
        RECT -278.565 -84.055 -278.395 -83.885 ;
        RECT -277.625 -83.135 -277.455 -82.965 ;
        RECT -268.645 -83.135 -268.475 -82.965 ;
        RECT -268.175 -83.060 -268.005 -82.890 ;
        RECT -277.625 -83.595 -277.455 -83.425 ;
        RECT -268.645 -83.595 -268.475 -83.425 ;
        RECT -277.625 -84.055 -277.455 -83.885 ;
        RECT -268.645 -84.055 -268.475 -83.885 ;
        RECT -267.705 -83.135 -267.535 -82.965 ;
        RECT -258.725 -83.135 -258.555 -82.965 ;
        RECT -258.255 -83.060 -258.085 -82.890 ;
        RECT -267.705 -83.595 -267.535 -83.425 ;
        RECT -258.725 -83.595 -258.555 -83.425 ;
        RECT -267.705 -84.055 -267.535 -83.885 ;
        RECT -258.725 -84.055 -258.555 -83.885 ;
        RECT -257.785 -83.135 -257.615 -82.965 ;
        RECT -248.805 -83.135 -248.635 -82.965 ;
        RECT -248.335 -83.060 -248.165 -82.890 ;
        RECT -257.785 -83.595 -257.615 -83.425 ;
        RECT -248.805 -83.595 -248.635 -83.425 ;
        RECT -257.785 -84.055 -257.615 -83.885 ;
        RECT -248.805 -84.055 -248.635 -83.885 ;
        RECT -247.865 -83.135 -247.695 -82.965 ;
        RECT -238.885 -83.135 -238.715 -82.965 ;
        RECT -238.415 -83.060 -238.245 -82.890 ;
        RECT -247.865 -83.595 -247.695 -83.425 ;
        RECT -238.885 -83.595 -238.715 -83.425 ;
        RECT -247.865 -84.055 -247.695 -83.885 ;
        RECT -238.885 -84.055 -238.715 -83.885 ;
        RECT -237.945 -83.135 -237.775 -82.965 ;
        RECT -228.965 -83.135 -228.795 -82.965 ;
        RECT -228.495 -83.060 -228.325 -82.890 ;
        RECT -237.945 -83.595 -237.775 -83.425 ;
        RECT -228.965 -83.595 -228.795 -83.425 ;
        RECT -237.945 -84.055 -237.775 -83.885 ;
        RECT -228.965 -84.055 -228.795 -83.885 ;
        RECT -228.025 -83.135 -227.855 -82.965 ;
        RECT -219.045 -83.135 -218.875 -82.965 ;
        RECT -218.575 -83.060 -218.405 -82.890 ;
        RECT -228.025 -83.595 -227.855 -83.425 ;
        RECT -219.045 -83.595 -218.875 -83.425 ;
        RECT -228.025 -84.055 -227.855 -83.885 ;
        RECT -219.045 -84.055 -218.875 -83.885 ;
        RECT -218.105 -83.135 -217.935 -82.965 ;
        RECT -209.125 -83.135 -208.955 -82.965 ;
        RECT -208.655 -83.060 -208.485 -82.890 ;
        RECT -218.105 -83.595 -217.935 -83.425 ;
        RECT -209.125 -83.595 -208.955 -83.425 ;
        RECT -218.105 -84.055 -217.935 -83.885 ;
        RECT -209.125 -84.055 -208.955 -83.885 ;
        RECT -208.185 -83.135 -208.015 -82.965 ;
        RECT -199.205 -83.135 -199.035 -82.965 ;
        RECT -198.735 -83.060 -198.565 -82.890 ;
        RECT -208.185 -83.595 -208.015 -83.425 ;
        RECT -199.205 -83.595 -199.035 -83.425 ;
        RECT -208.185 -84.055 -208.015 -83.885 ;
        RECT -199.205 -84.055 -199.035 -83.885 ;
        RECT -198.265 -83.135 -198.095 -82.965 ;
        RECT -189.285 -83.135 -189.115 -82.965 ;
        RECT -188.815 -83.060 -188.645 -82.890 ;
        RECT -198.265 -83.595 -198.095 -83.425 ;
        RECT -189.285 -83.595 -189.115 -83.425 ;
        RECT -198.265 -84.055 -198.095 -83.885 ;
        RECT -189.285 -84.055 -189.115 -83.885 ;
        RECT -188.345 -83.135 -188.175 -82.965 ;
        RECT -179.365 -83.135 -179.195 -82.965 ;
        RECT -178.895 -83.060 -178.725 -82.890 ;
        RECT -188.345 -83.595 -188.175 -83.425 ;
        RECT -179.365 -83.595 -179.195 -83.425 ;
        RECT -188.345 -84.055 -188.175 -83.885 ;
        RECT -179.365 -84.055 -179.195 -83.885 ;
        RECT -178.425 -83.135 -178.255 -82.965 ;
        RECT -169.445 -83.135 -169.275 -82.965 ;
        RECT -168.975 -83.060 -168.805 -82.890 ;
        RECT -178.425 -83.595 -178.255 -83.425 ;
        RECT -169.445 -83.595 -169.275 -83.425 ;
        RECT -178.425 -84.055 -178.255 -83.885 ;
        RECT -169.445 -84.055 -169.275 -83.885 ;
        RECT -168.505 -83.135 -168.335 -82.965 ;
        RECT -159.525 -83.135 -159.355 -82.965 ;
        RECT -159.055 -83.060 -158.885 -82.890 ;
        RECT -168.505 -83.595 -168.335 -83.425 ;
        RECT -159.525 -83.595 -159.355 -83.425 ;
        RECT -168.505 -84.055 -168.335 -83.885 ;
        RECT -159.525 -84.055 -159.355 -83.885 ;
        RECT -158.585 -83.135 -158.415 -82.965 ;
        RECT -149.605 -83.135 -149.435 -82.965 ;
        RECT -149.135 -83.060 -148.965 -82.890 ;
        RECT -158.585 -83.595 -158.415 -83.425 ;
        RECT -149.605 -83.595 -149.435 -83.425 ;
        RECT -158.585 -84.055 -158.415 -83.885 ;
        RECT -149.605 -84.055 -149.435 -83.885 ;
        RECT -148.665 -83.135 -148.495 -82.965 ;
        RECT -139.685 -83.135 -139.515 -82.965 ;
        RECT -139.215 -83.060 -139.045 -82.890 ;
        RECT -148.665 -83.595 -148.495 -83.425 ;
        RECT -139.685 -83.595 -139.515 -83.425 ;
        RECT -148.665 -84.055 -148.495 -83.885 ;
        RECT -139.685 -84.055 -139.515 -83.885 ;
        RECT -138.745 -83.135 -138.575 -82.965 ;
        RECT -129.765 -83.135 -129.595 -82.965 ;
        RECT -129.295 -83.060 -129.125 -82.890 ;
        RECT -138.745 -83.595 -138.575 -83.425 ;
        RECT -129.765 -83.595 -129.595 -83.425 ;
        RECT -138.745 -84.055 -138.575 -83.885 ;
        RECT -129.765 -84.055 -129.595 -83.885 ;
        RECT -128.825 -83.135 -128.655 -82.965 ;
        RECT -119.845 -83.135 -119.675 -82.965 ;
        RECT -119.375 -83.060 -119.205 -82.890 ;
        RECT -128.825 -83.595 -128.655 -83.425 ;
        RECT -119.845 -83.595 -119.675 -83.425 ;
        RECT -128.825 -84.055 -128.655 -83.885 ;
        RECT -119.845 -84.055 -119.675 -83.885 ;
        RECT -118.905 -83.135 -118.735 -82.965 ;
        RECT -109.925 -83.135 -109.755 -82.965 ;
        RECT -109.455 -83.060 -109.285 -82.890 ;
        RECT -118.905 -83.595 -118.735 -83.425 ;
        RECT -109.925 -83.595 -109.755 -83.425 ;
        RECT -118.905 -84.055 -118.735 -83.885 ;
        RECT -109.925 -84.055 -109.755 -83.885 ;
        RECT -108.985 -83.135 -108.815 -82.965 ;
        RECT -100.005 -83.135 -99.835 -82.965 ;
        RECT -99.535 -83.060 -99.365 -82.890 ;
        RECT -108.985 -83.595 -108.815 -83.425 ;
        RECT -100.005 -83.595 -99.835 -83.425 ;
        RECT -108.985 -84.055 -108.815 -83.885 ;
        RECT -100.005 -84.055 -99.835 -83.885 ;
        RECT -99.065 -83.135 -98.895 -82.965 ;
        RECT -90.085 -83.135 -89.915 -82.965 ;
        RECT -89.615 -83.060 -89.445 -82.890 ;
        RECT -99.065 -83.595 -98.895 -83.425 ;
        RECT -90.085 -83.595 -89.915 -83.425 ;
        RECT -99.065 -84.055 -98.895 -83.885 ;
        RECT -90.085 -84.055 -89.915 -83.885 ;
        RECT -89.145 -83.135 -88.975 -82.965 ;
        RECT -80.165 -83.135 -79.995 -82.965 ;
        RECT -79.695 -83.060 -79.525 -82.890 ;
        RECT -89.145 -83.595 -88.975 -83.425 ;
        RECT -80.165 -83.595 -79.995 -83.425 ;
        RECT -89.145 -84.055 -88.975 -83.885 ;
        RECT -80.165 -84.055 -79.995 -83.885 ;
        RECT -79.225 -83.135 -79.055 -82.965 ;
        RECT -70.245 -83.135 -70.075 -82.965 ;
        RECT -69.775 -83.060 -69.605 -82.890 ;
        RECT -79.225 -83.595 -79.055 -83.425 ;
        RECT -70.245 -83.595 -70.075 -83.425 ;
        RECT -79.225 -84.055 -79.055 -83.885 ;
        RECT -70.245 -84.055 -70.075 -83.885 ;
        RECT -69.305 -83.135 -69.135 -82.965 ;
        RECT -60.325 -83.135 -60.155 -82.965 ;
        RECT -59.855 -83.060 -59.685 -82.890 ;
        RECT -69.305 -83.595 -69.135 -83.425 ;
        RECT -60.325 -83.595 -60.155 -83.425 ;
        RECT -69.305 -84.055 -69.135 -83.885 ;
        RECT -60.325 -84.055 -60.155 -83.885 ;
        RECT -59.385 -83.135 -59.215 -82.965 ;
        RECT -50.405 -83.135 -50.235 -82.965 ;
        RECT -49.935 -83.060 -49.765 -82.890 ;
        RECT -59.385 -83.595 -59.215 -83.425 ;
        RECT -50.405 -83.595 -50.235 -83.425 ;
        RECT -59.385 -84.055 -59.215 -83.885 ;
        RECT -50.405 -84.055 -50.235 -83.885 ;
        RECT -49.465 -83.135 -49.295 -82.965 ;
        RECT -40.485 -83.135 -40.315 -82.965 ;
        RECT -40.015 -83.060 -39.845 -82.890 ;
        RECT -49.465 -83.595 -49.295 -83.425 ;
        RECT -40.485 -83.595 -40.315 -83.425 ;
        RECT -49.465 -84.055 -49.295 -83.885 ;
        RECT -40.485 -84.055 -40.315 -83.885 ;
        RECT -39.545 -83.135 -39.375 -82.965 ;
        RECT -30.565 -83.135 -30.395 -82.965 ;
        RECT -30.095 -83.060 -29.925 -82.890 ;
        RECT -39.545 -83.595 -39.375 -83.425 ;
        RECT -30.565 -83.595 -30.395 -83.425 ;
        RECT -39.545 -84.055 -39.375 -83.885 ;
        RECT -30.565 -84.055 -30.395 -83.885 ;
        RECT -29.625 -83.135 -29.455 -82.965 ;
        RECT -20.645 -83.135 -20.475 -82.965 ;
        RECT -20.175 -83.060 -20.005 -82.890 ;
        RECT -29.625 -83.595 -29.455 -83.425 ;
        RECT -20.645 -83.595 -20.475 -83.425 ;
        RECT -29.625 -84.055 -29.455 -83.885 ;
        RECT -20.645 -84.055 -20.475 -83.885 ;
        RECT -19.705 -83.135 -19.535 -82.965 ;
        RECT -10.725 -83.135 -10.555 -82.965 ;
        RECT -10.255 -83.060 -10.085 -82.890 ;
        RECT -19.705 -83.595 -19.535 -83.425 ;
        RECT -10.725 -83.595 -10.555 -83.425 ;
        RECT -19.705 -84.055 -19.535 -83.885 ;
        RECT -10.725 -84.055 -10.555 -83.885 ;
        RECT -9.785 -83.135 -9.615 -82.965 ;
        RECT -0.805 -83.135 -0.635 -82.965 ;
        RECT -0.335 -83.060 -0.165 -82.890 ;
        RECT -9.785 -83.595 -9.615 -83.425 ;
        RECT -0.805 -83.595 -0.635 -83.425 ;
        RECT -9.785 -84.055 -9.615 -83.885 ;
        RECT -0.805 -84.055 -0.635 -83.885 ;
        RECT 0.135 -83.135 0.305 -82.965 ;
        RECT 9.115 -83.135 9.285 -82.965 ;
        RECT 9.585 -83.060 9.755 -82.890 ;
        RECT 0.135 -83.595 0.305 -83.425 ;
        RECT 9.115 -83.595 9.285 -83.425 ;
        RECT 0.135 -84.055 0.305 -83.885 ;
        RECT 9.115 -84.055 9.285 -83.885 ;
        RECT 10.055 -83.135 10.225 -82.965 ;
        RECT 19.035 -83.135 19.205 -82.965 ;
        RECT 19.505 -83.060 19.675 -82.890 ;
        RECT 10.055 -83.595 10.225 -83.425 ;
        RECT 19.035 -83.595 19.205 -83.425 ;
        RECT 10.055 -84.055 10.225 -83.885 ;
        RECT 19.035 -84.055 19.205 -83.885 ;
        RECT 19.975 -83.135 20.145 -82.965 ;
        RECT 19.975 -83.595 20.145 -83.425 ;
        RECT 19.975 -84.055 20.145 -83.885 ;
        RECT -285.285 -172.755 -285.115 -172.585 ;
        RECT -284.815 -172.760 -284.645 -172.590 ;
        RECT -284.345 -172.755 -284.175 -172.585 ;
        RECT -285.285 -173.215 -285.115 -173.045 ;
        RECT -285.285 -173.675 -285.115 -173.505 ;
        RECT -275.365 -172.755 -275.195 -172.585 ;
        RECT -274.895 -172.760 -274.725 -172.590 ;
        RECT -274.425 -172.755 -274.255 -172.585 ;
        RECT -284.345 -173.215 -284.175 -173.045 ;
        RECT -275.365 -173.215 -275.195 -173.045 ;
        RECT -284.345 -173.675 -284.175 -173.505 ;
        RECT -275.365 -173.675 -275.195 -173.505 ;
        RECT -265.445 -172.755 -265.275 -172.585 ;
        RECT -264.975 -172.760 -264.805 -172.590 ;
        RECT -264.505 -172.755 -264.335 -172.585 ;
        RECT -274.425 -173.215 -274.255 -173.045 ;
        RECT -265.445 -173.215 -265.275 -173.045 ;
        RECT -274.425 -173.675 -274.255 -173.505 ;
        RECT -265.445 -173.675 -265.275 -173.505 ;
        RECT -255.525 -172.755 -255.355 -172.585 ;
        RECT -255.055 -172.760 -254.885 -172.590 ;
        RECT -254.585 -172.755 -254.415 -172.585 ;
        RECT -264.505 -173.215 -264.335 -173.045 ;
        RECT -255.525 -173.215 -255.355 -173.045 ;
        RECT -264.505 -173.675 -264.335 -173.505 ;
        RECT -255.525 -173.675 -255.355 -173.505 ;
        RECT -245.605 -172.755 -245.435 -172.585 ;
        RECT -245.135 -172.760 -244.965 -172.590 ;
        RECT -244.665 -172.755 -244.495 -172.585 ;
        RECT -254.585 -173.215 -254.415 -173.045 ;
        RECT -245.605 -173.215 -245.435 -173.045 ;
        RECT -254.585 -173.675 -254.415 -173.505 ;
        RECT -245.605 -173.675 -245.435 -173.505 ;
        RECT -235.685 -172.755 -235.515 -172.585 ;
        RECT -235.215 -172.760 -235.045 -172.590 ;
        RECT -234.745 -172.755 -234.575 -172.585 ;
        RECT -244.665 -173.215 -244.495 -173.045 ;
        RECT -235.685 -173.215 -235.515 -173.045 ;
        RECT -244.665 -173.675 -244.495 -173.505 ;
        RECT -235.685 -173.675 -235.515 -173.505 ;
        RECT -225.765 -172.755 -225.595 -172.585 ;
        RECT -225.295 -172.760 -225.125 -172.590 ;
        RECT -224.825 -172.755 -224.655 -172.585 ;
        RECT -234.745 -173.215 -234.575 -173.045 ;
        RECT -225.765 -173.215 -225.595 -173.045 ;
        RECT -234.745 -173.675 -234.575 -173.505 ;
        RECT -225.765 -173.675 -225.595 -173.505 ;
        RECT -215.845 -172.755 -215.675 -172.585 ;
        RECT -215.375 -172.760 -215.205 -172.590 ;
        RECT -214.905 -172.755 -214.735 -172.585 ;
        RECT -224.825 -173.215 -224.655 -173.045 ;
        RECT -215.845 -173.215 -215.675 -173.045 ;
        RECT -224.825 -173.675 -224.655 -173.505 ;
        RECT -215.845 -173.675 -215.675 -173.505 ;
        RECT -205.925 -172.755 -205.755 -172.585 ;
        RECT -205.455 -172.760 -205.285 -172.590 ;
        RECT -204.985 -172.755 -204.815 -172.585 ;
        RECT -214.905 -173.215 -214.735 -173.045 ;
        RECT -205.925 -173.215 -205.755 -173.045 ;
        RECT -214.905 -173.675 -214.735 -173.505 ;
        RECT -205.925 -173.675 -205.755 -173.505 ;
        RECT -196.005 -172.755 -195.835 -172.585 ;
        RECT -195.535 -172.760 -195.365 -172.590 ;
        RECT -195.065 -172.755 -194.895 -172.585 ;
        RECT -204.985 -173.215 -204.815 -173.045 ;
        RECT -196.005 -173.215 -195.835 -173.045 ;
        RECT -204.985 -173.675 -204.815 -173.505 ;
        RECT -196.005 -173.675 -195.835 -173.505 ;
        RECT -186.085 -172.755 -185.915 -172.585 ;
        RECT -185.615 -172.760 -185.445 -172.590 ;
        RECT -185.145 -172.755 -184.975 -172.585 ;
        RECT -195.065 -173.215 -194.895 -173.045 ;
        RECT -186.085 -173.215 -185.915 -173.045 ;
        RECT -195.065 -173.675 -194.895 -173.505 ;
        RECT -186.085 -173.675 -185.915 -173.505 ;
        RECT -176.165 -172.755 -175.995 -172.585 ;
        RECT -175.695 -172.760 -175.525 -172.590 ;
        RECT -175.225 -172.755 -175.055 -172.585 ;
        RECT -185.145 -173.215 -184.975 -173.045 ;
        RECT -176.165 -173.215 -175.995 -173.045 ;
        RECT -185.145 -173.675 -184.975 -173.505 ;
        RECT -176.165 -173.675 -175.995 -173.505 ;
        RECT -166.245 -172.755 -166.075 -172.585 ;
        RECT -165.775 -172.760 -165.605 -172.590 ;
        RECT -165.305 -172.755 -165.135 -172.585 ;
        RECT -175.225 -173.215 -175.055 -173.045 ;
        RECT -166.245 -173.215 -166.075 -173.045 ;
        RECT -175.225 -173.675 -175.055 -173.505 ;
        RECT -166.245 -173.675 -166.075 -173.505 ;
        RECT -156.325 -172.755 -156.155 -172.585 ;
        RECT -155.855 -172.760 -155.685 -172.590 ;
        RECT -155.385 -172.755 -155.215 -172.585 ;
        RECT -165.305 -173.215 -165.135 -173.045 ;
        RECT -156.325 -173.215 -156.155 -173.045 ;
        RECT -165.305 -173.675 -165.135 -173.505 ;
        RECT -156.325 -173.675 -156.155 -173.505 ;
        RECT -146.405 -172.755 -146.235 -172.585 ;
        RECT -145.935 -172.760 -145.765 -172.590 ;
        RECT -145.465 -172.755 -145.295 -172.585 ;
        RECT -155.385 -173.215 -155.215 -173.045 ;
        RECT -146.405 -173.215 -146.235 -173.045 ;
        RECT -155.385 -173.675 -155.215 -173.505 ;
        RECT -146.405 -173.675 -146.235 -173.505 ;
        RECT -136.485 -172.755 -136.315 -172.585 ;
        RECT -136.015 -172.760 -135.845 -172.590 ;
        RECT -135.545 -172.755 -135.375 -172.585 ;
        RECT -145.465 -173.215 -145.295 -173.045 ;
        RECT -136.485 -173.215 -136.315 -173.045 ;
        RECT -145.465 -173.675 -145.295 -173.505 ;
        RECT -136.485 -173.675 -136.315 -173.505 ;
        RECT -126.565 -172.755 -126.395 -172.585 ;
        RECT -126.095 -172.760 -125.925 -172.590 ;
        RECT -125.625 -172.755 -125.455 -172.585 ;
        RECT -135.545 -173.215 -135.375 -173.045 ;
        RECT -126.565 -173.215 -126.395 -173.045 ;
        RECT -135.545 -173.675 -135.375 -173.505 ;
        RECT -126.565 -173.675 -126.395 -173.505 ;
        RECT -116.645 -172.755 -116.475 -172.585 ;
        RECT -116.175 -172.760 -116.005 -172.590 ;
        RECT -115.705 -172.755 -115.535 -172.585 ;
        RECT -125.625 -173.215 -125.455 -173.045 ;
        RECT -116.645 -173.215 -116.475 -173.045 ;
        RECT -125.625 -173.675 -125.455 -173.505 ;
        RECT -116.645 -173.675 -116.475 -173.505 ;
        RECT -106.725 -172.755 -106.555 -172.585 ;
        RECT -106.255 -172.760 -106.085 -172.590 ;
        RECT -105.785 -172.755 -105.615 -172.585 ;
        RECT -115.705 -173.215 -115.535 -173.045 ;
        RECT -106.725 -173.215 -106.555 -173.045 ;
        RECT -115.705 -173.675 -115.535 -173.505 ;
        RECT -106.725 -173.675 -106.555 -173.505 ;
        RECT -96.805 -172.755 -96.635 -172.585 ;
        RECT -96.335 -172.760 -96.165 -172.590 ;
        RECT -95.865 -172.755 -95.695 -172.585 ;
        RECT -105.785 -173.215 -105.615 -173.045 ;
        RECT -96.805 -173.215 -96.635 -173.045 ;
        RECT -105.785 -173.675 -105.615 -173.505 ;
        RECT -96.805 -173.675 -96.635 -173.505 ;
        RECT -86.885 -172.755 -86.715 -172.585 ;
        RECT -86.415 -172.760 -86.245 -172.590 ;
        RECT -85.945 -172.755 -85.775 -172.585 ;
        RECT -95.865 -173.215 -95.695 -173.045 ;
        RECT -86.885 -173.215 -86.715 -173.045 ;
        RECT -95.865 -173.675 -95.695 -173.505 ;
        RECT -86.885 -173.675 -86.715 -173.505 ;
        RECT -76.965 -172.755 -76.795 -172.585 ;
        RECT -76.495 -172.760 -76.325 -172.590 ;
        RECT -76.025 -172.755 -75.855 -172.585 ;
        RECT -85.945 -173.215 -85.775 -173.045 ;
        RECT -76.965 -173.215 -76.795 -173.045 ;
        RECT -85.945 -173.675 -85.775 -173.505 ;
        RECT -76.965 -173.675 -76.795 -173.505 ;
        RECT -67.045 -172.755 -66.875 -172.585 ;
        RECT -66.575 -172.760 -66.405 -172.590 ;
        RECT -66.105 -172.755 -65.935 -172.585 ;
        RECT -76.025 -173.215 -75.855 -173.045 ;
        RECT -67.045 -173.215 -66.875 -173.045 ;
        RECT -76.025 -173.675 -75.855 -173.505 ;
        RECT -67.045 -173.675 -66.875 -173.505 ;
        RECT -57.125 -172.755 -56.955 -172.585 ;
        RECT -56.655 -172.760 -56.485 -172.590 ;
        RECT -56.185 -172.755 -56.015 -172.585 ;
        RECT -66.105 -173.215 -65.935 -173.045 ;
        RECT -57.125 -173.215 -56.955 -173.045 ;
        RECT -66.105 -173.675 -65.935 -173.505 ;
        RECT -57.125 -173.675 -56.955 -173.505 ;
        RECT -47.205 -172.755 -47.035 -172.585 ;
        RECT -46.735 -172.760 -46.565 -172.590 ;
        RECT -46.265 -172.755 -46.095 -172.585 ;
        RECT -56.185 -173.215 -56.015 -173.045 ;
        RECT -47.205 -173.215 -47.035 -173.045 ;
        RECT -56.185 -173.675 -56.015 -173.505 ;
        RECT -47.205 -173.675 -47.035 -173.505 ;
        RECT -37.285 -172.755 -37.115 -172.585 ;
        RECT -36.815 -172.760 -36.645 -172.590 ;
        RECT -36.345 -172.755 -36.175 -172.585 ;
        RECT -46.265 -173.215 -46.095 -173.045 ;
        RECT -37.285 -173.215 -37.115 -173.045 ;
        RECT -46.265 -173.675 -46.095 -173.505 ;
        RECT -37.285 -173.675 -37.115 -173.505 ;
        RECT -27.365 -172.755 -27.195 -172.585 ;
        RECT -26.895 -172.760 -26.725 -172.590 ;
        RECT -26.425 -172.755 -26.255 -172.585 ;
        RECT -36.345 -173.215 -36.175 -173.045 ;
        RECT -27.365 -173.215 -27.195 -173.045 ;
        RECT -36.345 -173.675 -36.175 -173.505 ;
        RECT -27.365 -173.675 -27.195 -173.505 ;
        RECT -17.445 -172.755 -17.275 -172.585 ;
        RECT -16.975 -172.760 -16.805 -172.590 ;
        RECT -16.505 -172.755 -16.335 -172.585 ;
        RECT -26.425 -173.215 -26.255 -173.045 ;
        RECT -17.445 -173.215 -17.275 -173.045 ;
        RECT -26.425 -173.675 -26.255 -173.505 ;
        RECT -17.445 -173.675 -17.275 -173.505 ;
        RECT -7.525 -172.755 -7.355 -172.585 ;
        RECT -7.055 -172.760 -6.885 -172.590 ;
        RECT -6.585 -172.755 -6.415 -172.585 ;
        RECT -16.505 -173.215 -16.335 -173.045 ;
        RECT -7.525 -173.215 -7.355 -173.045 ;
        RECT -16.505 -173.675 -16.335 -173.505 ;
        RECT -7.525 -173.675 -7.355 -173.505 ;
        RECT 2.395 -172.755 2.565 -172.585 ;
        RECT 2.865 -172.760 3.035 -172.590 ;
        RECT 3.335 -172.755 3.505 -172.585 ;
        RECT -6.585 -173.215 -6.415 -173.045 ;
        RECT 2.395 -173.215 2.565 -173.045 ;
        RECT -6.585 -173.675 -6.415 -173.505 ;
        RECT 2.395 -173.675 2.565 -173.505 ;
        RECT 12.315 -172.755 12.485 -172.585 ;
        RECT 12.785 -172.760 12.955 -172.590 ;
        RECT 13.255 -172.755 13.425 -172.585 ;
        RECT 3.335 -173.215 3.505 -173.045 ;
        RECT 12.315 -173.215 12.485 -173.045 ;
        RECT 3.335 -173.675 3.505 -173.505 ;
        RECT 12.315 -173.675 12.485 -173.505 ;
        RECT 22.235 -172.755 22.405 -172.585 ;
        RECT 22.705 -172.760 22.875 -172.590 ;
        RECT 13.255 -173.215 13.425 -173.045 ;
        RECT 22.235 -173.215 22.405 -173.045 ;
        RECT 13.255 -173.675 13.425 -173.505 ;
        RECT 22.235 -173.675 22.405 -173.505 ;
        RECT -291.155 -174.335 -290.985 -174.165 ;
        RECT -290.695 -174.335 -290.525 -174.165 ;
        RECT -290.235 -174.335 -290.065 -174.165 ;
        RECT -289.775 -174.335 -289.605 -174.165 ;
        RECT -289.315 -174.335 -289.145 -174.165 ;
        RECT -288.855 -174.335 -288.685 -174.165 ;
        RECT -288.395 -174.335 -288.225 -174.165 ;
        RECT -281.235 -174.335 -281.065 -174.165 ;
        RECT -280.775 -174.335 -280.605 -174.165 ;
        RECT -280.315 -174.335 -280.145 -174.165 ;
        RECT -279.855 -174.335 -279.685 -174.165 ;
        RECT -279.395 -174.335 -279.225 -174.165 ;
        RECT -278.935 -174.335 -278.765 -174.165 ;
        RECT -278.475 -174.335 -278.305 -174.165 ;
        RECT -271.315 -174.335 -271.145 -174.165 ;
        RECT -270.855 -174.335 -270.685 -174.165 ;
        RECT -270.395 -174.335 -270.225 -174.165 ;
        RECT -269.935 -174.335 -269.765 -174.165 ;
        RECT -269.475 -174.335 -269.305 -174.165 ;
        RECT -269.015 -174.335 -268.845 -174.165 ;
        RECT -268.555 -174.335 -268.385 -174.165 ;
        RECT -261.395 -174.335 -261.225 -174.165 ;
        RECT -260.935 -174.335 -260.765 -174.165 ;
        RECT -260.475 -174.335 -260.305 -174.165 ;
        RECT -260.015 -174.335 -259.845 -174.165 ;
        RECT -259.555 -174.335 -259.385 -174.165 ;
        RECT -259.095 -174.335 -258.925 -174.165 ;
        RECT -258.635 -174.335 -258.465 -174.165 ;
        RECT -251.475 -174.335 -251.305 -174.165 ;
        RECT -251.015 -174.335 -250.845 -174.165 ;
        RECT -250.555 -174.335 -250.385 -174.165 ;
        RECT -250.095 -174.335 -249.925 -174.165 ;
        RECT -249.635 -174.335 -249.465 -174.165 ;
        RECT -249.175 -174.335 -249.005 -174.165 ;
        RECT -248.715 -174.335 -248.545 -174.165 ;
        RECT -241.555 -174.335 -241.385 -174.165 ;
        RECT -241.095 -174.335 -240.925 -174.165 ;
        RECT -240.635 -174.335 -240.465 -174.165 ;
        RECT -240.175 -174.335 -240.005 -174.165 ;
        RECT -239.715 -174.335 -239.545 -174.165 ;
        RECT -239.255 -174.335 -239.085 -174.165 ;
        RECT -238.795 -174.335 -238.625 -174.165 ;
        RECT -231.635 -174.335 -231.465 -174.165 ;
        RECT -231.175 -174.335 -231.005 -174.165 ;
        RECT -230.715 -174.335 -230.545 -174.165 ;
        RECT -230.255 -174.335 -230.085 -174.165 ;
        RECT -229.795 -174.335 -229.625 -174.165 ;
        RECT -229.335 -174.335 -229.165 -174.165 ;
        RECT -228.875 -174.335 -228.705 -174.165 ;
        RECT -221.715 -174.335 -221.545 -174.165 ;
        RECT -221.255 -174.335 -221.085 -174.165 ;
        RECT -220.795 -174.335 -220.625 -174.165 ;
        RECT -220.335 -174.335 -220.165 -174.165 ;
        RECT -219.875 -174.335 -219.705 -174.165 ;
        RECT -219.415 -174.335 -219.245 -174.165 ;
        RECT -218.955 -174.335 -218.785 -174.165 ;
        RECT -211.795 -174.335 -211.625 -174.165 ;
        RECT -211.335 -174.335 -211.165 -174.165 ;
        RECT -210.875 -174.335 -210.705 -174.165 ;
        RECT -210.415 -174.335 -210.245 -174.165 ;
        RECT -209.955 -174.335 -209.785 -174.165 ;
        RECT -209.495 -174.335 -209.325 -174.165 ;
        RECT -209.035 -174.335 -208.865 -174.165 ;
        RECT -201.875 -174.335 -201.705 -174.165 ;
        RECT -201.415 -174.335 -201.245 -174.165 ;
        RECT -200.955 -174.335 -200.785 -174.165 ;
        RECT -200.495 -174.335 -200.325 -174.165 ;
        RECT -200.035 -174.335 -199.865 -174.165 ;
        RECT -199.575 -174.335 -199.405 -174.165 ;
        RECT -199.115 -174.335 -198.945 -174.165 ;
        RECT -191.955 -174.335 -191.785 -174.165 ;
        RECT -191.495 -174.335 -191.325 -174.165 ;
        RECT -191.035 -174.335 -190.865 -174.165 ;
        RECT -190.575 -174.335 -190.405 -174.165 ;
        RECT -190.115 -174.335 -189.945 -174.165 ;
        RECT -189.655 -174.335 -189.485 -174.165 ;
        RECT -189.195 -174.335 -189.025 -174.165 ;
        RECT -182.035 -174.335 -181.865 -174.165 ;
        RECT -181.575 -174.335 -181.405 -174.165 ;
        RECT -181.115 -174.335 -180.945 -174.165 ;
        RECT -180.655 -174.335 -180.485 -174.165 ;
        RECT -180.195 -174.335 -180.025 -174.165 ;
        RECT -179.735 -174.335 -179.565 -174.165 ;
        RECT -179.275 -174.335 -179.105 -174.165 ;
        RECT -172.115 -174.335 -171.945 -174.165 ;
        RECT -171.655 -174.335 -171.485 -174.165 ;
        RECT -171.195 -174.335 -171.025 -174.165 ;
        RECT -170.735 -174.335 -170.565 -174.165 ;
        RECT -170.275 -174.335 -170.105 -174.165 ;
        RECT -169.815 -174.335 -169.645 -174.165 ;
        RECT -169.355 -174.335 -169.185 -174.165 ;
        RECT -162.195 -174.335 -162.025 -174.165 ;
        RECT -161.735 -174.335 -161.565 -174.165 ;
        RECT -161.275 -174.335 -161.105 -174.165 ;
        RECT -160.815 -174.335 -160.645 -174.165 ;
        RECT -160.355 -174.335 -160.185 -174.165 ;
        RECT -159.895 -174.335 -159.725 -174.165 ;
        RECT -159.435 -174.335 -159.265 -174.165 ;
        RECT -152.275 -174.335 -152.105 -174.165 ;
        RECT -151.815 -174.335 -151.645 -174.165 ;
        RECT -151.355 -174.335 -151.185 -174.165 ;
        RECT -150.895 -174.335 -150.725 -174.165 ;
        RECT -150.435 -174.335 -150.265 -174.165 ;
        RECT -149.975 -174.335 -149.805 -174.165 ;
        RECT -149.515 -174.335 -149.345 -174.165 ;
        RECT -142.355 -174.335 -142.185 -174.165 ;
        RECT -141.895 -174.335 -141.725 -174.165 ;
        RECT -141.435 -174.335 -141.265 -174.165 ;
        RECT -140.975 -174.335 -140.805 -174.165 ;
        RECT -140.515 -174.335 -140.345 -174.165 ;
        RECT -140.055 -174.335 -139.885 -174.165 ;
        RECT -139.595 -174.335 -139.425 -174.165 ;
        RECT -132.435 -174.335 -132.265 -174.165 ;
        RECT -131.975 -174.335 -131.805 -174.165 ;
        RECT -131.515 -174.335 -131.345 -174.165 ;
        RECT -131.055 -174.335 -130.885 -174.165 ;
        RECT -130.595 -174.335 -130.425 -174.165 ;
        RECT -130.135 -174.335 -129.965 -174.165 ;
        RECT -129.675 -174.335 -129.505 -174.165 ;
        RECT -122.515 -174.335 -122.345 -174.165 ;
        RECT -122.055 -174.335 -121.885 -174.165 ;
        RECT -121.595 -174.335 -121.425 -174.165 ;
        RECT -121.135 -174.335 -120.965 -174.165 ;
        RECT -120.675 -174.335 -120.505 -174.165 ;
        RECT -120.215 -174.335 -120.045 -174.165 ;
        RECT -119.755 -174.335 -119.585 -174.165 ;
        RECT -112.595 -174.335 -112.425 -174.165 ;
        RECT -112.135 -174.335 -111.965 -174.165 ;
        RECT -111.675 -174.335 -111.505 -174.165 ;
        RECT -111.215 -174.335 -111.045 -174.165 ;
        RECT -110.755 -174.335 -110.585 -174.165 ;
        RECT -110.295 -174.335 -110.125 -174.165 ;
        RECT -109.835 -174.335 -109.665 -174.165 ;
        RECT -102.675 -174.335 -102.505 -174.165 ;
        RECT -102.215 -174.335 -102.045 -174.165 ;
        RECT -101.755 -174.335 -101.585 -174.165 ;
        RECT -101.295 -174.335 -101.125 -174.165 ;
        RECT -100.835 -174.335 -100.665 -174.165 ;
        RECT -100.375 -174.335 -100.205 -174.165 ;
        RECT -99.915 -174.335 -99.745 -174.165 ;
        RECT -92.755 -174.335 -92.585 -174.165 ;
        RECT -92.295 -174.335 -92.125 -174.165 ;
        RECT -91.835 -174.335 -91.665 -174.165 ;
        RECT -91.375 -174.335 -91.205 -174.165 ;
        RECT -90.915 -174.335 -90.745 -174.165 ;
        RECT -90.455 -174.335 -90.285 -174.165 ;
        RECT -89.995 -174.335 -89.825 -174.165 ;
        RECT -82.835 -174.335 -82.665 -174.165 ;
        RECT -82.375 -174.335 -82.205 -174.165 ;
        RECT -81.915 -174.335 -81.745 -174.165 ;
        RECT -81.455 -174.335 -81.285 -174.165 ;
        RECT -80.995 -174.335 -80.825 -174.165 ;
        RECT -80.535 -174.335 -80.365 -174.165 ;
        RECT -80.075 -174.335 -79.905 -174.165 ;
        RECT -72.915 -174.335 -72.745 -174.165 ;
        RECT -72.455 -174.335 -72.285 -174.165 ;
        RECT -71.995 -174.335 -71.825 -174.165 ;
        RECT -71.535 -174.335 -71.365 -174.165 ;
        RECT -71.075 -174.335 -70.905 -174.165 ;
        RECT -70.615 -174.335 -70.445 -174.165 ;
        RECT -70.155 -174.335 -69.985 -174.165 ;
        RECT -62.995 -174.335 -62.825 -174.165 ;
        RECT -62.535 -174.335 -62.365 -174.165 ;
        RECT -62.075 -174.335 -61.905 -174.165 ;
        RECT -61.615 -174.335 -61.445 -174.165 ;
        RECT -61.155 -174.335 -60.985 -174.165 ;
        RECT -60.695 -174.335 -60.525 -174.165 ;
        RECT -60.235 -174.335 -60.065 -174.165 ;
        RECT -53.075 -174.335 -52.905 -174.165 ;
        RECT -52.615 -174.335 -52.445 -174.165 ;
        RECT -52.155 -174.335 -51.985 -174.165 ;
        RECT -51.695 -174.335 -51.525 -174.165 ;
        RECT -51.235 -174.335 -51.065 -174.165 ;
        RECT -50.775 -174.335 -50.605 -174.165 ;
        RECT -50.315 -174.335 -50.145 -174.165 ;
        RECT -43.155 -174.335 -42.985 -174.165 ;
        RECT -42.695 -174.335 -42.525 -174.165 ;
        RECT -42.235 -174.335 -42.065 -174.165 ;
        RECT -41.775 -174.335 -41.605 -174.165 ;
        RECT -41.315 -174.335 -41.145 -174.165 ;
        RECT -40.855 -174.335 -40.685 -174.165 ;
        RECT -40.395 -174.335 -40.225 -174.165 ;
        RECT -33.235 -174.335 -33.065 -174.165 ;
        RECT -32.775 -174.335 -32.605 -174.165 ;
        RECT -32.315 -174.335 -32.145 -174.165 ;
        RECT -31.855 -174.335 -31.685 -174.165 ;
        RECT -31.395 -174.335 -31.225 -174.165 ;
        RECT -30.935 -174.335 -30.765 -174.165 ;
        RECT -30.475 -174.335 -30.305 -174.165 ;
        RECT -23.315 -174.335 -23.145 -174.165 ;
        RECT -22.855 -174.335 -22.685 -174.165 ;
        RECT -22.395 -174.335 -22.225 -174.165 ;
        RECT -21.935 -174.335 -21.765 -174.165 ;
        RECT -21.475 -174.335 -21.305 -174.165 ;
        RECT -21.015 -174.335 -20.845 -174.165 ;
        RECT -20.555 -174.335 -20.385 -174.165 ;
        RECT -13.395 -174.335 -13.225 -174.165 ;
        RECT -12.935 -174.335 -12.765 -174.165 ;
        RECT -12.475 -174.335 -12.305 -174.165 ;
        RECT -12.015 -174.335 -11.845 -174.165 ;
        RECT -11.555 -174.335 -11.385 -174.165 ;
        RECT -11.095 -174.335 -10.925 -174.165 ;
        RECT -10.635 -174.335 -10.465 -174.165 ;
        RECT -3.475 -174.335 -3.305 -174.165 ;
        RECT -3.015 -174.335 -2.845 -174.165 ;
        RECT -2.555 -174.335 -2.385 -174.165 ;
        RECT -2.095 -174.335 -1.925 -174.165 ;
        RECT -1.635 -174.335 -1.465 -174.165 ;
        RECT -1.175 -174.335 -1.005 -174.165 ;
        RECT -0.715 -174.335 -0.545 -174.165 ;
        RECT 6.445 -174.335 6.615 -174.165 ;
        RECT 6.905 -174.335 7.075 -174.165 ;
        RECT 7.365 -174.335 7.535 -174.165 ;
        RECT 7.825 -174.335 7.995 -174.165 ;
        RECT 8.285 -174.335 8.455 -174.165 ;
        RECT 8.745 -174.335 8.915 -174.165 ;
        RECT 9.205 -174.335 9.375 -174.165 ;
        RECT 16.365 -174.335 16.535 -174.165 ;
        RECT 16.825 -174.335 16.995 -174.165 ;
        RECT 17.285 -174.335 17.455 -174.165 ;
        RECT 17.745 -174.335 17.915 -174.165 ;
        RECT 18.205 -174.335 18.375 -174.165 ;
        RECT 18.665 -174.335 18.835 -174.165 ;
        RECT 19.125 -174.335 19.295 -174.165 ;
        RECT -286.195 -177.055 -286.025 -176.885 ;
        RECT -285.735 -177.055 -285.565 -176.885 ;
        RECT -285.275 -177.055 -285.105 -176.885 ;
        RECT -284.815 -177.055 -284.645 -176.885 ;
        RECT -284.355 -177.055 -284.185 -176.885 ;
        RECT -283.895 -177.055 -283.725 -176.885 ;
        RECT -283.435 -177.055 -283.265 -176.885 ;
        RECT -276.275 -177.055 -276.105 -176.885 ;
        RECT -275.815 -177.055 -275.645 -176.885 ;
        RECT -275.355 -177.055 -275.185 -176.885 ;
        RECT -274.895 -177.055 -274.725 -176.885 ;
        RECT -274.435 -177.055 -274.265 -176.885 ;
        RECT -273.975 -177.055 -273.805 -176.885 ;
        RECT -273.515 -177.055 -273.345 -176.885 ;
        RECT -266.355 -177.055 -266.185 -176.885 ;
        RECT -265.895 -177.055 -265.725 -176.885 ;
        RECT -265.435 -177.055 -265.265 -176.885 ;
        RECT -264.975 -177.055 -264.805 -176.885 ;
        RECT -264.515 -177.055 -264.345 -176.885 ;
        RECT -264.055 -177.055 -263.885 -176.885 ;
        RECT -263.595 -177.055 -263.425 -176.885 ;
        RECT -256.435 -177.055 -256.265 -176.885 ;
        RECT -255.975 -177.055 -255.805 -176.885 ;
        RECT -255.515 -177.055 -255.345 -176.885 ;
        RECT -255.055 -177.055 -254.885 -176.885 ;
        RECT -254.595 -177.055 -254.425 -176.885 ;
        RECT -254.135 -177.055 -253.965 -176.885 ;
        RECT -253.675 -177.055 -253.505 -176.885 ;
        RECT -246.515 -177.055 -246.345 -176.885 ;
        RECT -246.055 -177.055 -245.885 -176.885 ;
        RECT -245.595 -177.055 -245.425 -176.885 ;
        RECT -245.135 -177.055 -244.965 -176.885 ;
        RECT -244.675 -177.055 -244.505 -176.885 ;
        RECT -244.215 -177.055 -244.045 -176.885 ;
        RECT -243.755 -177.055 -243.585 -176.885 ;
        RECT -236.595 -177.055 -236.425 -176.885 ;
        RECT -236.135 -177.055 -235.965 -176.885 ;
        RECT -235.675 -177.055 -235.505 -176.885 ;
        RECT -235.215 -177.055 -235.045 -176.885 ;
        RECT -234.755 -177.055 -234.585 -176.885 ;
        RECT -234.295 -177.055 -234.125 -176.885 ;
        RECT -233.835 -177.055 -233.665 -176.885 ;
        RECT -226.675 -177.055 -226.505 -176.885 ;
        RECT -226.215 -177.055 -226.045 -176.885 ;
        RECT -225.755 -177.055 -225.585 -176.885 ;
        RECT -225.295 -177.055 -225.125 -176.885 ;
        RECT -224.835 -177.055 -224.665 -176.885 ;
        RECT -224.375 -177.055 -224.205 -176.885 ;
        RECT -223.915 -177.055 -223.745 -176.885 ;
        RECT -216.755 -177.055 -216.585 -176.885 ;
        RECT -216.295 -177.055 -216.125 -176.885 ;
        RECT -215.835 -177.055 -215.665 -176.885 ;
        RECT -215.375 -177.055 -215.205 -176.885 ;
        RECT -214.915 -177.055 -214.745 -176.885 ;
        RECT -214.455 -177.055 -214.285 -176.885 ;
        RECT -213.995 -177.055 -213.825 -176.885 ;
        RECT -206.835 -177.055 -206.665 -176.885 ;
        RECT -206.375 -177.055 -206.205 -176.885 ;
        RECT -205.915 -177.055 -205.745 -176.885 ;
        RECT -205.455 -177.055 -205.285 -176.885 ;
        RECT -204.995 -177.055 -204.825 -176.885 ;
        RECT -204.535 -177.055 -204.365 -176.885 ;
        RECT -204.075 -177.055 -203.905 -176.885 ;
        RECT -196.915 -177.055 -196.745 -176.885 ;
        RECT -196.455 -177.055 -196.285 -176.885 ;
        RECT -195.995 -177.055 -195.825 -176.885 ;
        RECT -195.535 -177.055 -195.365 -176.885 ;
        RECT -195.075 -177.055 -194.905 -176.885 ;
        RECT -194.615 -177.055 -194.445 -176.885 ;
        RECT -194.155 -177.055 -193.985 -176.885 ;
        RECT -186.995 -177.055 -186.825 -176.885 ;
        RECT -186.535 -177.055 -186.365 -176.885 ;
        RECT -186.075 -177.055 -185.905 -176.885 ;
        RECT -185.615 -177.055 -185.445 -176.885 ;
        RECT -185.155 -177.055 -184.985 -176.885 ;
        RECT -184.695 -177.055 -184.525 -176.885 ;
        RECT -184.235 -177.055 -184.065 -176.885 ;
        RECT -177.075 -177.055 -176.905 -176.885 ;
        RECT -176.615 -177.055 -176.445 -176.885 ;
        RECT -176.155 -177.055 -175.985 -176.885 ;
        RECT -175.695 -177.055 -175.525 -176.885 ;
        RECT -175.235 -177.055 -175.065 -176.885 ;
        RECT -174.775 -177.055 -174.605 -176.885 ;
        RECT -174.315 -177.055 -174.145 -176.885 ;
        RECT -167.155 -177.055 -166.985 -176.885 ;
        RECT -166.695 -177.055 -166.525 -176.885 ;
        RECT -166.235 -177.055 -166.065 -176.885 ;
        RECT -165.775 -177.055 -165.605 -176.885 ;
        RECT -165.315 -177.055 -165.145 -176.885 ;
        RECT -164.855 -177.055 -164.685 -176.885 ;
        RECT -164.395 -177.055 -164.225 -176.885 ;
        RECT -157.235 -177.055 -157.065 -176.885 ;
        RECT -156.775 -177.055 -156.605 -176.885 ;
        RECT -156.315 -177.055 -156.145 -176.885 ;
        RECT -155.855 -177.055 -155.685 -176.885 ;
        RECT -155.395 -177.055 -155.225 -176.885 ;
        RECT -154.935 -177.055 -154.765 -176.885 ;
        RECT -154.475 -177.055 -154.305 -176.885 ;
        RECT -147.315 -177.055 -147.145 -176.885 ;
        RECT -146.855 -177.055 -146.685 -176.885 ;
        RECT -146.395 -177.055 -146.225 -176.885 ;
        RECT -145.935 -177.055 -145.765 -176.885 ;
        RECT -145.475 -177.055 -145.305 -176.885 ;
        RECT -145.015 -177.055 -144.845 -176.885 ;
        RECT -144.555 -177.055 -144.385 -176.885 ;
        RECT -137.395 -177.055 -137.225 -176.885 ;
        RECT -136.935 -177.055 -136.765 -176.885 ;
        RECT -136.475 -177.055 -136.305 -176.885 ;
        RECT -136.015 -177.055 -135.845 -176.885 ;
        RECT -135.555 -177.055 -135.385 -176.885 ;
        RECT -135.095 -177.055 -134.925 -176.885 ;
        RECT -134.635 -177.055 -134.465 -176.885 ;
        RECT -127.475 -177.055 -127.305 -176.885 ;
        RECT -127.015 -177.055 -126.845 -176.885 ;
        RECT -126.555 -177.055 -126.385 -176.885 ;
        RECT -126.095 -177.055 -125.925 -176.885 ;
        RECT -125.635 -177.055 -125.465 -176.885 ;
        RECT -125.175 -177.055 -125.005 -176.885 ;
        RECT -124.715 -177.055 -124.545 -176.885 ;
        RECT -117.555 -177.055 -117.385 -176.885 ;
        RECT -117.095 -177.055 -116.925 -176.885 ;
        RECT -116.635 -177.055 -116.465 -176.885 ;
        RECT -116.175 -177.055 -116.005 -176.885 ;
        RECT -115.715 -177.055 -115.545 -176.885 ;
        RECT -115.255 -177.055 -115.085 -176.885 ;
        RECT -114.795 -177.055 -114.625 -176.885 ;
        RECT -107.635 -177.055 -107.465 -176.885 ;
        RECT -107.175 -177.055 -107.005 -176.885 ;
        RECT -106.715 -177.055 -106.545 -176.885 ;
        RECT -106.255 -177.055 -106.085 -176.885 ;
        RECT -105.795 -177.055 -105.625 -176.885 ;
        RECT -105.335 -177.055 -105.165 -176.885 ;
        RECT -104.875 -177.055 -104.705 -176.885 ;
        RECT -97.715 -177.055 -97.545 -176.885 ;
        RECT -97.255 -177.055 -97.085 -176.885 ;
        RECT -96.795 -177.055 -96.625 -176.885 ;
        RECT -96.335 -177.055 -96.165 -176.885 ;
        RECT -95.875 -177.055 -95.705 -176.885 ;
        RECT -95.415 -177.055 -95.245 -176.885 ;
        RECT -94.955 -177.055 -94.785 -176.885 ;
        RECT -87.795 -177.055 -87.625 -176.885 ;
        RECT -87.335 -177.055 -87.165 -176.885 ;
        RECT -86.875 -177.055 -86.705 -176.885 ;
        RECT -86.415 -177.055 -86.245 -176.885 ;
        RECT -85.955 -177.055 -85.785 -176.885 ;
        RECT -85.495 -177.055 -85.325 -176.885 ;
        RECT -85.035 -177.055 -84.865 -176.885 ;
        RECT -77.875 -177.055 -77.705 -176.885 ;
        RECT -77.415 -177.055 -77.245 -176.885 ;
        RECT -76.955 -177.055 -76.785 -176.885 ;
        RECT -76.495 -177.055 -76.325 -176.885 ;
        RECT -76.035 -177.055 -75.865 -176.885 ;
        RECT -75.575 -177.055 -75.405 -176.885 ;
        RECT -75.115 -177.055 -74.945 -176.885 ;
        RECT -67.955 -177.055 -67.785 -176.885 ;
        RECT -67.495 -177.055 -67.325 -176.885 ;
        RECT -67.035 -177.055 -66.865 -176.885 ;
        RECT -66.575 -177.055 -66.405 -176.885 ;
        RECT -66.115 -177.055 -65.945 -176.885 ;
        RECT -65.655 -177.055 -65.485 -176.885 ;
        RECT -65.195 -177.055 -65.025 -176.885 ;
        RECT -58.035 -177.055 -57.865 -176.885 ;
        RECT -57.575 -177.055 -57.405 -176.885 ;
        RECT -57.115 -177.055 -56.945 -176.885 ;
        RECT -56.655 -177.055 -56.485 -176.885 ;
        RECT -56.195 -177.055 -56.025 -176.885 ;
        RECT -55.735 -177.055 -55.565 -176.885 ;
        RECT -55.275 -177.055 -55.105 -176.885 ;
        RECT -48.115 -177.055 -47.945 -176.885 ;
        RECT -47.655 -177.055 -47.485 -176.885 ;
        RECT -47.195 -177.055 -47.025 -176.885 ;
        RECT -46.735 -177.055 -46.565 -176.885 ;
        RECT -46.275 -177.055 -46.105 -176.885 ;
        RECT -45.815 -177.055 -45.645 -176.885 ;
        RECT -45.355 -177.055 -45.185 -176.885 ;
        RECT -38.195 -177.055 -38.025 -176.885 ;
        RECT -37.735 -177.055 -37.565 -176.885 ;
        RECT -37.275 -177.055 -37.105 -176.885 ;
        RECT -36.815 -177.055 -36.645 -176.885 ;
        RECT -36.355 -177.055 -36.185 -176.885 ;
        RECT -35.895 -177.055 -35.725 -176.885 ;
        RECT -35.435 -177.055 -35.265 -176.885 ;
        RECT -28.275 -177.055 -28.105 -176.885 ;
        RECT -27.815 -177.055 -27.645 -176.885 ;
        RECT -27.355 -177.055 -27.185 -176.885 ;
        RECT -26.895 -177.055 -26.725 -176.885 ;
        RECT -26.435 -177.055 -26.265 -176.885 ;
        RECT -25.975 -177.055 -25.805 -176.885 ;
        RECT -25.515 -177.055 -25.345 -176.885 ;
        RECT -18.355 -177.055 -18.185 -176.885 ;
        RECT -17.895 -177.055 -17.725 -176.885 ;
        RECT -17.435 -177.055 -17.265 -176.885 ;
        RECT -16.975 -177.055 -16.805 -176.885 ;
        RECT -16.515 -177.055 -16.345 -176.885 ;
        RECT -16.055 -177.055 -15.885 -176.885 ;
        RECT -15.595 -177.055 -15.425 -176.885 ;
        RECT -8.435 -177.055 -8.265 -176.885 ;
        RECT -7.975 -177.055 -7.805 -176.885 ;
        RECT -7.515 -177.055 -7.345 -176.885 ;
        RECT -7.055 -177.055 -6.885 -176.885 ;
        RECT -6.595 -177.055 -6.425 -176.885 ;
        RECT -6.135 -177.055 -5.965 -176.885 ;
        RECT -5.675 -177.055 -5.505 -176.885 ;
        RECT 1.485 -177.055 1.655 -176.885 ;
        RECT 1.945 -177.055 2.115 -176.885 ;
        RECT 2.405 -177.055 2.575 -176.885 ;
        RECT 2.865 -177.055 3.035 -176.885 ;
        RECT 3.325 -177.055 3.495 -176.885 ;
        RECT 3.785 -177.055 3.955 -176.885 ;
        RECT 4.245 -177.055 4.415 -176.885 ;
        RECT 11.405 -177.055 11.575 -176.885 ;
        RECT 11.865 -177.055 12.035 -176.885 ;
        RECT 12.325 -177.055 12.495 -176.885 ;
        RECT 12.785 -177.055 12.955 -176.885 ;
        RECT 13.245 -177.055 13.415 -176.885 ;
        RECT 13.705 -177.055 13.875 -176.885 ;
        RECT 14.165 -177.055 14.335 -176.885 ;
        RECT 21.325 -177.055 21.495 -176.885 ;
        RECT 21.785 -177.055 21.955 -176.885 ;
        RECT 22.245 -177.055 22.415 -176.885 ;
        RECT 22.705 -177.055 22.875 -176.885 ;
        RECT -290.245 -177.715 -290.075 -177.545 ;
        RECT -289.775 -177.640 -289.605 -177.470 ;
        RECT -290.245 -178.175 -290.075 -178.005 ;
        RECT -290.245 -178.635 -290.075 -178.465 ;
        RECT -289.305 -177.715 -289.135 -177.545 ;
        RECT -280.325 -177.715 -280.155 -177.545 ;
        RECT -279.855 -177.640 -279.685 -177.470 ;
        RECT -289.305 -178.175 -289.135 -178.005 ;
        RECT -280.325 -178.175 -280.155 -178.005 ;
        RECT -289.305 -178.635 -289.135 -178.465 ;
        RECT -280.325 -178.635 -280.155 -178.465 ;
        RECT -279.385 -177.715 -279.215 -177.545 ;
        RECT -270.405 -177.715 -270.235 -177.545 ;
        RECT -269.935 -177.640 -269.765 -177.470 ;
        RECT -279.385 -178.175 -279.215 -178.005 ;
        RECT -270.405 -178.175 -270.235 -178.005 ;
        RECT -279.385 -178.635 -279.215 -178.465 ;
        RECT -270.405 -178.635 -270.235 -178.465 ;
        RECT -269.465 -177.715 -269.295 -177.545 ;
        RECT -260.485 -177.715 -260.315 -177.545 ;
        RECT -260.015 -177.640 -259.845 -177.470 ;
        RECT -269.465 -178.175 -269.295 -178.005 ;
        RECT -260.485 -178.175 -260.315 -178.005 ;
        RECT -269.465 -178.635 -269.295 -178.465 ;
        RECT -260.485 -178.635 -260.315 -178.465 ;
        RECT -259.545 -177.715 -259.375 -177.545 ;
        RECT -250.565 -177.715 -250.395 -177.545 ;
        RECT -250.095 -177.640 -249.925 -177.470 ;
        RECT -259.545 -178.175 -259.375 -178.005 ;
        RECT -250.565 -178.175 -250.395 -178.005 ;
        RECT -259.545 -178.635 -259.375 -178.465 ;
        RECT -250.565 -178.635 -250.395 -178.465 ;
        RECT -249.625 -177.715 -249.455 -177.545 ;
        RECT -240.645 -177.715 -240.475 -177.545 ;
        RECT -240.175 -177.640 -240.005 -177.470 ;
        RECT -249.625 -178.175 -249.455 -178.005 ;
        RECT -240.645 -178.175 -240.475 -178.005 ;
        RECT -249.625 -178.635 -249.455 -178.465 ;
        RECT -240.645 -178.635 -240.475 -178.465 ;
        RECT -239.705 -177.715 -239.535 -177.545 ;
        RECT -230.725 -177.715 -230.555 -177.545 ;
        RECT -230.255 -177.640 -230.085 -177.470 ;
        RECT -239.705 -178.175 -239.535 -178.005 ;
        RECT -230.725 -178.175 -230.555 -178.005 ;
        RECT -239.705 -178.635 -239.535 -178.465 ;
        RECT -230.725 -178.635 -230.555 -178.465 ;
        RECT -229.785 -177.715 -229.615 -177.545 ;
        RECT -220.805 -177.715 -220.635 -177.545 ;
        RECT -220.335 -177.640 -220.165 -177.470 ;
        RECT -229.785 -178.175 -229.615 -178.005 ;
        RECT -220.805 -178.175 -220.635 -178.005 ;
        RECT -229.785 -178.635 -229.615 -178.465 ;
        RECT -220.805 -178.635 -220.635 -178.465 ;
        RECT -219.865 -177.715 -219.695 -177.545 ;
        RECT -210.885 -177.715 -210.715 -177.545 ;
        RECT -210.415 -177.640 -210.245 -177.470 ;
        RECT -219.865 -178.175 -219.695 -178.005 ;
        RECT -210.885 -178.175 -210.715 -178.005 ;
        RECT -219.865 -178.635 -219.695 -178.465 ;
        RECT -210.885 -178.635 -210.715 -178.465 ;
        RECT -209.945 -177.715 -209.775 -177.545 ;
        RECT -200.965 -177.715 -200.795 -177.545 ;
        RECT -200.495 -177.640 -200.325 -177.470 ;
        RECT -209.945 -178.175 -209.775 -178.005 ;
        RECT -200.965 -178.175 -200.795 -178.005 ;
        RECT -209.945 -178.635 -209.775 -178.465 ;
        RECT -200.965 -178.635 -200.795 -178.465 ;
        RECT -200.025 -177.715 -199.855 -177.545 ;
        RECT -191.045 -177.715 -190.875 -177.545 ;
        RECT -190.575 -177.640 -190.405 -177.470 ;
        RECT -200.025 -178.175 -199.855 -178.005 ;
        RECT -191.045 -178.175 -190.875 -178.005 ;
        RECT -200.025 -178.635 -199.855 -178.465 ;
        RECT -191.045 -178.635 -190.875 -178.465 ;
        RECT -190.105 -177.715 -189.935 -177.545 ;
        RECT -181.125 -177.715 -180.955 -177.545 ;
        RECT -180.655 -177.640 -180.485 -177.470 ;
        RECT -190.105 -178.175 -189.935 -178.005 ;
        RECT -181.125 -178.175 -180.955 -178.005 ;
        RECT -190.105 -178.635 -189.935 -178.465 ;
        RECT -181.125 -178.635 -180.955 -178.465 ;
        RECT -180.185 -177.715 -180.015 -177.545 ;
        RECT -171.205 -177.715 -171.035 -177.545 ;
        RECT -170.735 -177.640 -170.565 -177.470 ;
        RECT -180.185 -178.175 -180.015 -178.005 ;
        RECT -171.205 -178.175 -171.035 -178.005 ;
        RECT -180.185 -178.635 -180.015 -178.465 ;
        RECT -171.205 -178.635 -171.035 -178.465 ;
        RECT -170.265 -177.715 -170.095 -177.545 ;
        RECT -161.285 -177.715 -161.115 -177.545 ;
        RECT -160.815 -177.640 -160.645 -177.470 ;
        RECT -170.265 -178.175 -170.095 -178.005 ;
        RECT -161.285 -178.175 -161.115 -178.005 ;
        RECT -170.265 -178.635 -170.095 -178.465 ;
        RECT -161.285 -178.635 -161.115 -178.465 ;
        RECT -160.345 -177.715 -160.175 -177.545 ;
        RECT -151.365 -177.715 -151.195 -177.545 ;
        RECT -150.895 -177.640 -150.725 -177.470 ;
        RECT -160.345 -178.175 -160.175 -178.005 ;
        RECT -151.365 -178.175 -151.195 -178.005 ;
        RECT -160.345 -178.635 -160.175 -178.465 ;
        RECT -151.365 -178.635 -151.195 -178.465 ;
        RECT -150.425 -177.715 -150.255 -177.545 ;
        RECT -141.445 -177.715 -141.275 -177.545 ;
        RECT -140.975 -177.640 -140.805 -177.470 ;
        RECT -150.425 -178.175 -150.255 -178.005 ;
        RECT -141.445 -178.175 -141.275 -178.005 ;
        RECT -150.425 -178.635 -150.255 -178.465 ;
        RECT -141.445 -178.635 -141.275 -178.465 ;
        RECT -140.505 -177.715 -140.335 -177.545 ;
        RECT -131.525 -177.715 -131.355 -177.545 ;
        RECT -131.055 -177.640 -130.885 -177.470 ;
        RECT -140.505 -178.175 -140.335 -178.005 ;
        RECT -131.525 -178.175 -131.355 -178.005 ;
        RECT -140.505 -178.635 -140.335 -178.465 ;
        RECT -131.525 -178.635 -131.355 -178.465 ;
        RECT -130.585 -177.715 -130.415 -177.545 ;
        RECT -121.605 -177.715 -121.435 -177.545 ;
        RECT -121.135 -177.640 -120.965 -177.470 ;
        RECT -130.585 -178.175 -130.415 -178.005 ;
        RECT -121.605 -178.175 -121.435 -178.005 ;
        RECT -130.585 -178.635 -130.415 -178.465 ;
        RECT -121.605 -178.635 -121.435 -178.465 ;
        RECT -120.665 -177.715 -120.495 -177.545 ;
        RECT -111.685 -177.715 -111.515 -177.545 ;
        RECT -111.215 -177.640 -111.045 -177.470 ;
        RECT -120.665 -178.175 -120.495 -178.005 ;
        RECT -111.685 -178.175 -111.515 -178.005 ;
        RECT -120.665 -178.635 -120.495 -178.465 ;
        RECT -111.685 -178.635 -111.515 -178.465 ;
        RECT -110.745 -177.715 -110.575 -177.545 ;
        RECT -101.765 -177.715 -101.595 -177.545 ;
        RECT -101.295 -177.640 -101.125 -177.470 ;
        RECT -110.745 -178.175 -110.575 -178.005 ;
        RECT -101.765 -178.175 -101.595 -178.005 ;
        RECT -110.745 -178.635 -110.575 -178.465 ;
        RECT -101.765 -178.635 -101.595 -178.465 ;
        RECT -100.825 -177.715 -100.655 -177.545 ;
        RECT -91.845 -177.715 -91.675 -177.545 ;
        RECT -91.375 -177.640 -91.205 -177.470 ;
        RECT -100.825 -178.175 -100.655 -178.005 ;
        RECT -91.845 -178.175 -91.675 -178.005 ;
        RECT -100.825 -178.635 -100.655 -178.465 ;
        RECT -91.845 -178.635 -91.675 -178.465 ;
        RECT -90.905 -177.715 -90.735 -177.545 ;
        RECT -81.925 -177.715 -81.755 -177.545 ;
        RECT -81.455 -177.640 -81.285 -177.470 ;
        RECT -90.905 -178.175 -90.735 -178.005 ;
        RECT -81.925 -178.175 -81.755 -178.005 ;
        RECT -90.905 -178.635 -90.735 -178.465 ;
        RECT -81.925 -178.635 -81.755 -178.465 ;
        RECT -80.985 -177.715 -80.815 -177.545 ;
        RECT -72.005 -177.715 -71.835 -177.545 ;
        RECT -71.535 -177.640 -71.365 -177.470 ;
        RECT -80.985 -178.175 -80.815 -178.005 ;
        RECT -72.005 -178.175 -71.835 -178.005 ;
        RECT -80.985 -178.635 -80.815 -178.465 ;
        RECT -72.005 -178.635 -71.835 -178.465 ;
        RECT -71.065 -177.715 -70.895 -177.545 ;
        RECT -62.085 -177.715 -61.915 -177.545 ;
        RECT -61.615 -177.640 -61.445 -177.470 ;
        RECT -71.065 -178.175 -70.895 -178.005 ;
        RECT -62.085 -178.175 -61.915 -178.005 ;
        RECT -71.065 -178.635 -70.895 -178.465 ;
        RECT -62.085 -178.635 -61.915 -178.465 ;
        RECT -61.145 -177.715 -60.975 -177.545 ;
        RECT -52.165 -177.715 -51.995 -177.545 ;
        RECT -51.695 -177.640 -51.525 -177.470 ;
        RECT -61.145 -178.175 -60.975 -178.005 ;
        RECT -52.165 -178.175 -51.995 -178.005 ;
        RECT -61.145 -178.635 -60.975 -178.465 ;
        RECT -52.165 -178.635 -51.995 -178.465 ;
        RECT -51.225 -177.715 -51.055 -177.545 ;
        RECT -42.245 -177.715 -42.075 -177.545 ;
        RECT -41.775 -177.640 -41.605 -177.470 ;
        RECT -51.225 -178.175 -51.055 -178.005 ;
        RECT -42.245 -178.175 -42.075 -178.005 ;
        RECT -51.225 -178.635 -51.055 -178.465 ;
        RECT -42.245 -178.635 -42.075 -178.465 ;
        RECT -41.305 -177.715 -41.135 -177.545 ;
        RECT -32.325 -177.715 -32.155 -177.545 ;
        RECT -31.855 -177.640 -31.685 -177.470 ;
        RECT -41.305 -178.175 -41.135 -178.005 ;
        RECT -32.325 -178.175 -32.155 -178.005 ;
        RECT -41.305 -178.635 -41.135 -178.465 ;
        RECT -32.325 -178.635 -32.155 -178.465 ;
        RECT -31.385 -177.715 -31.215 -177.545 ;
        RECT -22.405 -177.715 -22.235 -177.545 ;
        RECT -21.935 -177.640 -21.765 -177.470 ;
        RECT -31.385 -178.175 -31.215 -178.005 ;
        RECT -22.405 -178.175 -22.235 -178.005 ;
        RECT -31.385 -178.635 -31.215 -178.465 ;
        RECT -22.405 -178.635 -22.235 -178.465 ;
        RECT -21.465 -177.715 -21.295 -177.545 ;
        RECT -12.485 -177.715 -12.315 -177.545 ;
        RECT -12.015 -177.640 -11.845 -177.470 ;
        RECT -21.465 -178.175 -21.295 -178.005 ;
        RECT -12.485 -178.175 -12.315 -178.005 ;
        RECT -21.465 -178.635 -21.295 -178.465 ;
        RECT -12.485 -178.635 -12.315 -178.465 ;
        RECT -11.545 -177.715 -11.375 -177.545 ;
        RECT -2.565 -177.715 -2.395 -177.545 ;
        RECT -2.095 -177.640 -1.925 -177.470 ;
        RECT -11.545 -178.175 -11.375 -178.005 ;
        RECT -2.565 -178.175 -2.395 -178.005 ;
        RECT -11.545 -178.635 -11.375 -178.465 ;
        RECT -2.565 -178.635 -2.395 -178.465 ;
        RECT -1.625 -177.715 -1.455 -177.545 ;
        RECT 7.355 -177.715 7.525 -177.545 ;
        RECT 7.825 -177.640 7.995 -177.470 ;
        RECT -1.625 -178.175 -1.455 -178.005 ;
        RECT 7.355 -178.175 7.525 -178.005 ;
        RECT -1.625 -178.635 -1.455 -178.465 ;
        RECT 7.355 -178.635 7.525 -178.465 ;
        RECT 8.295 -177.715 8.465 -177.545 ;
        RECT 17.275 -177.715 17.445 -177.545 ;
        RECT 17.745 -177.640 17.915 -177.470 ;
        RECT 8.295 -178.175 8.465 -178.005 ;
        RECT 17.275 -178.175 17.445 -178.005 ;
        RECT 8.295 -178.635 8.465 -178.465 ;
        RECT 17.275 -178.635 17.445 -178.465 ;
        RECT 18.215 -177.715 18.385 -177.545 ;
        RECT 18.215 -178.175 18.385 -178.005 ;
        RECT 18.215 -178.635 18.385 -178.465 ;
      LAYER met1 ;
        RECT -281.540 95.140 -281.080 95.145 ;
        RECT -271.620 95.140 -271.160 95.145 ;
        RECT -261.700 95.140 -261.240 95.145 ;
        RECT -251.780 95.140 -251.320 95.145 ;
        RECT -241.860 95.140 -241.400 95.145 ;
        RECT -231.940 95.140 -231.480 95.145 ;
        RECT -222.020 95.140 -221.560 95.145 ;
        RECT -212.100 95.140 -211.640 95.145 ;
        RECT -202.180 95.140 -201.720 95.145 ;
        RECT -192.260 95.140 -191.800 95.145 ;
        RECT -182.340 95.140 -181.880 95.145 ;
        RECT -172.420 95.140 -171.960 95.145 ;
        RECT -162.500 95.140 -162.040 95.145 ;
        RECT -152.580 95.140 -152.120 95.145 ;
        RECT -142.660 95.140 -142.200 95.145 ;
        RECT -132.740 95.140 -132.280 95.145 ;
        RECT -122.820 95.140 -122.360 95.145 ;
        RECT -112.900 95.140 -112.440 95.145 ;
        RECT -102.980 95.140 -102.520 95.145 ;
        RECT -93.060 95.140 -92.600 95.145 ;
        RECT -83.140 95.140 -82.680 95.145 ;
        RECT -73.220 95.140 -72.760 95.145 ;
        RECT -63.300 95.140 -62.840 95.145 ;
        RECT -53.380 95.140 -52.920 95.145 ;
        RECT -43.460 95.140 -43.000 95.145 ;
        RECT -33.540 95.140 -33.080 95.145 ;
        RECT -23.620 95.140 -23.160 95.145 ;
        RECT -13.700 95.140 -13.240 95.145 ;
        RECT -3.780 95.140 -3.320 95.145 ;
        RECT 6.140 95.140 6.600 95.145 ;
        RECT 16.060 95.140 16.520 95.145 ;
        RECT 25.980 95.140 26.440 95.145 ;
        RECT -282.020 93.760 -280.600 95.140 ;
        RECT -272.100 93.760 -270.680 95.140 ;
        RECT -262.180 93.760 -260.760 95.140 ;
        RECT -252.260 93.760 -250.840 95.140 ;
        RECT -242.340 93.760 -240.920 95.140 ;
        RECT -232.420 93.760 -231.000 95.140 ;
        RECT -222.500 93.760 -221.080 95.140 ;
        RECT -212.580 93.760 -211.160 95.140 ;
        RECT -202.660 93.760 -201.240 95.140 ;
        RECT -192.740 93.760 -191.320 95.140 ;
        RECT -182.820 93.760 -181.400 95.140 ;
        RECT -172.900 93.760 -171.480 95.140 ;
        RECT -162.980 93.760 -161.560 95.140 ;
        RECT -153.060 93.760 -151.640 95.140 ;
        RECT -143.140 93.760 -141.720 95.140 ;
        RECT -133.220 93.760 -131.800 95.140 ;
        RECT -123.300 93.760 -121.880 95.140 ;
        RECT -113.380 93.760 -111.960 95.140 ;
        RECT -103.460 93.760 -102.040 95.140 ;
        RECT -93.540 93.760 -92.120 95.140 ;
        RECT -83.620 93.760 -82.200 95.140 ;
        RECT -73.700 93.760 -72.280 95.140 ;
        RECT -63.780 93.760 -62.360 95.140 ;
        RECT -53.860 93.760 -52.440 95.140 ;
        RECT -43.940 93.760 -42.520 95.140 ;
        RECT -34.020 93.760 -32.600 95.140 ;
        RECT -24.100 93.760 -22.680 95.140 ;
        RECT -14.180 93.760 -12.760 95.140 ;
        RECT -4.260 93.760 -2.840 95.140 ;
        RECT 5.660 93.760 7.080 95.140 ;
        RECT 15.580 93.760 17.000 95.140 ;
        RECT 25.500 93.760 26.440 95.140 ;
        RECT -287.880 93.090 -284.660 93.570 ;
        RECT -277.960 93.090 -274.740 93.570 ;
        RECT -268.040 93.090 -264.820 93.570 ;
        RECT -258.120 93.090 -254.900 93.570 ;
        RECT -248.200 93.090 -244.980 93.570 ;
        RECT -238.280 93.090 -235.060 93.570 ;
        RECT -228.360 93.090 -225.140 93.570 ;
        RECT -218.440 93.090 -215.220 93.570 ;
        RECT -208.520 93.090 -205.300 93.570 ;
        RECT -198.600 93.090 -195.380 93.570 ;
        RECT -188.680 93.090 -185.460 93.570 ;
        RECT -178.760 93.090 -175.540 93.570 ;
        RECT -168.840 93.090 -165.620 93.570 ;
        RECT -158.920 93.090 -155.700 93.570 ;
        RECT -149.000 93.090 -145.780 93.570 ;
        RECT -139.080 93.090 -135.860 93.570 ;
        RECT -129.160 93.090 -125.940 93.570 ;
        RECT -119.240 93.090 -116.020 93.570 ;
        RECT -109.320 93.090 -106.100 93.570 ;
        RECT -99.400 93.090 -96.180 93.570 ;
        RECT -89.480 93.090 -86.260 93.570 ;
        RECT -79.560 93.090 -76.340 93.570 ;
        RECT -69.640 93.090 -66.420 93.570 ;
        RECT -59.720 93.090 -56.500 93.570 ;
        RECT -49.800 93.090 -46.580 93.570 ;
        RECT -39.880 93.090 -36.660 93.570 ;
        RECT -29.960 93.090 -26.740 93.570 ;
        RECT -20.040 93.090 -16.820 93.570 ;
        RECT -10.120 93.090 -6.900 93.570 ;
        RECT -0.200 93.090 3.020 93.570 ;
        RECT 9.720 93.090 12.940 93.570 ;
        RECT 19.640 93.090 22.860 93.570 ;
        RECT -282.920 90.370 -279.700 90.850 ;
        RECT -273.000 90.370 -269.780 90.850 ;
        RECT -263.080 90.370 -259.860 90.850 ;
        RECT -253.160 90.370 -249.940 90.850 ;
        RECT -243.240 90.370 -240.020 90.850 ;
        RECT -233.320 90.370 -230.100 90.850 ;
        RECT -223.400 90.370 -220.180 90.850 ;
        RECT -213.480 90.370 -210.260 90.850 ;
        RECT -203.560 90.370 -200.340 90.850 ;
        RECT -193.640 90.370 -190.420 90.850 ;
        RECT -183.720 90.370 -180.500 90.850 ;
        RECT -173.800 90.370 -170.580 90.850 ;
        RECT -163.880 90.370 -160.660 90.850 ;
        RECT -153.960 90.370 -150.740 90.850 ;
        RECT -144.040 90.370 -140.820 90.850 ;
        RECT -134.120 90.370 -130.900 90.850 ;
        RECT -124.200 90.370 -120.980 90.850 ;
        RECT -114.280 90.370 -111.060 90.850 ;
        RECT -104.360 90.370 -101.140 90.850 ;
        RECT -94.440 90.370 -91.220 90.850 ;
        RECT -84.520 90.370 -81.300 90.850 ;
        RECT -74.600 90.370 -71.380 90.850 ;
        RECT -64.680 90.370 -61.460 90.850 ;
        RECT -54.760 90.370 -51.540 90.850 ;
        RECT -44.840 90.370 -41.620 90.850 ;
        RECT -34.920 90.370 -31.700 90.850 ;
        RECT -25.000 90.370 -21.780 90.850 ;
        RECT -15.080 90.370 -11.860 90.850 ;
        RECT -5.160 90.370 -1.940 90.850 ;
        RECT 4.760 90.370 7.980 90.850 ;
        RECT 14.680 90.370 17.900 90.850 ;
        RECT 24.600 90.370 26.440 90.850 ;
        RECT -286.980 88.800 -285.560 90.180 ;
        RECT -277.060 88.800 -275.640 90.180 ;
        RECT -267.140 88.800 -265.720 90.180 ;
        RECT -257.220 88.800 -255.800 90.180 ;
        RECT -247.300 88.800 -245.880 90.180 ;
        RECT -237.380 88.800 -235.960 90.180 ;
        RECT -227.460 88.800 -226.040 90.180 ;
        RECT -217.540 88.800 -216.120 90.180 ;
        RECT -207.620 88.800 -206.200 90.180 ;
        RECT -197.700 88.800 -196.280 90.180 ;
        RECT -187.780 88.800 -186.360 90.180 ;
        RECT -177.860 88.800 -176.440 90.180 ;
        RECT -167.940 88.800 -166.520 90.180 ;
        RECT -158.020 88.800 -156.600 90.180 ;
        RECT -148.100 88.800 -146.680 90.180 ;
        RECT -138.180 88.800 -136.760 90.180 ;
        RECT -128.260 88.800 -126.840 90.180 ;
        RECT -118.340 88.800 -116.920 90.180 ;
        RECT -108.420 88.800 -107.000 90.180 ;
        RECT -98.500 88.800 -97.080 90.180 ;
        RECT -88.580 88.800 -87.160 90.180 ;
        RECT -78.660 88.800 -77.240 90.180 ;
        RECT -68.740 88.800 -67.320 90.180 ;
        RECT -58.820 88.800 -57.400 90.180 ;
        RECT -48.900 88.800 -47.480 90.180 ;
        RECT -38.980 88.800 -37.560 90.180 ;
        RECT -29.060 88.800 -27.640 90.180 ;
        RECT -19.140 88.800 -17.720 90.180 ;
        RECT -9.220 88.800 -7.800 90.180 ;
        RECT 0.700 88.800 2.120 90.180 ;
        RECT 10.620 88.800 12.040 90.180 ;
        RECT 20.540 88.800 21.960 90.180 ;
        RECT -283.560 11.090 -283.100 11.095 ;
        RECT -273.640 11.090 -273.180 11.095 ;
        RECT -263.720 11.090 -263.260 11.095 ;
        RECT -253.800 11.090 -253.340 11.095 ;
        RECT -243.880 11.090 -243.420 11.095 ;
        RECT -233.960 11.090 -233.500 11.095 ;
        RECT -224.040 11.090 -223.580 11.095 ;
        RECT -214.120 11.090 -213.660 11.095 ;
        RECT -204.200 11.090 -203.740 11.095 ;
        RECT -194.280 11.090 -193.820 11.095 ;
        RECT -184.360 11.090 -183.900 11.095 ;
        RECT -174.440 11.090 -173.980 11.095 ;
        RECT -164.520 11.090 -164.060 11.095 ;
        RECT -154.600 11.090 -154.140 11.095 ;
        RECT -144.680 11.090 -144.220 11.095 ;
        RECT -134.760 11.090 -134.300 11.095 ;
        RECT -124.840 11.090 -124.380 11.095 ;
        RECT -114.920 11.090 -114.460 11.095 ;
        RECT -105.000 11.090 -104.540 11.095 ;
        RECT -95.080 11.090 -94.620 11.095 ;
        RECT -85.160 11.090 -84.700 11.095 ;
        RECT -75.240 11.090 -74.780 11.095 ;
        RECT -65.320 11.090 -64.860 11.095 ;
        RECT -55.400 11.090 -54.940 11.095 ;
        RECT -45.480 11.090 -45.020 11.095 ;
        RECT -35.560 11.090 -35.100 11.095 ;
        RECT -25.640 11.090 -25.180 11.095 ;
        RECT -15.720 11.090 -15.260 11.095 ;
        RECT -5.800 11.090 -5.340 11.095 ;
        RECT 4.120 11.090 4.580 11.095 ;
        RECT 14.040 11.090 14.500 11.095 ;
        RECT 23.960 11.090 24.420 11.095 ;
        RECT -284.040 9.710 -282.620 11.090 ;
        RECT -274.120 9.710 -272.700 11.090 ;
        RECT -264.200 9.710 -262.780 11.090 ;
        RECT -254.280 9.710 -252.860 11.090 ;
        RECT -244.360 9.710 -242.940 11.090 ;
        RECT -234.440 9.710 -233.020 11.090 ;
        RECT -224.520 9.710 -223.100 11.090 ;
        RECT -214.600 9.710 -213.180 11.090 ;
        RECT -204.680 9.710 -203.260 11.090 ;
        RECT -194.760 9.710 -193.340 11.090 ;
        RECT -184.840 9.710 -183.420 11.090 ;
        RECT -174.920 9.710 -173.500 11.090 ;
        RECT -165.000 9.710 -163.580 11.090 ;
        RECT -155.080 9.710 -153.660 11.090 ;
        RECT -145.160 9.710 -143.740 11.090 ;
        RECT -135.240 9.710 -133.820 11.090 ;
        RECT -125.320 9.710 -123.900 11.090 ;
        RECT -115.400 9.710 -113.980 11.090 ;
        RECT -105.480 9.710 -104.060 11.090 ;
        RECT -95.560 9.710 -94.140 11.090 ;
        RECT -85.640 9.710 -84.220 11.090 ;
        RECT -75.720 9.710 -74.300 11.090 ;
        RECT -65.800 9.710 -64.380 11.090 ;
        RECT -55.880 9.710 -54.460 11.090 ;
        RECT -45.960 9.710 -44.540 11.090 ;
        RECT -36.040 9.710 -34.620 11.090 ;
        RECT -26.120 9.710 -24.700 11.090 ;
        RECT -16.200 9.710 -14.780 11.090 ;
        RECT -6.280 9.710 -4.860 11.090 ;
        RECT 3.640 9.710 5.060 11.090 ;
        RECT 13.560 9.710 14.980 11.090 ;
        RECT 23.480 9.710 24.420 11.090 ;
        RECT -289.900 9.040 -286.680 9.520 ;
        RECT -279.980 9.040 -276.760 9.520 ;
        RECT -270.060 9.040 -266.840 9.520 ;
        RECT -260.140 9.040 -256.920 9.520 ;
        RECT -250.220 9.040 -247.000 9.520 ;
        RECT -240.300 9.040 -237.080 9.520 ;
        RECT -230.380 9.040 -227.160 9.520 ;
        RECT -220.460 9.040 -217.240 9.520 ;
        RECT -210.540 9.040 -207.320 9.520 ;
        RECT -200.620 9.040 -197.400 9.520 ;
        RECT -190.700 9.040 -187.480 9.520 ;
        RECT -180.780 9.040 -177.560 9.520 ;
        RECT -170.860 9.040 -167.640 9.520 ;
        RECT -160.940 9.040 -157.720 9.520 ;
        RECT -151.020 9.040 -147.800 9.520 ;
        RECT -141.100 9.040 -137.880 9.520 ;
        RECT -131.180 9.040 -127.960 9.520 ;
        RECT -121.260 9.040 -118.040 9.520 ;
        RECT -111.340 9.040 -108.120 9.520 ;
        RECT -101.420 9.040 -98.200 9.520 ;
        RECT -91.500 9.040 -88.280 9.520 ;
        RECT -81.580 9.040 -78.360 9.520 ;
        RECT -71.660 9.040 -68.440 9.520 ;
        RECT -61.740 9.040 -58.520 9.520 ;
        RECT -51.820 9.040 -48.600 9.520 ;
        RECT -41.900 9.040 -38.680 9.520 ;
        RECT -31.980 9.040 -28.760 9.520 ;
        RECT -22.060 9.040 -18.840 9.520 ;
        RECT -12.140 9.040 -8.920 9.520 ;
        RECT -2.220 9.040 1.000 9.520 ;
        RECT 7.700 9.040 10.920 9.520 ;
        RECT 17.620 9.040 20.840 9.520 ;
        RECT -284.940 6.320 -281.720 6.800 ;
        RECT -275.020 6.320 -271.800 6.800 ;
        RECT -265.100 6.320 -261.880 6.800 ;
        RECT -255.180 6.320 -251.960 6.800 ;
        RECT -245.260 6.320 -242.040 6.800 ;
        RECT -235.340 6.320 -232.120 6.800 ;
        RECT -225.420 6.320 -222.200 6.800 ;
        RECT -215.500 6.320 -212.280 6.800 ;
        RECT -205.580 6.320 -202.360 6.800 ;
        RECT -195.660 6.320 -192.440 6.800 ;
        RECT -185.740 6.320 -182.520 6.800 ;
        RECT -175.820 6.320 -172.600 6.800 ;
        RECT -165.900 6.320 -162.680 6.800 ;
        RECT -155.980 6.320 -152.760 6.800 ;
        RECT -146.060 6.320 -142.840 6.800 ;
        RECT -136.140 6.320 -132.920 6.800 ;
        RECT -126.220 6.320 -123.000 6.800 ;
        RECT -116.300 6.320 -113.080 6.800 ;
        RECT -106.380 6.320 -103.160 6.800 ;
        RECT -96.460 6.320 -93.240 6.800 ;
        RECT -86.540 6.320 -83.320 6.800 ;
        RECT -76.620 6.320 -73.400 6.800 ;
        RECT -66.700 6.320 -63.480 6.800 ;
        RECT -56.780 6.320 -53.560 6.800 ;
        RECT -46.860 6.320 -43.640 6.800 ;
        RECT -36.940 6.320 -33.720 6.800 ;
        RECT -27.020 6.320 -23.800 6.800 ;
        RECT -17.100 6.320 -13.880 6.800 ;
        RECT -7.180 6.320 -3.960 6.800 ;
        RECT 2.740 6.320 5.960 6.800 ;
        RECT 12.660 6.320 15.880 6.800 ;
        RECT 22.580 6.320 24.420 6.800 ;
        RECT -289.000 4.750 -287.580 6.130 ;
        RECT -279.080 4.750 -277.660 6.130 ;
        RECT -269.160 4.750 -267.740 6.130 ;
        RECT -259.240 4.750 -257.820 6.130 ;
        RECT -249.320 4.750 -247.900 6.130 ;
        RECT -239.400 4.750 -237.980 6.130 ;
        RECT -229.480 4.750 -228.060 6.130 ;
        RECT -219.560 4.750 -218.140 6.130 ;
        RECT -209.640 4.750 -208.220 6.130 ;
        RECT -199.720 4.750 -198.300 6.130 ;
        RECT -189.800 4.750 -188.380 6.130 ;
        RECT -179.880 4.750 -178.460 6.130 ;
        RECT -169.960 4.750 -168.540 6.130 ;
        RECT -160.040 4.750 -158.620 6.130 ;
        RECT -150.120 4.750 -148.700 6.130 ;
        RECT -140.200 4.750 -138.780 6.130 ;
        RECT -130.280 4.750 -128.860 6.130 ;
        RECT -120.360 4.750 -118.940 6.130 ;
        RECT -110.440 4.750 -109.020 6.130 ;
        RECT -100.520 4.750 -99.100 6.130 ;
        RECT -90.600 4.750 -89.180 6.130 ;
        RECT -80.680 4.750 -79.260 6.130 ;
        RECT -70.760 4.750 -69.340 6.130 ;
        RECT -60.840 4.750 -59.420 6.130 ;
        RECT -50.920 4.750 -49.500 6.130 ;
        RECT -41.000 4.750 -39.580 6.130 ;
        RECT -31.080 4.750 -29.660 6.130 ;
        RECT -21.160 4.750 -19.740 6.130 ;
        RECT -11.240 4.750 -9.820 6.130 ;
        RECT -1.320 4.750 0.100 6.130 ;
        RECT 8.600 4.750 10.020 6.130 ;
        RECT 18.520 4.750 19.940 6.130 ;
        RECT -283.200 -77.860 -282.740 -77.855 ;
        RECT -273.280 -77.860 -272.820 -77.855 ;
        RECT -263.360 -77.860 -262.900 -77.855 ;
        RECT -253.440 -77.860 -252.980 -77.855 ;
        RECT -243.520 -77.860 -243.060 -77.855 ;
        RECT -233.600 -77.860 -233.140 -77.855 ;
        RECT -223.680 -77.860 -223.220 -77.855 ;
        RECT -213.760 -77.860 -213.300 -77.855 ;
        RECT -203.840 -77.860 -203.380 -77.855 ;
        RECT -193.920 -77.860 -193.460 -77.855 ;
        RECT -184.000 -77.860 -183.540 -77.855 ;
        RECT -174.080 -77.860 -173.620 -77.855 ;
        RECT -164.160 -77.860 -163.700 -77.855 ;
        RECT -154.240 -77.860 -153.780 -77.855 ;
        RECT -144.320 -77.860 -143.860 -77.855 ;
        RECT -134.400 -77.860 -133.940 -77.855 ;
        RECT -124.480 -77.860 -124.020 -77.855 ;
        RECT -114.560 -77.860 -114.100 -77.855 ;
        RECT -104.640 -77.860 -104.180 -77.855 ;
        RECT -94.720 -77.860 -94.260 -77.855 ;
        RECT -84.800 -77.860 -84.340 -77.855 ;
        RECT -74.880 -77.860 -74.420 -77.855 ;
        RECT -64.960 -77.860 -64.500 -77.855 ;
        RECT -55.040 -77.860 -54.580 -77.855 ;
        RECT -45.120 -77.860 -44.660 -77.855 ;
        RECT -35.200 -77.860 -34.740 -77.855 ;
        RECT -25.280 -77.860 -24.820 -77.855 ;
        RECT -15.360 -77.860 -14.900 -77.855 ;
        RECT -5.440 -77.860 -4.980 -77.855 ;
        RECT 4.480 -77.860 4.940 -77.855 ;
        RECT 14.400 -77.860 14.860 -77.855 ;
        RECT 24.320 -77.860 24.780 -77.855 ;
        RECT -283.680 -79.240 -282.260 -77.860 ;
        RECT -273.760 -79.240 -272.340 -77.860 ;
        RECT -263.840 -79.240 -262.420 -77.860 ;
        RECT -253.920 -79.240 -252.500 -77.860 ;
        RECT -244.000 -79.240 -242.580 -77.860 ;
        RECT -234.080 -79.240 -232.660 -77.860 ;
        RECT -224.160 -79.240 -222.740 -77.860 ;
        RECT -214.240 -79.240 -212.820 -77.860 ;
        RECT -204.320 -79.240 -202.900 -77.860 ;
        RECT -194.400 -79.240 -192.980 -77.860 ;
        RECT -184.480 -79.240 -183.060 -77.860 ;
        RECT -174.560 -79.240 -173.140 -77.860 ;
        RECT -164.640 -79.240 -163.220 -77.860 ;
        RECT -154.720 -79.240 -153.300 -77.860 ;
        RECT -144.800 -79.240 -143.380 -77.860 ;
        RECT -134.880 -79.240 -133.460 -77.860 ;
        RECT -124.960 -79.240 -123.540 -77.860 ;
        RECT -115.040 -79.240 -113.620 -77.860 ;
        RECT -105.120 -79.240 -103.700 -77.860 ;
        RECT -95.200 -79.240 -93.780 -77.860 ;
        RECT -85.280 -79.240 -83.860 -77.860 ;
        RECT -75.360 -79.240 -73.940 -77.860 ;
        RECT -65.440 -79.240 -64.020 -77.860 ;
        RECT -55.520 -79.240 -54.100 -77.860 ;
        RECT -45.600 -79.240 -44.180 -77.860 ;
        RECT -35.680 -79.240 -34.260 -77.860 ;
        RECT -25.760 -79.240 -24.340 -77.860 ;
        RECT -15.840 -79.240 -14.420 -77.860 ;
        RECT -5.920 -79.240 -4.500 -77.860 ;
        RECT 4.000 -79.240 5.420 -77.860 ;
        RECT 13.920 -79.240 15.340 -77.860 ;
        RECT 23.840 -79.240 24.780 -77.860 ;
        RECT -289.540 -79.910 -286.320 -79.430 ;
        RECT -279.620 -79.910 -276.400 -79.430 ;
        RECT -269.700 -79.910 -266.480 -79.430 ;
        RECT -259.780 -79.910 -256.560 -79.430 ;
        RECT -249.860 -79.910 -246.640 -79.430 ;
        RECT -239.940 -79.910 -236.720 -79.430 ;
        RECT -230.020 -79.910 -226.800 -79.430 ;
        RECT -220.100 -79.910 -216.880 -79.430 ;
        RECT -210.180 -79.910 -206.960 -79.430 ;
        RECT -200.260 -79.910 -197.040 -79.430 ;
        RECT -190.340 -79.910 -187.120 -79.430 ;
        RECT -180.420 -79.910 -177.200 -79.430 ;
        RECT -170.500 -79.910 -167.280 -79.430 ;
        RECT -160.580 -79.910 -157.360 -79.430 ;
        RECT -150.660 -79.910 -147.440 -79.430 ;
        RECT -140.740 -79.910 -137.520 -79.430 ;
        RECT -130.820 -79.910 -127.600 -79.430 ;
        RECT -120.900 -79.910 -117.680 -79.430 ;
        RECT -110.980 -79.910 -107.760 -79.430 ;
        RECT -101.060 -79.910 -97.840 -79.430 ;
        RECT -91.140 -79.910 -87.920 -79.430 ;
        RECT -81.220 -79.910 -78.000 -79.430 ;
        RECT -71.300 -79.910 -68.080 -79.430 ;
        RECT -61.380 -79.910 -58.160 -79.430 ;
        RECT -51.460 -79.910 -48.240 -79.430 ;
        RECT -41.540 -79.910 -38.320 -79.430 ;
        RECT -31.620 -79.910 -28.400 -79.430 ;
        RECT -21.700 -79.910 -18.480 -79.430 ;
        RECT -11.780 -79.910 -8.560 -79.430 ;
        RECT -1.860 -79.910 1.360 -79.430 ;
        RECT 8.060 -79.910 11.280 -79.430 ;
        RECT 17.980 -79.910 21.200 -79.430 ;
        RECT -284.580 -82.630 -281.360 -82.150 ;
        RECT -274.660 -82.630 -271.440 -82.150 ;
        RECT -264.740 -82.630 -261.520 -82.150 ;
        RECT -254.820 -82.630 -251.600 -82.150 ;
        RECT -244.900 -82.630 -241.680 -82.150 ;
        RECT -234.980 -82.630 -231.760 -82.150 ;
        RECT -225.060 -82.630 -221.840 -82.150 ;
        RECT -215.140 -82.630 -211.920 -82.150 ;
        RECT -205.220 -82.630 -202.000 -82.150 ;
        RECT -195.300 -82.630 -192.080 -82.150 ;
        RECT -185.380 -82.630 -182.160 -82.150 ;
        RECT -175.460 -82.630 -172.240 -82.150 ;
        RECT -165.540 -82.630 -162.320 -82.150 ;
        RECT -155.620 -82.630 -152.400 -82.150 ;
        RECT -145.700 -82.630 -142.480 -82.150 ;
        RECT -135.780 -82.630 -132.560 -82.150 ;
        RECT -125.860 -82.630 -122.640 -82.150 ;
        RECT -115.940 -82.630 -112.720 -82.150 ;
        RECT -106.020 -82.630 -102.800 -82.150 ;
        RECT -96.100 -82.630 -92.880 -82.150 ;
        RECT -86.180 -82.630 -82.960 -82.150 ;
        RECT -76.260 -82.630 -73.040 -82.150 ;
        RECT -66.340 -82.630 -63.120 -82.150 ;
        RECT -56.420 -82.630 -53.200 -82.150 ;
        RECT -46.500 -82.630 -43.280 -82.150 ;
        RECT -36.580 -82.630 -33.360 -82.150 ;
        RECT -26.660 -82.630 -23.440 -82.150 ;
        RECT -16.740 -82.630 -13.520 -82.150 ;
        RECT -6.820 -82.630 -3.600 -82.150 ;
        RECT 3.100 -82.630 6.320 -82.150 ;
        RECT 13.020 -82.630 16.240 -82.150 ;
        RECT 22.940 -82.630 24.780 -82.150 ;
        RECT -288.640 -84.200 -287.220 -82.820 ;
        RECT -278.720 -84.200 -277.300 -82.820 ;
        RECT -268.800 -84.200 -267.380 -82.820 ;
        RECT -258.880 -84.200 -257.460 -82.820 ;
        RECT -248.960 -84.200 -247.540 -82.820 ;
        RECT -239.040 -84.200 -237.620 -82.820 ;
        RECT -229.120 -84.200 -227.700 -82.820 ;
        RECT -219.200 -84.200 -217.780 -82.820 ;
        RECT -209.280 -84.200 -207.860 -82.820 ;
        RECT -199.360 -84.200 -197.940 -82.820 ;
        RECT -189.440 -84.200 -188.020 -82.820 ;
        RECT -179.520 -84.200 -178.100 -82.820 ;
        RECT -169.600 -84.200 -168.180 -82.820 ;
        RECT -159.680 -84.200 -158.260 -82.820 ;
        RECT -149.760 -84.200 -148.340 -82.820 ;
        RECT -139.840 -84.200 -138.420 -82.820 ;
        RECT -129.920 -84.200 -128.500 -82.820 ;
        RECT -120.000 -84.200 -118.580 -82.820 ;
        RECT -110.080 -84.200 -108.660 -82.820 ;
        RECT -100.160 -84.200 -98.740 -82.820 ;
        RECT -90.240 -84.200 -88.820 -82.820 ;
        RECT -80.320 -84.200 -78.900 -82.820 ;
        RECT -70.400 -84.200 -68.980 -82.820 ;
        RECT -60.480 -84.200 -59.060 -82.820 ;
        RECT -50.560 -84.200 -49.140 -82.820 ;
        RECT -40.640 -84.200 -39.220 -82.820 ;
        RECT -30.720 -84.200 -29.300 -82.820 ;
        RECT -20.800 -84.200 -19.380 -82.820 ;
        RECT -10.880 -84.200 -9.460 -82.820 ;
        RECT -0.960 -84.200 0.460 -82.820 ;
        RECT 8.960 -84.200 10.380 -82.820 ;
        RECT 18.880 -84.200 20.300 -82.820 ;
        RECT -284.960 -172.440 -284.500 -172.435 ;
        RECT -275.040 -172.440 -274.580 -172.435 ;
        RECT -265.120 -172.440 -264.660 -172.435 ;
        RECT -255.200 -172.440 -254.740 -172.435 ;
        RECT -245.280 -172.440 -244.820 -172.435 ;
        RECT -235.360 -172.440 -234.900 -172.435 ;
        RECT -225.440 -172.440 -224.980 -172.435 ;
        RECT -215.520 -172.440 -215.060 -172.435 ;
        RECT -205.600 -172.440 -205.140 -172.435 ;
        RECT -195.680 -172.440 -195.220 -172.435 ;
        RECT -185.760 -172.440 -185.300 -172.435 ;
        RECT -175.840 -172.440 -175.380 -172.435 ;
        RECT -165.920 -172.440 -165.460 -172.435 ;
        RECT -156.000 -172.440 -155.540 -172.435 ;
        RECT -146.080 -172.440 -145.620 -172.435 ;
        RECT -136.160 -172.440 -135.700 -172.435 ;
        RECT -126.240 -172.440 -125.780 -172.435 ;
        RECT -116.320 -172.440 -115.860 -172.435 ;
        RECT -106.400 -172.440 -105.940 -172.435 ;
        RECT -96.480 -172.440 -96.020 -172.435 ;
        RECT -86.560 -172.440 -86.100 -172.435 ;
        RECT -76.640 -172.440 -76.180 -172.435 ;
        RECT -66.720 -172.440 -66.260 -172.435 ;
        RECT -56.800 -172.440 -56.340 -172.435 ;
        RECT -46.880 -172.440 -46.420 -172.435 ;
        RECT -36.960 -172.440 -36.500 -172.435 ;
        RECT -27.040 -172.440 -26.580 -172.435 ;
        RECT -17.120 -172.440 -16.660 -172.435 ;
        RECT -7.200 -172.440 -6.740 -172.435 ;
        RECT 2.720 -172.440 3.180 -172.435 ;
        RECT 12.640 -172.440 13.100 -172.435 ;
        RECT 22.560 -172.440 23.020 -172.435 ;
        RECT -285.440 -173.820 -284.020 -172.440 ;
        RECT -275.520 -173.820 -274.100 -172.440 ;
        RECT -265.600 -173.820 -264.180 -172.440 ;
        RECT -255.680 -173.820 -254.260 -172.440 ;
        RECT -245.760 -173.820 -244.340 -172.440 ;
        RECT -235.840 -173.820 -234.420 -172.440 ;
        RECT -225.920 -173.820 -224.500 -172.440 ;
        RECT -216.000 -173.820 -214.580 -172.440 ;
        RECT -206.080 -173.820 -204.660 -172.440 ;
        RECT -196.160 -173.820 -194.740 -172.440 ;
        RECT -186.240 -173.820 -184.820 -172.440 ;
        RECT -176.320 -173.820 -174.900 -172.440 ;
        RECT -166.400 -173.820 -164.980 -172.440 ;
        RECT -156.480 -173.820 -155.060 -172.440 ;
        RECT -146.560 -173.820 -145.140 -172.440 ;
        RECT -136.640 -173.820 -135.220 -172.440 ;
        RECT -126.720 -173.820 -125.300 -172.440 ;
        RECT -116.800 -173.820 -115.380 -172.440 ;
        RECT -106.880 -173.820 -105.460 -172.440 ;
        RECT -96.960 -173.820 -95.540 -172.440 ;
        RECT -87.040 -173.820 -85.620 -172.440 ;
        RECT -77.120 -173.820 -75.700 -172.440 ;
        RECT -67.200 -173.820 -65.780 -172.440 ;
        RECT -57.280 -173.820 -55.860 -172.440 ;
        RECT -47.360 -173.820 -45.940 -172.440 ;
        RECT -37.440 -173.820 -36.020 -172.440 ;
        RECT -27.520 -173.820 -26.100 -172.440 ;
        RECT -17.600 -173.820 -16.180 -172.440 ;
        RECT -7.680 -173.820 -6.260 -172.440 ;
        RECT 2.240 -173.820 3.660 -172.440 ;
        RECT 12.160 -173.820 13.580 -172.440 ;
        RECT 22.080 -173.820 23.020 -172.440 ;
        RECT -291.300 -174.490 -288.080 -174.010 ;
        RECT -281.380 -174.490 -278.160 -174.010 ;
        RECT -271.460 -174.490 -268.240 -174.010 ;
        RECT -261.540 -174.490 -258.320 -174.010 ;
        RECT -251.620 -174.490 -248.400 -174.010 ;
        RECT -241.700 -174.490 -238.480 -174.010 ;
        RECT -231.780 -174.490 -228.560 -174.010 ;
        RECT -221.860 -174.490 -218.640 -174.010 ;
        RECT -211.940 -174.490 -208.720 -174.010 ;
        RECT -202.020 -174.490 -198.800 -174.010 ;
        RECT -192.100 -174.490 -188.880 -174.010 ;
        RECT -182.180 -174.490 -178.960 -174.010 ;
        RECT -172.260 -174.490 -169.040 -174.010 ;
        RECT -162.340 -174.490 -159.120 -174.010 ;
        RECT -152.420 -174.490 -149.200 -174.010 ;
        RECT -142.500 -174.490 -139.280 -174.010 ;
        RECT -132.580 -174.490 -129.360 -174.010 ;
        RECT -122.660 -174.490 -119.440 -174.010 ;
        RECT -112.740 -174.490 -109.520 -174.010 ;
        RECT -102.820 -174.490 -99.600 -174.010 ;
        RECT -92.900 -174.490 -89.680 -174.010 ;
        RECT -82.980 -174.490 -79.760 -174.010 ;
        RECT -73.060 -174.490 -69.840 -174.010 ;
        RECT -63.140 -174.490 -59.920 -174.010 ;
        RECT -53.220 -174.490 -50.000 -174.010 ;
        RECT -43.300 -174.490 -40.080 -174.010 ;
        RECT -33.380 -174.490 -30.160 -174.010 ;
        RECT -23.460 -174.490 -20.240 -174.010 ;
        RECT -13.540 -174.490 -10.320 -174.010 ;
        RECT -3.620 -174.490 -0.400 -174.010 ;
        RECT 6.300 -174.490 9.520 -174.010 ;
        RECT 16.220 -174.490 19.440 -174.010 ;
        RECT -286.340 -177.210 -283.120 -176.730 ;
        RECT -276.420 -177.210 -273.200 -176.730 ;
        RECT -266.500 -177.210 -263.280 -176.730 ;
        RECT -256.580 -177.210 -253.360 -176.730 ;
        RECT -246.660 -177.210 -243.440 -176.730 ;
        RECT -236.740 -177.210 -233.520 -176.730 ;
        RECT -226.820 -177.210 -223.600 -176.730 ;
        RECT -216.900 -177.210 -213.680 -176.730 ;
        RECT -206.980 -177.210 -203.760 -176.730 ;
        RECT -197.060 -177.210 -193.840 -176.730 ;
        RECT -187.140 -177.210 -183.920 -176.730 ;
        RECT -177.220 -177.210 -174.000 -176.730 ;
        RECT -167.300 -177.210 -164.080 -176.730 ;
        RECT -157.380 -177.210 -154.160 -176.730 ;
        RECT -147.460 -177.210 -144.240 -176.730 ;
        RECT -137.540 -177.210 -134.320 -176.730 ;
        RECT -127.620 -177.210 -124.400 -176.730 ;
        RECT -117.700 -177.210 -114.480 -176.730 ;
        RECT -107.780 -177.210 -104.560 -176.730 ;
        RECT -97.860 -177.210 -94.640 -176.730 ;
        RECT -87.940 -177.210 -84.720 -176.730 ;
        RECT -78.020 -177.210 -74.800 -176.730 ;
        RECT -68.100 -177.210 -64.880 -176.730 ;
        RECT -58.180 -177.210 -54.960 -176.730 ;
        RECT -48.260 -177.210 -45.040 -176.730 ;
        RECT -38.340 -177.210 -35.120 -176.730 ;
        RECT -28.420 -177.210 -25.200 -176.730 ;
        RECT -18.500 -177.210 -15.280 -176.730 ;
        RECT -8.580 -177.210 -5.360 -176.730 ;
        RECT 1.340 -177.210 4.560 -176.730 ;
        RECT 11.260 -177.210 14.480 -176.730 ;
        RECT 21.180 -177.210 23.020 -176.730 ;
        RECT -290.400 -178.780 -288.980 -177.400 ;
        RECT -280.480 -178.780 -279.060 -177.400 ;
        RECT -270.560 -178.780 -269.140 -177.400 ;
        RECT -260.640 -178.780 -259.220 -177.400 ;
        RECT -250.720 -178.780 -249.300 -177.400 ;
        RECT -240.800 -178.780 -239.380 -177.400 ;
        RECT -230.880 -178.780 -229.460 -177.400 ;
        RECT -220.960 -178.780 -219.540 -177.400 ;
        RECT -211.040 -178.780 -209.620 -177.400 ;
        RECT -201.120 -178.780 -199.700 -177.400 ;
        RECT -191.200 -178.780 -189.780 -177.400 ;
        RECT -181.280 -178.780 -179.860 -177.400 ;
        RECT -171.360 -178.780 -169.940 -177.400 ;
        RECT -161.440 -178.780 -160.020 -177.400 ;
        RECT -151.520 -178.780 -150.100 -177.400 ;
        RECT -141.600 -178.780 -140.180 -177.400 ;
        RECT -131.680 -178.780 -130.260 -177.400 ;
        RECT -121.760 -178.780 -120.340 -177.400 ;
        RECT -111.840 -178.780 -110.420 -177.400 ;
        RECT -101.920 -178.780 -100.500 -177.400 ;
        RECT -92.000 -178.780 -90.580 -177.400 ;
        RECT -82.080 -178.780 -80.660 -177.400 ;
        RECT -72.160 -178.780 -70.740 -177.400 ;
        RECT -62.240 -178.780 -60.820 -177.400 ;
        RECT -52.320 -178.780 -50.900 -177.400 ;
        RECT -42.400 -178.780 -40.980 -177.400 ;
        RECT -32.480 -178.780 -31.060 -177.400 ;
        RECT -22.560 -178.780 -21.140 -177.400 ;
        RECT -12.640 -178.780 -11.220 -177.400 ;
        RECT -2.720 -178.780 -1.300 -177.400 ;
        RECT 7.200 -178.780 8.620 -177.400 ;
        RECT 17.120 -178.780 18.540 -177.400 ;
      LAYER via ;
        RECT -281.920 94.780 -281.645 95.045 ;
        RECT -280.980 94.770 -280.705 95.035 ;
        RECT -271.290 95.035 -271.020 95.040 ;
        RECT -271.290 94.770 -270.785 95.035 ;
        RECT -262.080 94.780 -261.805 95.045 ;
        RECT -261.140 94.770 -260.865 95.035 ;
        RECT -252.160 94.780 -251.885 95.045 ;
        RECT -251.220 94.770 -250.945 95.035 ;
        RECT -242.240 94.780 -241.965 95.045 ;
        RECT -241.300 94.770 -241.025 95.035 ;
        RECT -232.320 94.780 -232.045 95.045 ;
        RECT -231.380 94.770 -231.105 95.035 ;
        RECT -222.400 94.780 -222.125 95.045 ;
        RECT -221.460 94.770 -221.185 95.035 ;
        RECT -212.480 94.780 -212.205 95.045 ;
        RECT -211.540 94.770 -211.265 95.035 ;
        RECT -202.560 94.780 -202.285 95.045 ;
        RECT -201.620 94.770 -201.345 95.035 ;
        RECT -192.640 94.780 -192.365 95.045 ;
        RECT -191.700 94.770 -191.425 95.035 ;
        RECT -182.720 94.780 -182.445 95.045 ;
        RECT -181.780 94.770 -181.505 95.035 ;
        RECT -172.800 94.780 -172.525 95.045 ;
        RECT -171.860 94.770 -171.585 95.035 ;
        RECT -162.880 94.780 -162.605 95.045 ;
        RECT -161.940 94.770 -161.665 95.035 ;
        RECT -152.960 94.780 -152.685 95.045 ;
        RECT -152.020 94.770 -151.745 95.035 ;
        RECT -143.040 94.780 -142.765 95.045 ;
        RECT -142.100 94.770 -141.825 95.035 ;
        RECT -133.120 94.780 -132.845 95.045 ;
        RECT -132.180 94.770 -131.905 95.035 ;
        RECT -123.200 94.780 -122.925 95.045 ;
        RECT -122.260 94.770 -121.985 95.035 ;
        RECT -113.280 94.780 -113.005 95.045 ;
        RECT -112.340 94.770 -112.065 95.035 ;
        RECT -103.360 94.780 -103.085 95.045 ;
        RECT -102.420 94.770 -102.145 95.035 ;
        RECT -93.440 94.780 -93.165 95.045 ;
        RECT -92.500 94.770 -92.225 95.035 ;
        RECT -83.520 94.780 -83.245 95.045 ;
        RECT -82.580 94.770 -82.305 95.035 ;
        RECT -73.600 94.780 -73.325 95.045 ;
        RECT -72.660 94.770 -72.385 95.035 ;
        RECT -63.680 94.780 -63.405 95.045 ;
        RECT -62.740 94.770 -62.465 95.035 ;
        RECT -53.760 94.780 -53.485 95.045 ;
        RECT -52.820 94.770 -52.545 95.035 ;
        RECT -43.840 94.780 -43.565 95.045 ;
        RECT -42.900 94.770 -42.625 95.035 ;
        RECT -33.920 94.780 -33.645 95.045 ;
        RECT -32.980 94.770 -32.705 95.035 ;
        RECT -24.000 94.780 -23.725 95.045 ;
        RECT -23.060 94.770 -22.785 95.035 ;
        RECT -14.080 94.780 -13.805 95.045 ;
        RECT -13.140 94.770 -12.865 95.035 ;
        RECT -4.160 94.780 -3.885 95.045 ;
        RECT -3.220 94.770 -2.945 95.035 ;
        RECT 5.760 94.780 6.035 95.045 ;
        RECT 6.700 94.770 6.975 95.035 ;
        RECT 15.680 94.780 15.955 95.045 ;
        RECT 16.620 94.770 16.895 95.035 ;
        RECT 25.600 94.780 25.875 95.045 ;
        RECT -286.640 93.190 -286.365 93.455 ;
        RECT -286.180 93.190 -285.905 93.455 ;
        RECT -276.720 93.190 -276.445 93.455 ;
        RECT -276.260 93.190 -275.985 93.455 ;
        RECT -266.800 93.190 -266.525 93.455 ;
        RECT -266.340 93.190 -266.065 93.455 ;
        RECT -256.880 93.190 -256.605 93.455 ;
        RECT -256.420 93.190 -256.145 93.455 ;
        RECT -246.960 93.190 -246.685 93.455 ;
        RECT -246.500 93.190 -246.225 93.455 ;
        RECT -237.040 93.190 -236.765 93.455 ;
        RECT -236.580 93.190 -236.305 93.455 ;
        RECT -227.120 93.190 -226.845 93.455 ;
        RECT -226.660 93.190 -226.385 93.455 ;
        RECT -217.200 93.190 -216.925 93.455 ;
        RECT -216.740 93.190 -216.465 93.455 ;
        RECT -207.280 93.190 -207.005 93.455 ;
        RECT -206.820 93.190 -206.545 93.455 ;
        RECT -197.360 93.190 -197.085 93.455 ;
        RECT -196.900 93.190 -196.625 93.455 ;
        RECT -187.440 93.190 -187.165 93.455 ;
        RECT -186.980 93.190 -186.705 93.455 ;
        RECT -177.520 93.190 -177.245 93.455 ;
        RECT -177.060 93.190 -176.785 93.455 ;
        RECT -167.600 93.190 -167.325 93.455 ;
        RECT -167.140 93.190 -166.865 93.455 ;
        RECT -157.680 93.190 -157.405 93.455 ;
        RECT -157.220 93.190 -156.945 93.455 ;
        RECT -147.760 93.190 -147.485 93.455 ;
        RECT -147.300 93.190 -147.025 93.455 ;
        RECT -137.840 93.190 -137.565 93.455 ;
        RECT -137.380 93.190 -137.105 93.455 ;
        RECT -127.920 93.190 -127.645 93.455 ;
        RECT -127.460 93.190 -127.185 93.455 ;
        RECT -118.000 93.190 -117.725 93.455 ;
        RECT -117.540 93.190 -117.265 93.455 ;
        RECT -108.080 93.190 -107.805 93.455 ;
        RECT -107.620 93.190 -107.345 93.455 ;
        RECT -98.160 93.190 -97.885 93.455 ;
        RECT -97.700 93.190 -97.425 93.455 ;
        RECT -88.240 93.190 -87.965 93.455 ;
        RECT -87.780 93.190 -87.505 93.455 ;
        RECT -78.320 93.190 -78.045 93.455 ;
        RECT -77.860 93.190 -77.585 93.455 ;
        RECT -68.400 93.190 -68.125 93.455 ;
        RECT -67.940 93.190 -67.665 93.455 ;
        RECT -58.480 93.190 -58.205 93.455 ;
        RECT -58.020 93.190 -57.745 93.455 ;
        RECT -48.560 93.190 -48.285 93.455 ;
        RECT -48.100 93.190 -47.825 93.455 ;
        RECT -38.640 93.190 -38.365 93.455 ;
        RECT -38.180 93.190 -37.905 93.455 ;
        RECT -28.720 93.190 -28.445 93.455 ;
        RECT -28.260 93.190 -27.985 93.455 ;
        RECT -18.800 93.190 -18.525 93.455 ;
        RECT -18.340 93.190 -18.065 93.455 ;
        RECT -8.880 93.190 -8.605 93.455 ;
        RECT -8.420 93.190 -8.145 93.455 ;
        RECT 1.040 93.190 1.315 93.455 ;
        RECT 1.500 93.190 1.775 93.455 ;
        RECT 10.960 93.190 11.235 93.455 ;
        RECT 11.420 93.190 11.695 93.455 ;
        RECT 20.880 93.190 21.155 93.455 ;
        RECT 21.340 93.190 21.615 93.455 ;
        RECT -281.680 90.480 -281.405 90.745 ;
        RECT -281.220 90.480 -280.945 90.745 ;
        RECT -271.760 90.480 -271.485 90.745 ;
        RECT -271.300 90.480 -271.025 90.745 ;
        RECT -261.840 90.480 -261.565 90.745 ;
        RECT -261.380 90.480 -261.105 90.745 ;
        RECT -251.920 90.480 -251.645 90.745 ;
        RECT -251.460 90.480 -251.185 90.745 ;
        RECT -242.000 90.480 -241.725 90.745 ;
        RECT -241.540 90.480 -241.265 90.745 ;
        RECT -232.080 90.480 -231.805 90.745 ;
        RECT -231.620 90.480 -231.345 90.745 ;
        RECT -222.160 90.480 -221.885 90.745 ;
        RECT -221.700 90.480 -221.425 90.745 ;
        RECT -212.240 90.480 -211.965 90.745 ;
        RECT -211.780 90.480 -211.505 90.745 ;
        RECT -202.320 90.480 -202.045 90.745 ;
        RECT -201.860 90.480 -201.585 90.745 ;
        RECT -192.400 90.480 -192.125 90.745 ;
        RECT -191.940 90.480 -191.665 90.745 ;
        RECT -182.480 90.480 -182.205 90.745 ;
        RECT -182.020 90.480 -181.745 90.745 ;
        RECT -172.560 90.480 -172.285 90.745 ;
        RECT -172.100 90.480 -171.825 90.745 ;
        RECT -162.640 90.480 -162.365 90.745 ;
        RECT -162.180 90.480 -161.905 90.745 ;
        RECT -152.720 90.480 -152.445 90.745 ;
        RECT -152.260 90.480 -151.985 90.745 ;
        RECT -142.800 90.480 -142.525 90.745 ;
        RECT -142.340 90.480 -142.065 90.745 ;
        RECT -132.880 90.480 -132.605 90.745 ;
        RECT -132.420 90.480 -132.145 90.745 ;
        RECT -122.960 90.480 -122.685 90.745 ;
        RECT -122.500 90.480 -122.225 90.745 ;
        RECT -113.040 90.480 -112.765 90.745 ;
        RECT -112.580 90.480 -112.305 90.745 ;
        RECT -103.120 90.480 -102.845 90.745 ;
        RECT -102.660 90.480 -102.385 90.745 ;
        RECT -93.200 90.480 -92.925 90.745 ;
        RECT -92.740 90.480 -92.465 90.745 ;
        RECT -83.280 90.480 -83.005 90.745 ;
        RECT -82.820 90.480 -82.545 90.745 ;
        RECT -73.360 90.480 -73.085 90.745 ;
        RECT -72.900 90.480 -72.625 90.745 ;
        RECT -63.440 90.480 -63.165 90.745 ;
        RECT -62.980 90.480 -62.705 90.745 ;
        RECT -53.520 90.480 -53.245 90.745 ;
        RECT -53.060 90.480 -52.785 90.745 ;
        RECT -43.600 90.480 -43.325 90.745 ;
        RECT -43.140 90.480 -42.865 90.745 ;
        RECT -33.680 90.480 -33.405 90.745 ;
        RECT -33.220 90.480 -32.945 90.745 ;
        RECT -23.760 90.480 -23.485 90.745 ;
        RECT -23.300 90.480 -23.025 90.745 ;
        RECT -13.840 90.480 -13.565 90.745 ;
        RECT -13.380 90.480 -13.105 90.745 ;
        RECT -3.920 90.480 -3.645 90.745 ;
        RECT -3.460 90.480 -3.185 90.745 ;
        RECT 6.000 90.480 6.275 90.745 ;
        RECT 6.460 90.480 6.735 90.745 ;
        RECT 15.920 90.480 16.195 90.745 ;
        RECT 16.380 90.480 16.655 90.745 ;
        RECT 25.840 90.480 26.115 90.745 ;
        RECT -286.870 88.890 -286.595 89.155 ;
        RECT -285.940 88.890 -285.665 89.155 ;
        RECT -276.950 88.890 -276.675 89.155 ;
        RECT -276.020 88.890 -275.745 89.155 ;
        RECT -267.030 88.890 -266.755 89.155 ;
        RECT -266.100 88.890 -265.825 89.155 ;
        RECT -257.110 88.890 -256.835 89.155 ;
        RECT -256.180 88.890 -255.905 89.155 ;
        RECT -247.190 88.890 -246.915 89.155 ;
        RECT -246.260 88.890 -245.985 89.155 ;
        RECT -237.270 88.890 -236.995 89.155 ;
        RECT -236.340 88.890 -236.065 89.155 ;
        RECT -227.350 88.890 -227.075 89.155 ;
        RECT -226.420 88.890 -226.145 89.155 ;
        RECT -217.430 88.890 -217.155 89.155 ;
        RECT -216.500 88.890 -216.225 89.155 ;
        RECT -207.510 88.890 -207.235 89.155 ;
        RECT -206.580 88.890 -206.305 89.155 ;
        RECT -197.590 88.890 -197.315 89.155 ;
        RECT -196.660 88.890 -196.385 89.155 ;
        RECT -187.670 88.890 -187.395 89.155 ;
        RECT -186.740 88.890 -186.465 89.155 ;
        RECT -177.750 88.890 -177.475 89.155 ;
        RECT -176.820 88.890 -176.545 89.155 ;
        RECT -167.830 88.890 -167.555 89.155 ;
        RECT -166.900 88.890 -166.625 89.155 ;
        RECT -157.910 88.890 -157.635 89.155 ;
        RECT -156.980 88.890 -156.705 89.155 ;
        RECT -147.990 88.890 -147.715 89.155 ;
        RECT -147.060 88.890 -146.785 89.155 ;
        RECT -138.070 88.890 -137.795 89.155 ;
        RECT -137.140 88.890 -136.865 89.155 ;
        RECT -128.150 88.890 -127.875 89.155 ;
        RECT -127.220 88.890 -126.945 89.155 ;
        RECT -118.230 88.890 -117.955 89.155 ;
        RECT -117.300 88.890 -117.025 89.155 ;
        RECT -108.310 88.890 -108.035 89.155 ;
        RECT -107.380 88.890 -107.105 89.155 ;
        RECT -98.390 88.890 -98.115 89.155 ;
        RECT -97.460 88.890 -97.185 89.155 ;
        RECT -88.470 88.890 -88.195 89.155 ;
        RECT -87.540 88.890 -87.265 89.155 ;
        RECT -78.550 88.890 -78.275 89.155 ;
        RECT -77.620 88.890 -77.345 89.155 ;
        RECT -68.630 88.890 -68.355 89.155 ;
        RECT -67.700 88.890 -67.425 89.155 ;
        RECT -58.710 88.890 -58.435 89.155 ;
        RECT -57.780 88.890 -57.505 89.155 ;
        RECT -48.790 88.890 -48.515 89.155 ;
        RECT -47.860 88.890 -47.585 89.155 ;
        RECT -38.870 88.890 -38.595 89.155 ;
        RECT -37.940 88.890 -37.665 89.155 ;
        RECT -28.950 88.890 -28.675 89.155 ;
        RECT -28.020 88.890 -27.745 89.155 ;
        RECT -19.030 88.890 -18.755 89.155 ;
        RECT -18.100 88.890 -17.825 89.155 ;
        RECT -9.110 88.890 -8.835 89.155 ;
        RECT -8.180 88.890 -7.905 89.155 ;
        RECT 0.810 88.890 1.085 89.155 ;
        RECT 1.740 88.890 2.015 89.155 ;
        RECT 10.730 88.890 11.005 89.155 ;
        RECT 11.660 88.890 11.935 89.155 ;
        RECT 20.650 88.890 20.925 89.155 ;
        RECT 21.580 88.890 21.855 89.155 ;
        RECT -283.940 10.730 -283.665 10.995 ;
        RECT -283.000 10.720 -282.725 10.985 ;
        RECT -273.310 10.985 -273.040 10.990 ;
        RECT -273.310 10.720 -272.805 10.985 ;
        RECT -264.100 10.730 -263.825 10.995 ;
        RECT -263.160 10.720 -262.885 10.985 ;
        RECT -254.180 10.730 -253.905 10.995 ;
        RECT -253.240 10.720 -252.965 10.985 ;
        RECT -244.260 10.730 -243.985 10.995 ;
        RECT -243.320 10.720 -243.045 10.985 ;
        RECT -234.340 10.730 -234.065 10.995 ;
        RECT -233.400 10.720 -233.125 10.985 ;
        RECT -224.420 10.730 -224.145 10.995 ;
        RECT -223.480 10.720 -223.205 10.985 ;
        RECT -214.500 10.730 -214.225 10.995 ;
        RECT -213.560 10.720 -213.285 10.985 ;
        RECT -204.580 10.730 -204.305 10.995 ;
        RECT -203.640 10.720 -203.365 10.985 ;
        RECT -194.660 10.730 -194.385 10.995 ;
        RECT -193.720 10.720 -193.445 10.985 ;
        RECT -184.740 10.730 -184.465 10.995 ;
        RECT -183.800 10.720 -183.525 10.985 ;
        RECT -174.820 10.730 -174.545 10.995 ;
        RECT -173.880 10.720 -173.605 10.985 ;
        RECT -164.900 10.730 -164.625 10.995 ;
        RECT -163.960 10.720 -163.685 10.985 ;
        RECT -154.980 10.730 -154.705 10.995 ;
        RECT -154.040 10.720 -153.765 10.985 ;
        RECT -145.060 10.730 -144.785 10.995 ;
        RECT -144.120 10.720 -143.845 10.985 ;
        RECT -135.140 10.730 -134.865 10.995 ;
        RECT -134.200 10.720 -133.925 10.985 ;
        RECT -125.220 10.730 -124.945 10.995 ;
        RECT -124.280 10.720 -124.005 10.985 ;
        RECT -115.300 10.730 -115.025 10.995 ;
        RECT -114.360 10.720 -114.085 10.985 ;
        RECT -105.380 10.730 -105.105 10.995 ;
        RECT -104.440 10.720 -104.165 10.985 ;
        RECT -95.460 10.730 -95.185 10.995 ;
        RECT -94.520 10.720 -94.245 10.985 ;
        RECT -85.540 10.730 -85.265 10.995 ;
        RECT -84.600 10.720 -84.325 10.985 ;
        RECT -75.620 10.730 -75.345 10.995 ;
        RECT -74.680 10.720 -74.405 10.985 ;
        RECT -65.700 10.730 -65.425 10.995 ;
        RECT -64.760 10.720 -64.485 10.985 ;
        RECT -55.780 10.730 -55.505 10.995 ;
        RECT -54.840 10.720 -54.565 10.985 ;
        RECT -45.860 10.730 -45.585 10.995 ;
        RECT -44.920 10.720 -44.645 10.985 ;
        RECT -35.940 10.730 -35.665 10.995 ;
        RECT -35.000 10.720 -34.725 10.985 ;
        RECT -26.020 10.730 -25.745 10.995 ;
        RECT -25.080 10.720 -24.805 10.985 ;
        RECT -16.100 10.730 -15.825 10.995 ;
        RECT -15.160 10.720 -14.885 10.985 ;
        RECT -6.180 10.730 -5.905 10.995 ;
        RECT -5.240 10.720 -4.965 10.985 ;
        RECT 3.740 10.730 4.015 10.995 ;
        RECT 4.680 10.720 4.955 10.985 ;
        RECT 13.660 10.730 13.935 10.995 ;
        RECT 14.600 10.720 14.875 10.985 ;
        RECT 23.580 10.730 23.855 10.995 ;
        RECT -288.660 9.140 -288.385 9.405 ;
        RECT -288.200 9.140 -287.925 9.405 ;
        RECT -278.740 9.140 -278.465 9.405 ;
        RECT -278.280 9.140 -278.005 9.405 ;
        RECT -268.820 9.140 -268.545 9.405 ;
        RECT -268.360 9.140 -268.085 9.405 ;
        RECT -258.900 9.140 -258.625 9.405 ;
        RECT -258.440 9.140 -258.165 9.405 ;
        RECT -248.980 9.140 -248.705 9.405 ;
        RECT -248.520 9.140 -248.245 9.405 ;
        RECT -239.060 9.140 -238.785 9.405 ;
        RECT -238.600 9.140 -238.325 9.405 ;
        RECT -229.140 9.140 -228.865 9.405 ;
        RECT -228.680 9.140 -228.405 9.405 ;
        RECT -219.220 9.140 -218.945 9.405 ;
        RECT -218.760 9.140 -218.485 9.405 ;
        RECT -209.300 9.140 -209.025 9.405 ;
        RECT -208.840 9.140 -208.565 9.405 ;
        RECT -199.380 9.140 -199.105 9.405 ;
        RECT -198.920 9.140 -198.645 9.405 ;
        RECT -189.460 9.140 -189.185 9.405 ;
        RECT -189.000 9.140 -188.725 9.405 ;
        RECT -179.540 9.140 -179.265 9.405 ;
        RECT -179.080 9.140 -178.805 9.405 ;
        RECT -169.620 9.140 -169.345 9.405 ;
        RECT -169.160 9.140 -168.885 9.405 ;
        RECT -159.700 9.140 -159.425 9.405 ;
        RECT -159.240 9.140 -158.965 9.405 ;
        RECT -149.780 9.140 -149.505 9.405 ;
        RECT -149.320 9.140 -149.045 9.405 ;
        RECT -139.860 9.140 -139.585 9.405 ;
        RECT -139.400 9.140 -139.125 9.405 ;
        RECT -129.940 9.140 -129.665 9.405 ;
        RECT -129.480 9.140 -129.205 9.405 ;
        RECT -120.020 9.140 -119.745 9.405 ;
        RECT -119.560 9.140 -119.285 9.405 ;
        RECT -110.100 9.140 -109.825 9.405 ;
        RECT -109.640 9.140 -109.365 9.405 ;
        RECT -100.180 9.140 -99.905 9.405 ;
        RECT -99.720 9.140 -99.445 9.405 ;
        RECT -90.260 9.140 -89.985 9.405 ;
        RECT -89.800 9.140 -89.525 9.405 ;
        RECT -80.340 9.140 -80.065 9.405 ;
        RECT -79.880 9.140 -79.605 9.405 ;
        RECT -70.420 9.140 -70.145 9.405 ;
        RECT -69.960 9.140 -69.685 9.405 ;
        RECT -60.500 9.140 -60.225 9.405 ;
        RECT -60.040 9.140 -59.765 9.405 ;
        RECT -50.580 9.140 -50.305 9.405 ;
        RECT -50.120 9.140 -49.845 9.405 ;
        RECT -40.660 9.140 -40.385 9.405 ;
        RECT -40.200 9.140 -39.925 9.405 ;
        RECT -30.740 9.140 -30.465 9.405 ;
        RECT -30.280 9.140 -30.005 9.405 ;
        RECT -20.820 9.140 -20.545 9.405 ;
        RECT -20.360 9.140 -20.085 9.405 ;
        RECT -10.900 9.140 -10.625 9.405 ;
        RECT -10.440 9.140 -10.165 9.405 ;
        RECT -0.980 9.140 -0.705 9.405 ;
        RECT -0.520 9.140 -0.245 9.405 ;
        RECT 8.940 9.140 9.215 9.405 ;
        RECT 9.400 9.140 9.675 9.405 ;
        RECT 18.860 9.140 19.135 9.405 ;
        RECT 19.320 9.140 19.595 9.405 ;
        RECT -283.700 6.430 -283.425 6.695 ;
        RECT -283.240 6.430 -282.965 6.695 ;
        RECT -273.780 6.430 -273.505 6.695 ;
        RECT -273.320 6.430 -273.045 6.695 ;
        RECT -263.860 6.430 -263.585 6.695 ;
        RECT -263.400 6.430 -263.125 6.695 ;
        RECT -253.940 6.430 -253.665 6.695 ;
        RECT -253.480 6.430 -253.205 6.695 ;
        RECT -244.020 6.430 -243.745 6.695 ;
        RECT -243.560 6.430 -243.285 6.695 ;
        RECT -234.100 6.430 -233.825 6.695 ;
        RECT -233.640 6.430 -233.365 6.695 ;
        RECT -224.180 6.430 -223.905 6.695 ;
        RECT -223.720 6.430 -223.445 6.695 ;
        RECT -214.260 6.430 -213.985 6.695 ;
        RECT -213.800 6.430 -213.525 6.695 ;
        RECT -204.340 6.430 -204.065 6.695 ;
        RECT -203.880 6.430 -203.605 6.695 ;
        RECT -194.420 6.430 -194.145 6.695 ;
        RECT -193.960 6.430 -193.685 6.695 ;
        RECT -184.500 6.430 -184.225 6.695 ;
        RECT -184.040 6.430 -183.765 6.695 ;
        RECT -174.580 6.430 -174.305 6.695 ;
        RECT -174.120 6.430 -173.845 6.695 ;
        RECT -164.660 6.430 -164.385 6.695 ;
        RECT -164.200 6.430 -163.925 6.695 ;
        RECT -154.740 6.430 -154.465 6.695 ;
        RECT -154.280 6.430 -154.005 6.695 ;
        RECT -144.820 6.430 -144.545 6.695 ;
        RECT -144.360 6.430 -144.085 6.695 ;
        RECT -134.900 6.430 -134.625 6.695 ;
        RECT -134.440 6.430 -134.165 6.695 ;
        RECT -124.980 6.430 -124.705 6.695 ;
        RECT -124.520 6.430 -124.245 6.695 ;
        RECT -115.060 6.430 -114.785 6.695 ;
        RECT -114.600 6.430 -114.325 6.695 ;
        RECT -105.140 6.430 -104.865 6.695 ;
        RECT -104.680 6.430 -104.405 6.695 ;
        RECT -95.220 6.430 -94.945 6.695 ;
        RECT -94.760 6.430 -94.485 6.695 ;
        RECT -85.300 6.430 -85.025 6.695 ;
        RECT -84.840 6.430 -84.565 6.695 ;
        RECT -75.380 6.430 -75.105 6.695 ;
        RECT -74.920 6.430 -74.645 6.695 ;
        RECT -65.460 6.430 -65.185 6.695 ;
        RECT -65.000 6.430 -64.725 6.695 ;
        RECT -55.540 6.430 -55.265 6.695 ;
        RECT -55.080 6.430 -54.805 6.695 ;
        RECT -45.620 6.430 -45.345 6.695 ;
        RECT -45.160 6.430 -44.885 6.695 ;
        RECT -35.700 6.430 -35.425 6.695 ;
        RECT -35.240 6.430 -34.965 6.695 ;
        RECT -25.780 6.430 -25.505 6.695 ;
        RECT -25.320 6.430 -25.045 6.695 ;
        RECT -15.860 6.430 -15.585 6.695 ;
        RECT -15.400 6.430 -15.125 6.695 ;
        RECT -5.940 6.430 -5.665 6.695 ;
        RECT -5.480 6.430 -5.205 6.695 ;
        RECT 3.980 6.430 4.255 6.695 ;
        RECT 4.440 6.430 4.715 6.695 ;
        RECT 13.900 6.430 14.175 6.695 ;
        RECT 14.360 6.430 14.635 6.695 ;
        RECT 23.820 6.430 24.095 6.695 ;
        RECT -288.890 4.840 -288.615 5.105 ;
        RECT -287.960 4.840 -287.685 5.105 ;
        RECT -278.970 4.840 -278.695 5.105 ;
        RECT -278.040 4.840 -277.765 5.105 ;
        RECT -269.050 4.840 -268.775 5.105 ;
        RECT -268.120 4.840 -267.845 5.105 ;
        RECT -259.130 4.840 -258.855 5.105 ;
        RECT -258.200 4.840 -257.925 5.105 ;
        RECT -249.210 4.840 -248.935 5.105 ;
        RECT -248.280 4.840 -248.005 5.105 ;
        RECT -239.290 4.840 -239.015 5.105 ;
        RECT -238.360 4.840 -238.085 5.105 ;
        RECT -229.370 4.840 -229.095 5.105 ;
        RECT -228.440 4.840 -228.165 5.105 ;
        RECT -219.450 4.840 -219.175 5.105 ;
        RECT -218.520 4.840 -218.245 5.105 ;
        RECT -209.530 4.840 -209.255 5.105 ;
        RECT -208.600 4.840 -208.325 5.105 ;
        RECT -199.610 4.840 -199.335 5.105 ;
        RECT -198.680 4.840 -198.405 5.105 ;
        RECT -189.690 4.840 -189.415 5.105 ;
        RECT -188.760 4.840 -188.485 5.105 ;
        RECT -179.770 4.840 -179.495 5.105 ;
        RECT -178.840 4.840 -178.565 5.105 ;
        RECT -169.850 4.840 -169.575 5.105 ;
        RECT -168.920 4.840 -168.645 5.105 ;
        RECT -159.930 4.840 -159.655 5.105 ;
        RECT -159.000 4.840 -158.725 5.105 ;
        RECT -150.010 4.840 -149.735 5.105 ;
        RECT -149.080 4.840 -148.805 5.105 ;
        RECT -140.090 4.840 -139.815 5.105 ;
        RECT -139.160 4.840 -138.885 5.105 ;
        RECT -130.170 4.840 -129.895 5.105 ;
        RECT -129.240 4.840 -128.965 5.105 ;
        RECT -120.250 4.840 -119.975 5.105 ;
        RECT -119.320 4.840 -119.045 5.105 ;
        RECT -110.330 4.840 -110.055 5.105 ;
        RECT -109.400 4.840 -109.125 5.105 ;
        RECT -100.410 4.840 -100.135 5.105 ;
        RECT -99.480 4.840 -99.205 5.105 ;
        RECT -90.490 4.840 -90.215 5.105 ;
        RECT -89.560 4.840 -89.285 5.105 ;
        RECT -80.570 4.840 -80.295 5.105 ;
        RECT -79.640 4.840 -79.365 5.105 ;
        RECT -70.650 4.840 -70.375 5.105 ;
        RECT -69.720 4.840 -69.445 5.105 ;
        RECT -60.730 4.840 -60.455 5.105 ;
        RECT -59.800 4.840 -59.525 5.105 ;
        RECT -50.810 4.840 -50.535 5.105 ;
        RECT -49.880 4.840 -49.605 5.105 ;
        RECT -40.890 4.840 -40.615 5.105 ;
        RECT -39.960 4.840 -39.685 5.105 ;
        RECT -30.970 4.840 -30.695 5.105 ;
        RECT -30.040 4.840 -29.765 5.105 ;
        RECT -21.050 4.840 -20.775 5.105 ;
        RECT -20.120 4.840 -19.845 5.105 ;
        RECT -11.130 4.840 -10.855 5.105 ;
        RECT -10.200 4.840 -9.925 5.105 ;
        RECT -1.210 4.840 -0.935 5.105 ;
        RECT -0.280 4.840 -0.005 5.105 ;
        RECT 8.710 4.840 8.985 5.105 ;
        RECT 9.640 4.840 9.915 5.105 ;
        RECT 18.630 4.840 18.905 5.105 ;
        RECT 19.560 4.840 19.835 5.105 ;
        RECT -283.580 -78.220 -283.305 -77.955 ;
        RECT -282.640 -78.230 -282.365 -77.965 ;
        RECT -272.950 -77.965 -272.680 -77.960 ;
        RECT -272.950 -78.230 -272.445 -77.965 ;
        RECT -263.740 -78.220 -263.465 -77.955 ;
        RECT -262.800 -78.230 -262.525 -77.965 ;
        RECT -253.820 -78.220 -253.545 -77.955 ;
        RECT -252.880 -78.230 -252.605 -77.965 ;
        RECT -243.900 -78.220 -243.625 -77.955 ;
        RECT -242.960 -78.230 -242.685 -77.965 ;
        RECT -233.980 -78.220 -233.705 -77.955 ;
        RECT -233.040 -78.230 -232.765 -77.965 ;
        RECT -224.060 -78.220 -223.785 -77.955 ;
        RECT -223.120 -78.230 -222.845 -77.965 ;
        RECT -214.140 -78.220 -213.865 -77.955 ;
        RECT -213.200 -78.230 -212.925 -77.965 ;
        RECT -204.220 -78.220 -203.945 -77.955 ;
        RECT -203.280 -78.230 -203.005 -77.965 ;
        RECT -194.300 -78.220 -194.025 -77.955 ;
        RECT -193.360 -78.230 -193.085 -77.965 ;
        RECT -184.380 -78.220 -184.105 -77.955 ;
        RECT -183.440 -78.230 -183.165 -77.965 ;
        RECT -174.460 -78.220 -174.185 -77.955 ;
        RECT -173.520 -78.230 -173.245 -77.965 ;
        RECT -164.540 -78.220 -164.265 -77.955 ;
        RECT -163.600 -78.230 -163.325 -77.965 ;
        RECT -154.620 -78.220 -154.345 -77.955 ;
        RECT -153.680 -78.230 -153.405 -77.965 ;
        RECT -144.700 -78.220 -144.425 -77.955 ;
        RECT -143.760 -78.230 -143.485 -77.965 ;
        RECT -134.780 -78.220 -134.505 -77.955 ;
        RECT -133.840 -78.230 -133.565 -77.965 ;
        RECT -124.860 -78.220 -124.585 -77.955 ;
        RECT -123.920 -78.230 -123.645 -77.965 ;
        RECT -114.940 -78.220 -114.665 -77.955 ;
        RECT -114.000 -78.230 -113.725 -77.965 ;
        RECT -105.020 -78.220 -104.745 -77.955 ;
        RECT -104.080 -78.230 -103.805 -77.965 ;
        RECT -95.100 -78.220 -94.825 -77.955 ;
        RECT -94.160 -78.230 -93.885 -77.965 ;
        RECT -85.180 -78.220 -84.905 -77.955 ;
        RECT -84.240 -78.230 -83.965 -77.965 ;
        RECT -75.260 -78.220 -74.985 -77.955 ;
        RECT -74.320 -78.230 -74.045 -77.965 ;
        RECT -65.340 -78.220 -65.065 -77.955 ;
        RECT -64.400 -78.230 -64.125 -77.965 ;
        RECT -55.420 -78.220 -55.145 -77.955 ;
        RECT -54.480 -78.230 -54.205 -77.965 ;
        RECT -45.500 -78.220 -45.225 -77.955 ;
        RECT -44.560 -78.230 -44.285 -77.965 ;
        RECT -35.580 -78.220 -35.305 -77.955 ;
        RECT -34.640 -78.230 -34.365 -77.965 ;
        RECT -25.660 -78.220 -25.385 -77.955 ;
        RECT -24.720 -78.230 -24.445 -77.965 ;
        RECT -15.740 -78.220 -15.465 -77.955 ;
        RECT -14.800 -78.230 -14.525 -77.965 ;
        RECT -5.820 -78.220 -5.545 -77.955 ;
        RECT -4.880 -78.230 -4.605 -77.965 ;
        RECT 4.100 -78.220 4.375 -77.955 ;
        RECT 5.040 -78.230 5.315 -77.965 ;
        RECT 14.020 -78.220 14.295 -77.955 ;
        RECT 14.960 -78.230 15.235 -77.965 ;
        RECT 23.940 -78.220 24.215 -77.955 ;
        RECT -288.300 -79.810 -288.025 -79.545 ;
        RECT -287.840 -79.810 -287.565 -79.545 ;
        RECT -278.380 -79.810 -278.105 -79.545 ;
        RECT -277.920 -79.810 -277.645 -79.545 ;
        RECT -268.460 -79.810 -268.185 -79.545 ;
        RECT -268.000 -79.810 -267.725 -79.545 ;
        RECT -258.540 -79.810 -258.265 -79.545 ;
        RECT -258.080 -79.810 -257.805 -79.545 ;
        RECT -248.620 -79.810 -248.345 -79.545 ;
        RECT -248.160 -79.810 -247.885 -79.545 ;
        RECT -238.700 -79.810 -238.425 -79.545 ;
        RECT -238.240 -79.810 -237.965 -79.545 ;
        RECT -228.780 -79.810 -228.505 -79.545 ;
        RECT -228.320 -79.810 -228.045 -79.545 ;
        RECT -218.860 -79.810 -218.585 -79.545 ;
        RECT -218.400 -79.810 -218.125 -79.545 ;
        RECT -208.940 -79.810 -208.665 -79.545 ;
        RECT -208.480 -79.810 -208.205 -79.545 ;
        RECT -199.020 -79.810 -198.745 -79.545 ;
        RECT -198.560 -79.810 -198.285 -79.545 ;
        RECT -189.100 -79.810 -188.825 -79.545 ;
        RECT -188.640 -79.810 -188.365 -79.545 ;
        RECT -179.180 -79.810 -178.905 -79.545 ;
        RECT -178.720 -79.810 -178.445 -79.545 ;
        RECT -169.260 -79.810 -168.985 -79.545 ;
        RECT -168.800 -79.810 -168.525 -79.545 ;
        RECT -159.340 -79.810 -159.065 -79.545 ;
        RECT -158.880 -79.810 -158.605 -79.545 ;
        RECT -149.420 -79.810 -149.145 -79.545 ;
        RECT -148.960 -79.810 -148.685 -79.545 ;
        RECT -139.500 -79.810 -139.225 -79.545 ;
        RECT -139.040 -79.810 -138.765 -79.545 ;
        RECT -129.580 -79.810 -129.305 -79.545 ;
        RECT -129.120 -79.810 -128.845 -79.545 ;
        RECT -119.660 -79.810 -119.385 -79.545 ;
        RECT -119.200 -79.810 -118.925 -79.545 ;
        RECT -109.740 -79.810 -109.465 -79.545 ;
        RECT -109.280 -79.810 -109.005 -79.545 ;
        RECT -99.820 -79.810 -99.545 -79.545 ;
        RECT -99.360 -79.810 -99.085 -79.545 ;
        RECT -89.900 -79.810 -89.625 -79.545 ;
        RECT -89.440 -79.810 -89.165 -79.545 ;
        RECT -79.980 -79.810 -79.705 -79.545 ;
        RECT -79.520 -79.810 -79.245 -79.545 ;
        RECT -70.060 -79.810 -69.785 -79.545 ;
        RECT -69.600 -79.810 -69.325 -79.545 ;
        RECT -60.140 -79.810 -59.865 -79.545 ;
        RECT -59.680 -79.810 -59.405 -79.545 ;
        RECT -50.220 -79.810 -49.945 -79.545 ;
        RECT -49.760 -79.810 -49.485 -79.545 ;
        RECT -40.300 -79.810 -40.025 -79.545 ;
        RECT -39.840 -79.810 -39.565 -79.545 ;
        RECT -30.380 -79.810 -30.105 -79.545 ;
        RECT -29.920 -79.810 -29.645 -79.545 ;
        RECT -20.460 -79.810 -20.185 -79.545 ;
        RECT -20.000 -79.810 -19.725 -79.545 ;
        RECT -10.540 -79.810 -10.265 -79.545 ;
        RECT -10.080 -79.810 -9.805 -79.545 ;
        RECT -0.620 -79.810 -0.345 -79.545 ;
        RECT -0.160 -79.810 0.115 -79.545 ;
        RECT 9.300 -79.810 9.575 -79.545 ;
        RECT 9.760 -79.810 10.035 -79.545 ;
        RECT 19.220 -79.810 19.495 -79.545 ;
        RECT 19.680 -79.810 19.955 -79.545 ;
        RECT -283.340 -82.520 -283.065 -82.255 ;
        RECT -282.880 -82.520 -282.605 -82.255 ;
        RECT -273.420 -82.520 -273.145 -82.255 ;
        RECT -272.960 -82.520 -272.685 -82.255 ;
        RECT -263.500 -82.520 -263.225 -82.255 ;
        RECT -263.040 -82.520 -262.765 -82.255 ;
        RECT -253.580 -82.520 -253.305 -82.255 ;
        RECT -253.120 -82.520 -252.845 -82.255 ;
        RECT -243.660 -82.520 -243.385 -82.255 ;
        RECT -243.200 -82.520 -242.925 -82.255 ;
        RECT -233.740 -82.520 -233.465 -82.255 ;
        RECT -233.280 -82.520 -233.005 -82.255 ;
        RECT -223.820 -82.520 -223.545 -82.255 ;
        RECT -223.360 -82.520 -223.085 -82.255 ;
        RECT -213.900 -82.520 -213.625 -82.255 ;
        RECT -213.440 -82.520 -213.165 -82.255 ;
        RECT -203.980 -82.520 -203.705 -82.255 ;
        RECT -203.520 -82.520 -203.245 -82.255 ;
        RECT -194.060 -82.520 -193.785 -82.255 ;
        RECT -193.600 -82.520 -193.325 -82.255 ;
        RECT -184.140 -82.520 -183.865 -82.255 ;
        RECT -183.680 -82.520 -183.405 -82.255 ;
        RECT -174.220 -82.520 -173.945 -82.255 ;
        RECT -173.760 -82.520 -173.485 -82.255 ;
        RECT -164.300 -82.520 -164.025 -82.255 ;
        RECT -163.840 -82.520 -163.565 -82.255 ;
        RECT -154.380 -82.520 -154.105 -82.255 ;
        RECT -153.920 -82.520 -153.645 -82.255 ;
        RECT -144.460 -82.520 -144.185 -82.255 ;
        RECT -144.000 -82.520 -143.725 -82.255 ;
        RECT -134.540 -82.520 -134.265 -82.255 ;
        RECT -134.080 -82.520 -133.805 -82.255 ;
        RECT -124.620 -82.520 -124.345 -82.255 ;
        RECT -124.160 -82.520 -123.885 -82.255 ;
        RECT -114.700 -82.520 -114.425 -82.255 ;
        RECT -114.240 -82.520 -113.965 -82.255 ;
        RECT -104.780 -82.520 -104.505 -82.255 ;
        RECT -104.320 -82.520 -104.045 -82.255 ;
        RECT -94.860 -82.520 -94.585 -82.255 ;
        RECT -94.400 -82.520 -94.125 -82.255 ;
        RECT -84.940 -82.520 -84.665 -82.255 ;
        RECT -84.480 -82.520 -84.205 -82.255 ;
        RECT -75.020 -82.520 -74.745 -82.255 ;
        RECT -74.560 -82.520 -74.285 -82.255 ;
        RECT -65.100 -82.520 -64.825 -82.255 ;
        RECT -64.640 -82.520 -64.365 -82.255 ;
        RECT -55.180 -82.520 -54.905 -82.255 ;
        RECT -54.720 -82.520 -54.445 -82.255 ;
        RECT -45.260 -82.520 -44.985 -82.255 ;
        RECT -44.800 -82.520 -44.525 -82.255 ;
        RECT -35.340 -82.520 -35.065 -82.255 ;
        RECT -34.880 -82.520 -34.605 -82.255 ;
        RECT -25.420 -82.520 -25.145 -82.255 ;
        RECT -24.960 -82.520 -24.685 -82.255 ;
        RECT -15.500 -82.520 -15.225 -82.255 ;
        RECT -15.040 -82.520 -14.765 -82.255 ;
        RECT -5.580 -82.520 -5.305 -82.255 ;
        RECT -5.120 -82.520 -4.845 -82.255 ;
        RECT 4.340 -82.520 4.615 -82.255 ;
        RECT 4.800 -82.520 5.075 -82.255 ;
        RECT 14.260 -82.520 14.535 -82.255 ;
        RECT 14.720 -82.520 14.995 -82.255 ;
        RECT 24.180 -82.520 24.455 -82.255 ;
        RECT -288.530 -84.110 -288.255 -83.845 ;
        RECT -287.600 -84.110 -287.325 -83.845 ;
        RECT -278.610 -84.110 -278.335 -83.845 ;
        RECT -277.680 -84.110 -277.405 -83.845 ;
        RECT -268.690 -84.110 -268.415 -83.845 ;
        RECT -267.760 -84.110 -267.485 -83.845 ;
        RECT -258.770 -84.110 -258.495 -83.845 ;
        RECT -257.840 -84.110 -257.565 -83.845 ;
        RECT -248.850 -84.110 -248.575 -83.845 ;
        RECT -247.920 -84.110 -247.645 -83.845 ;
        RECT -238.930 -84.110 -238.655 -83.845 ;
        RECT -238.000 -84.110 -237.725 -83.845 ;
        RECT -229.010 -84.110 -228.735 -83.845 ;
        RECT -228.080 -84.110 -227.805 -83.845 ;
        RECT -219.090 -84.110 -218.815 -83.845 ;
        RECT -218.160 -84.110 -217.885 -83.845 ;
        RECT -209.170 -84.110 -208.895 -83.845 ;
        RECT -208.240 -84.110 -207.965 -83.845 ;
        RECT -199.250 -84.110 -198.975 -83.845 ;
        RECT -198.320 -84.110 -198.045 -83.845 ;
        RECT -189.330 -84.110 -189.055 -83.845 ;
        RECT -188.400 -84.110 -188.125 -83.845 ;
        RECT -179.410 -84.110 -179.135 -83.845 ;
        RECT -178.480 -84.110 -178.205 -83.845 ;
        RECT -169.490 -84.110 -169.215 -83.845 ;
        RECT -168.560 -84.110 -168.285 -83.845 ;
        RECT -159.570 -84.110 -159.295 -83.845 ;
        RECT -158.640 -84.110 -158.365 -83.845 ;
        RECT -149.650 -84.110 -149.375 -83.845 ;
        RECT -148.720 -84.110 -148.445 -83.845 ;
        RECT -139.730 -84.110 -139.455 -83.845 ;
        RECT -138.800 -84.110 -138.525 -83.845 ;
        RECT -129.810 -84.110 -129.535 -83.845 ;
        RECT -128.880 -84.110 -128.605 -83.845 ;
        RECT -119.890 -84.110 -119.615 -83.845 ;
        RECT -118.960 -84.110 -118.685 -83.845 ;
        RECT -109.970 -84.110 -109.695 -83.845 ;
        RECT -109.040 -84.110 -108.765 -83.845 ;
        RECT -100.050 -84.110 -99.775 -83.845 ;
        RECT -99.120 -84.110 -98.845 -83.845 ;
        RECT -90.130 -84.110 -89.855 -83.845 ;
        RECT -89.200 -84.110 -88.925 -83.845 ;
        RECT -80.210 -84.110 -79.935 -83.845 ;
        RECT -79.280 -84.110 -79.005 -83.845 ;
        RECT -70.290 -84.110 -70.015 -83.845 ;
        RECT -69.360 -84.110 -69.085 -83.845 ;
        RECT -60.370 -84.110 -60.095 -83.845 ;
        RECT -59.440 -84.110 -59.165 -83.845 ;
        RECT -50.450 -84.110 -50.175 -83.845 ;
        RECT -49.520 -84.110 -49.245 -83.845 ;
        RECT -40.530 -84.110 -40.255 -83.845 ;
        RECT -39.600 -84.110 -39.325 -83.845 ;
        RECT -30.610 -84.110 -30.335 -83.845 ;
        RECT -29.680 -84.110 -29.405 -83.845 ;
        RECT -20.690 -84.110 -20.415 -83.845 ;
        RECT -19.760 -84.110 -19.485 -83.845 ;
        RECT -10.770 -84.110 -10.495 -83.845 ;
        RECT -9.840 -84.110 -9.565 -83.845 ;
        RECT -0.850 -84.110 -0.575 -83.845 ;
        RECT 0.080 -84.110 0.355 -83.845 ;
        RECT 9.070 -84.110 9.345 -83.845 ;
        RECT 10.000 -84.110 10.275 -83.845 ;
        RECT 18.990 -84.110 19.265 -83.845 ;
        RECT 19.920 -84.110 20.195 -83.845 ;
        RECT -285.340 -172.800 -285.065 -172.535 ;
        RECT -284.400 -172.810 -284.125 -172.545 ;
        RECT -274.710 -172.545 -274.440 -172.540 ;
        RECT -274.710 -172.810 -274.205 -172.545 ;
        RECT -265.500 -172.800 -265.225 -172.535 ;
        RECT -264.560 -172.810 -264.285 -172.545 ;
        RECT -255.580 -172.800 -255.305 -172.535 ;
        RECT -254.640 -172.810 -254.365 -172.545 ;
        RECT -245.660 -172.800 -245.385 -172.535 ;
        RECT -244.720 -172.810 -244.445 -172.545 ;
        RECT -235.740 -172.800 -235.465 -172.535 ;
        RECT -234.800 -172.810 -234.525 -172.545 ;
        RECT -225.820 -172.800 -225.545 -172.535 ;
        RECT -224.880 -172.810 -224.605 -172.545 ;
        RECT -215.900 -172.800 -215.625 -172.535 ;
        RECT -214.960 -172.810 -214.685 -172.545 ;
        RECT -205.980 -172.800 -205.705 -172.535 ;
        RECT -205.040 -172.810 -204.765 -172.545 ;
        RECT -196.060 -172.800 -195.785 -172.535 ;
        RECT -195.120 -172.810 -194.845 -172.545 ;
        RECT -186.140 -172.800 -185.865 -172.535 ;
        RECT -185.200 -172.810 -184.925 -172.545 ;
        RECT -176.220 -172.800 -175.945 -172.535 ;
        RECT -175.280 -172.810 -175.005 -172.545 ;
        RECT -166.300 -172.800 -166.025 -172.535 ;
        RECT -165.360 -172.810 -165.085 -172.545 ;
        RECT -156.380 -172.800 -156.105 -172.535 ;
        RECT -155.440 -172.810 -155.165 -172.545 ;
        RECT -146.460 -172.800 -146.185 -172.535 ;
        RECT -145.520 -172.810 -145.245 -172.545 ;
        RECT -136.540 -172.800 -136.265 -172.535 ;
        RECT -135.600 -172.810 -135.325 -172.545 ;
        RECT -126.620 -172.800 -126.345 -172.535 ;
        RECT -125.680 -172.810 -125.405 -172.545 ;
        RECT -116.700 -172.800 -116.425 -172.535 ;
        RECT -115.760 -172.810 -115.485 -172.545 ;
        RECT -106.780 -172.800 -106.505 -172.535 ;
        RECT -105.840 -172.810 -105.565 -172.545 ;
        RECT -96.860 -172.800 -96.585 -172.535 ;
        RECT -95.920 -172.810 -95.645 -172.545 ;
        RECT -86.940 -172.800 -86.665 -172.535 ;
        RECT -86.000 -172.810 -85.725 -172.545 ;
        RECT -77.020 -172.800 -76.745 -172.535 ;
        RECT -76.080 -172.810 -75.805 -172.545 ;
        RECT -67.100 -172.800 -66.825 -172.535 ;
        RECT -66.160 -172.810 -65.885 -172.545 ;
        RECT -57.180 -172.800 -56.905 -172.535 ;
        RECT -56.240 -172.810 -55.965 -172.545 ;
        RECT -47.260 -172.800 -46.985 -172.535 ;
        RECT -46.320 -172.810 -46.045 -172.545 ;
        RECT -37.340 -172.800 -37.065 -172.535 ;
        RECT -36.400 -172.810 -36.125 -172.545 ;
        RECT -27.420 -172.800 -27.145 -172.535 ;
        RECT -26.480 -172.810 -26.205 -172.545 ;
        RECT -17.500 -172.800 -17.225 -172.535 ;
        RECT -16.560 -172.810 -16.285 -172.545 ;
        RECT -7.580 -172.800 -7.305 -172.535 ;
        RECT -6.640 -172.810 -6.365 -172.545 ;
        RECT 2.340 -172.800 2.615 -172.535 ;
        RECT 3.280 -172.810 3.555 -172.545 ;
        RECT 12.260 -172.800 12.535 -172.535 ;
        RECT 13.200 -172.810 13.475 -172.545 ;
        RECT 22.180 -172.800 22.455 -172.535 ;
        RECT -290.060 -174.390 -289.785 -174.125 ;
        RECT -289.600 -174.390 -289.325 -174.125 ;
        RECT -280.140 -174.390 -279.865 -174.125 ;
        RECT -279.680 -174.390 -279.405 -174.125 ;
        RECT -270.220 -174.390 -269.945 -174.125 ;
        RECT -269.760 -174.390 -269.485 -174.125 ;
        RECT -260.300 -174.390 -260.025 -174.125 ;
        RECT -259.840 -174.390 -259.565 -174.125 ;
        RECT -250.380 -174.390 -250.105 -174.125 ;
        RECT -249.920 -174.390 -249.645 -174.125 ;
        RECT -240.460 -174.390 -240.185 -174.125 ;
        RECT -240.000 -174.390 -239.725 -174.125 ;
        RECT -230.540 -174.390 -230.265 -174.125 ;
        RECT -230.080 -174.390 -229.805 -174.125 ;
        RECT -220.620 -174.390 -220.345 -174.125 ;
        RECT -220.160 -174.390 -219.885 -174.125 ;
        RECT -210.700 -174.390 -210.425 -174.125 ;
        RECT -210.240 -174.390 -209.965 -174.125 ;
        RECT -200.780 -174.390 -200.505 -174.125 ;
        RECT -200.320 -174.390 -200.045 -174.125 ;
        RECT -190.860 -174.390 -190.585 -174.125 ;
        RECT -190.400 -174.390 -190.125 -174.125 ;
        RECT -180.940 -174.390 -180.665 -174.125 ;
        RECT -180.480 -174.390 -180.205 -174.125 ;
        RECT -171.020 -174.390 -170.745 -174.125 ;
        RECT -170.560 -174.390 -170.285 -174.125 ;
        RECT -161.100 -174.390 -160.825 -174.125 ;
        RECT -160.640 -174.390 -160.365 -174.125 ;
        RECT -151.180 -174.390 -150.905 -174.125 ;
        RECT -150.720 -174.390 -150.445 -174.125 ;
        RECT -141.260 -174.390 -140.985 -174.125 ;
        RECT -140.800 -174.390 -140.525 -174.125 ;
        RECT -131.340 -174.390 -131.065 -174.125 ;
        RECT -130.880 -174.390 -130.605 -174.125 ;
        RECT -121.420 -174.390 -121.145 -174.125 ;
        RECT -120.960 -174.390 -120.685 -174.125 ;
        RECT -111.500 -174.390 -111.225 -174.125 ;
        RECT -111.040 -174.390 -110.765 -174.125 ;
        RECT -101.580 -174.390 -101.305 -174.125 ;
        RECT -101.120 -174.390 -100.845 -174.125 ;
        RECT -91.660 -174.390 -91.385 -174.125 ;
        RECT -91.200 -174.390 -90.925 -174.125 ;
        RECT -81.740 -174.390 -81.465 -174.125 ;
        RECT -81.280 -174.390 -81.005 -174.125 ;
        RECT -71.820 -174.390 -71.545 -174.125 ;
        RECT -71.360 -174.390 -71.085 -174.125 ;
        RECT -61.900 -174.390 -61.625 -174.125 ;
        RECT -61.440 -174.390 -61.165 -174.125 ;
        RECT -51.980 -174.390 -51.705 -174.125 ;
        RECT -51.520 -174.390 -51.245 -174.125 ;
        RECT -42.060 -174.390 -41.785 -174.125 ;
        RECT -41.600 -174.390 -41.325 -174.125 ;
        RECT -32.140 -174.390 -31.865 -174.125 ;
        RECT -31.680 -174.390 -31.405 -174.125 ;
        RECT -22.220 -174.390 -21.945 -174.125 ;
        RECT -21.760 -174.390 -21.485 -174.125 ;
        RECT -12.300 -174.390 -12.025 -174.125 ;
        RECT -11.840 -174.390 -11.565 -174.125 ;
        RECT -2.380 -174.390 -2.105 -174.125 ;
        RECT -1.920 -174.390 -1.645 -174.125 ;
        RECT 7.540 -174.390 7.815 -174.125 ;
        RECT 8.000 -174.390 8.275 -174.125 ;
        RECT 17.460 -174.390 17.735 -174.125 ;
        RECT 17.920 -174.390 18.195 -174.125 ;
        RECT -285.100 -177.100 -284.825 -176.835 ;
        RECT -284.640 -177.100 -284.365 -176.835 ;
        RECT -275.180 -177.100 -274.905 -176.835 ;
        RECT -274.720 -177.100 -274.445 -176.835 ;
        RECT -265.260 -177.100 -264.985 -176.835 ;
        RECT -264.800 -177.100 -264.525 -176.835 ;
        RECT -255.340 -177.100 -255.065 -176.835 ;
        RECT -254.880 -177.100 -254.605 -176.835 ;
        RECT -245.420 -177.100 -245.145 -176.835 ;
        RECT -244.960 -177.100 -244.685 -176.835 ;
        RECT -235.500 -177.100 -235.225 -176.835 ;
        RECT -235.040 -177.100 -234.765 -176.835 ;
        RECT -225.580 -177.100 -225.305 -176.835 ;
        RECT -225.120 -177.100 -224.845 -176.835 ;
        RECT -215.660 -177.100 -215.385 -176.835 ;
        RECT -215.200 -177.100 -214.925 -176.835 ;
        RECT -205.740 -177.100 -205.465 -176.835 ;
        RECT -205.280 -177.100 -205.005 -176.835 ;
        RECT -195.820 -177.100 -195.545 -176.835 ;
        RECT -195.360 -177.100 -195.085 -176.835 ;
        RECT -185.900 -177.100 -185.625 -176.835 ;
        RECT -185.440 -177.100 -185.165 -176.835 ;
        RECT -175.980 -177.100 -175.705 -176.835 ;
        RECT -175.520 -177.100 -175.245 -176.835 ;
        RECT -166.060 -177.100 -165.785 -176.835 ;
        RECT -165.600 -177.100 -165.325 -176.835 ;
        RECT -156.140 -177.100 -155.865 -176.835 ;
        RECT -155.680 -177.100 -155.405 -176.835 ;
        RECT -146.220 -177.100 -145.945 -176.835 ;
        RECT -145.760 -177.100 -145.485 -176.835 ;
        RECT -136.300 -177.100 -136.025 -176.835 ;
        RECT -135.840 -177.100 -135.565 -176.835 ;
        RECT -126.380 -177.100 -126.105 -176.835 ;
        RECT -125.920 -177.100 -125.645 -176.835 ;
        RECT -116.460 -177.100 -116.185 -176.835 ;
        RECT -116.000 -177.100 -115.725 -176.835 ;
        RECT -106.540 -177.100 -106.265 -176.835 ;
        RECT -106.080 -177.100 -105.805 -176.835 ;
        RECT -96.620 -177.100 -96.345 -176.835 ;
        RECT -96.160 -177.100 -95.885 -176.835 ;
        RECT -86.700 -177.100 -86.425 -176.835 ;
        RECT -86.240 -177.100 -85.965 -176.835 ;
        RECT -76.780 -177.100 -76.505 -176.835 ;
        RECT -76.320 -177.100 -76.045 -176.835 ;
        RECT -66.860 -177.100 -66.585 -176.835 ;
        RECT -66.400 -177.100 -66.125 -176.835 ;
        RECT -56.940 -177.100 -56.665 -176.835 ;
        RECT -56.480 -177.100 -56.205 -176.835 ;
        RECT -47.020 -177.100 -46.745 -176.835 ;
        RECT -46.560 -177.100 -46.285 -176.835 ;
        RECT -37.100 -177.100 -36.825 -176.835 ;
        RECT -36.640 -177.100 -36.365 -176.835 ;
        RECT -27.180 -177.100 -26.905 -176.835 ;
        RECT -26.720 -177.100 -26.445 -176.835 ;
        RECT -17.260 -177.100 -16.985 -176.835 ;
        RECT -16.800 -177.100 -16.525 -176.835 ;
        RECT -7.340 -177.100 -7.065 -176.835 ;
        RECT -6.880 -177.100 -6.605 -176.835 ;
        RECT 2.580 -177.100 2.855 -176.835 ;
        RECT 3.040 -177.100 3.315 -176.835 ;
        RECT 12.500 -177.100 12.775 -176.835 ;
        RECT 12.960 -177.100 13.235 -176.835 ;
        RECT 22.420 -177.100 22.695 -176.835 ;
        RECT -290.290 -178.690 -290.015 -178.425 ;
        RECT -289.360 -178.690 -289.085 -178.425 ;
        RECT -280.370 -178.690 -280.095 -178.425 ;
        RECT -279.440 -178.690 -279.165 -178.425 ;
        RECT -270.450 -178.690 -270.175 -178.425 ;
        RECT -269.520 -178.690 -269.245 -178.425 ;
        RECT -260.530 -178.690 -260.255 -178.425 ;
        RECT -259.600 -178.690 -259.325 -178.425 ;
        RECT -250.610 -178.690 -250.335 -178.425 ;
        RECT -249.680 -178.690 -249.405 -178.425 ;
        RECT -240.690 -178.690 -240.415 -178.425 ;
        RECT -239.760 -178.690 -239.485 -178.425 ;
        RECT -230.770 -178.690 -230.495 -178.425 ;
        RECT -229.840 -178.690 -229.565 -178.425 ;
        RECT -220.850 -178.690 -220.575 -178.425 ;
        RECT -219.920 -178.690 -219.645 -178.425 ;
        RECT -210.930 -178.690 -210.655 -178.425 ;
        RECT -210.000 -178.690 -209.725 -178.425 ;
        RECT -201.010 -178.690 -200.735 -178.425 ;
        RECT -200.080 -178.690 -199.805 -178.425 ;
        RECT -191.090 -178.690 -190.815 -178.425 ;
        RECT -190.160 -178.690 -189.885 -178.425 ;
        RECT -181.170 -178.690 -180.895 -178.425 ;
        RECT -180.240 -178.690 -179.965 -178.425 ;
        RECT -171.250 -178.690 -170.975 -178.425 ;
        RECT -170.320 -178.690 -170.045 -178.425 ;
        RECT -161.330 -178.690 -161.055 -178.425 ;
        RECT -160.400 -178.690 -160.125 -178.425 ;
        RECT -151.410 -178.690 -151.135 -178.425 ;
        RECT -150.480 -178.690 -150.205 -178.425 ;
        RECT -141.490 -178.690 -141.215 -178.425 ;
        RECT -140.560 -178.690 -140.285 -178.425 ;
        RECT -131.570 -178.690 -131.295 -178.425 ;
        RECT -130.640 -178.690 -130.365 -178.425 ;
        RECT -121.650 -178.690 -121.375 -178.425 ;
        RECT -120.720 -178.690 -120.445 -178.425 ;
        RECT -111.730 -178.690 -111.455 -178.425 ;
        RECT -110.800 -178.690 -110.525 -178.425 ;
        RECT -101.810 -178.690 -101.535 -178.425 ;
        RECT -100.880 -178.690 -100.605 -178.425 ;
        RECT -91.890 -178.690 -91.615 -178.425 ;
        RECT -90.960 -178.690 -90.685 -178.425 ;
        RECT -81.970 -178.690 -81.695 -178.425 ;
        RECT -81.040 -178.690 -80.765 -178.425 ;
        RECT -72.050 -178.690 -71.775 -178.425 ;
        RECT -71.120 -178.690 -70.845 -178.425 ;
        RECT -62.130 -178.690 -61.855 -178.425 ;
        RECT -61.200 -178.690 -60.925 -178.425 ;
        RECT -52.210 -178.690 -51.935 -178.425 ;
        RECT -51.280 -178.690 -51.005 -178.425 ;
        RECT -42.290 -178.690 -42.015 -178.425 ;
        RECT -41.360 -178.690 -41.085 -178.425 ;
        RECT -32.370 -178.690 -32.095 -178.425 ;
        RECT -31.440 -178.690 -31.165 -178.425 ;
        RECT -22.450 -178.690 -22.175 -178.425 ;
        RECT -21.520 -178.690 -21.245 -178.425 ;
        RECT -12.530 -178.690 -12.255 -178.425 ;
        RECT -11.600 -178.690 -11.325 -178.425 ;
        RECT -2.610 -178.690 -2.335 -178.425 ;
        RECT -1.680 -178.690 -1.405 -178.425 ;
        RECT 7.310 -178.690 7.585 -178.425 ;
        RECT 8.240 -178.690 8.515 -178.425 ;
        RECT 17.230 -178.690 17.505 -178.425 ;
        RECT 18.160 -178.690 18.435 -178.425 ;
      LAYER met2 ;
        RECT -282.020 94.730 -280.600 95.140 ;
        RECT -272.100 94.730 -270.680 95.140 ;
        RECT -262.180 94.730 -260.760 95.140 ;
        RECT -252.260 94.730 -250.840 95.140 ;
        RECT -242.340 94.730 -240.920 95.140 ;
        RECT -232.420 94.730 -231.000 95.140 ;
        RECT -222.500 94.730 -221.080 95.140 ;
        RECT -212.580 94.730 -211.160 95.140 ;
        RECT -202.660 94.730 -201.240 95.140 ;
        RECT -192.740 94.730 -191.320 95.140 ;
        RECT -182.820 94.730 -181.400 95.140 ;
        RECT -172.900 94.730 -171.480 95.140 ;
        RECT -162.980 94.730 -161.560 95.140 ;
        RECT -153.060 94.730 -151.640 95.140 ;
        RECT -143.140 94.730 -141.720 95.140 ;
        RECT -133.220 94.730 -131.800 95.140 ;
        RECT -123.300 94.730 -121.880 95.140 ;
        RECT -113.380 94.730 -111.960 95.140 ;
        RECT -103.460 94.730 -102.040 95.140 ;
        RECT -93.540 94.730 -92.120 95.140 ;
        RECT -83.620 94.730 -82.200 95.140 ;
        RECT -73.700 94.730 -72.280 95.140 ;
        RECT -63.780 94.730 -62.360 95.140 ;
        RECT -53.860 94.730 -52.440 95.140 ;
        RECT -43.940 94.730 -42.520 95.140 ;
        RECT -34.020 94.730 -32.600 95.140 ;
        RECT -24.100 94.730 -22.680 95.140 ;
        RECT -14.180 94.730 -12.760 95.140 ;
        RECT -4.260 94.730 -2.840 95.140 ;
        RECT 5.660 94.730 7.080 95.140 ;
        RECT 15.580 94.730 17.000 95.140 ;
        RECT 25.500 94.730 26.440 95.140 ;
        RECT -272.100 94.360 -270.690 94.730 ;
        RECT -286.870 93.090 -285.670 93.570 ;
        RECT -276.950 93.090 -275.750 93.570 ;
        RECT -267.030 93.090 -265.830 93.570 ;
        RECT -257.110 93.090 -255.910 93.570 ;
        RECT -247.190 93.090 -245.990 93.570 ;
        RECT -237.270 93.090 -236.070 93.570 ;
        RECT -227.350 93.090 -226.150 93.570 ;
        RECT -217.430 93.090 -216.230 93.570 ;
        RECT -207.510 93.090 -206.310 93.570 ;
        RECT -197.590 93.090 -196.390 93.570 ;
        RECT -187.670 93.090 -186.470 93.570 ;
        RECT -177.750 93.090 -176.550 93.570 ;
        RECT -167.830 93.090 -166.630 93.570 ;
        RECT -157.910 93.090 -156.710 93.570 ;
        RECT -147.990 93.090 -146.790 93.570 ;
        RECT -138.070 93.090 -136.870 93.570 ;
        RECT -128.150 93.090 -126.950 93.570 ;
        RECT -118.230 93.090 -117.030 93.570 ;
        RECT -108.310 93.090 -107.110 93.570 ;
        RECT -98.390 93.090 -97.190 93.570 ;
        RECT -88.470 93.090 -87.270 93.570 ;
        RECT -78.550 93.090 -77.350 93.570 ;
        RECT -68.630 93.090 -67.430 93.570 ;
        RECT -58.710 93.090 -57.510 93.570 ;
        RECT -48.790 93.090 -47.590 93.570 ;
        RECT -38.870 93.090 -37.670 93.570 ;
        RECT -28.950 93.090 -27.750 93.570 ;
        RECT -19.030 93.090 -17.830 93.570 ;
        RECT -9.110 93.090 -7.910 93.570 ;
        RECT 0.810 93.090 2.010 93.570 ;
        RECT 10.730 93.090 11.930 93.570 ;
        RECT 20.650 93.090 21.850 93.570 ;
        RECT -281.910 90.370 -280.710 90.850 ;
        RECT -271.990 90.370 -270.790 90.850 ;
        RECT -262.070 90.370 -260.870 90.850 ;
        RECT -252.150 90.370 -250.950 90.850 ;
        RECT -242.230 90.370 -241.030 90.850 ;
        RECT -232.310 90.370 -231.110 90.850 ;
        RECT -222.390 90.370 -221.190 90.850 ;
        RECT -212.470 90.370 -211.270 90.850 ;
        RECT -202.550 90.370 -201.350 90.850 ;
        RECT -192.630 90.370 -191.430 90.850 ;
        RECT -182.710 90.370 -181.510 90.850 ;
        RECT -172.790 90.370 -171.590 90.850 ;
        RECT -162.870 90.370 -161.670 90.850 ;
        RECT -152.950 90.370 -151.750 90.850 ;
        RECT -143.030 90.370 -141.830 90.850 ;
        RECT -133.110 90.370 -131.910 90.850 ;
        RECT -123.190 90.370 -121.990 90.850 ;
        RECT -113.270 90.370 -112.070 90.850 ;
        RECT -103.350 90.370 -102.150 90.850 ;
        RECT -93.430 90.370 -92.230 90.850 ;
        RECT -83.510 90.370 -82.310 90.850 ;
        RECT -73.590 90.370 -72.390 90.850 ;
        RECT -63.670 90.370 -62.470 90.850 ;
        RECT -53.750 90.370 -52.550 90.850 ;
        RECT -43.830 90.370 -42.630 90.850 ;
        RECT -33.910 90.370 -32.710 90.850 ;
        RECT -23.990 90.370 -22.790 90.850 ;
        RECT -14.070 90.370 -12.870 90.850 ;
        RECT -4.150 90.370 -2.950 90.850 ;
        RECT 5.770 90.370 6.970 90.850 ;
        RECT 15.690 90.370 16.890 90.850 ;
        RECT 25.610 90.370 26.440 90.850 ;
        RECT -286.980 88.800 -285.560 89.210 ;
        RECT -277.060 88.800 -275.640 89.210 ;
        RECT -267.140 88.800 -265.720 89.210 ;
        RECT -257.220 88.800 -255.800 89.210 ;
        RECT -247.300 88.800 -245.880 89.210 ;
        RECT -237.380 88.800 -235.960 89.210 ;
        RECT -227.460 88.800 -226.040 89.210 ;
        RECT -217.540 88.800 -216.120 89.210 ;
        RECT -207.620 88.800 -206.200 89.210 ;
        RECT -197.700 88.800 -196.280 89.210 ;
        RECT -187.780 88.800 -186.360 89.210 ;
        RECT -177.860 88.800 -176.440 89.210 ;
        RECT -167.940 88.800 -166.520 89.210 ;
        RECT -158.020 88.800 -156.600 89.210 ;
        RECT -148.100 88.800 -146.680 89.210 ;
        RECT -138.180 88.800 -136.760 89.210 ;
        RECT -128.260 88.800 -126.840 89.210 ;
        RECT -118.340 88.800 -116.920 89.210 ;
        RECT -108.420 88.800 -107.000 89.210 ;
        RECT -98.500 88.800 -97.080 89.210 ;
        RECT -88.580 88.800 -87.160 89.210 ;
        RECT -78.660 88.800 -77.240 89.210 ;
        RECT -68.740 88.800 -67.320 89.210 ;
        RECT -58.820 88.800 -57.400 89.210 ;
        RECT -48.900 88.800 -47.480 89.210 ;
        RECT -38.980 88.800 -37.560 89.210 ;
        RECT -29.060 88.800 -27.640 89.210 ;
        RECT -19.140 88.800 -17.720 89.210 ;
        RECT -9.220 88.800 -7.800 89.210 ;
        RECT 0.700 88.800 2.120 89.210 ;
        RECT 10.620 88.800 12.040 89.210 ;
        RECT 20.540 88.800 21.960 89.210 ;
        RECT -284.040 10.680 -282.620 11.090 ;
        RECT -274.120 10.680 -272.700 11.090 ;
        RECT -264.200 10.680 -262.780 11.090 ;
        RECT -254.280 10.680 -252.860 11.090 ;
        RECT -244.360 10.680 -242.940 11.090 ;
        RECT -234.440 10.680 -233.020 11.090 ;
        RECT -224.520 10.680 -223.100 11.090 ;
        RECT -214.600 10.680 -213.180 11.090 ;
        RECT -204.680 10.680 -203.260 11.090 ;
        RECT -194.760 10.680 -193.340 11.090 ;
        RECT -184.840 10.680 -183.420 11.090 ;
        RECT -174.920 10.680 -173.500 11.090 ;
        RECT -165.000 10.680 -163.580 11.090 ;
        RECT -155.080 10.680 -153.660 11.090 ;
        RECT -145.160 10.680 -143.740 11.090 ;
        RECT -135.240 10.680 -133.820 11.090 ;
        RECT -125.320 10.680 -123.900 11.090 ;
        RECT -115.400 10.680 -113.980 11.090 ;
        RECT -105.480 10.680 -104.060 11.090 ;
        RECT -95.560 10.680 -94.140 11.090 ;
        RECT -85.640 10.680 -84.220 11.090 ;
        RECT -75.720 10.680 -74.300 11.090 ;
        RECT -65.800 10.680 -64.380 11.090 ;
        RECT -55.880 10.680 -54.460 11.090 ;
        RECT -45.960 10.680 -44.540 11.090 ;
        RECT -36.040 10.680 -34.620 11.090 ;
        RECT -26.120 10.680 -24.700 11.090 ;
        RECT -16.200 10.680 -14.780 11.090 ;
        RECT -6.280 10.680 -4.860 11.090 ;
        RECT 3.640 10.680 5.060 11.090 ;
        RECT 13.560 10.680 14.980 11.090 ;
        RECT 23.480 10.680 24.420 11.090 ;
        RECT -274.120 10.310 -272.710 10.680 ;
        RECT -288.890 9.040 -287.690 9.520 ;
        RECT -278.970 9.040 -277.770 9.520 ;
        RECT -269.050 9.040 -267.850 9.520 ;
        RECT -259.130 9.040 -257.930 9.520 ;
        RECT -249.210 9.040 -248.010 9.520 ;
        RECT -239.290 9.040 -238.090 9.520 ;
        RECT -229.370 9.040 -228.170 9.520 ;
        RECT -219.450 9.040 -218.250 9.520 ;
        RECT -209.530 9.040 -208.330 9.520 ;
        RECT -199.610 9.040 -198.410 9.520 ;
        RECT -189.690 9.040 -188.490 9.520 ;
        RECT -179.770 9.040 -178.570 9.520 ;
        RECT -169.850 9.040 -168.650 9.520 ;
        RECT -159.930 9.040 -158.730 9.520 ;
        RECT -150.010 9.040 -148.810 9.520 ;
        RECT -140.090 9.040 -138.890 9.520 ;
        RECT -130.170 9.040 -128.970 9.520 ;
        RECT -120.250 9.040 -119.050 9.520 ;
        RECT -110.330 9.040 -109.130 9.520 ;
        RECT -100.410 9.040 -99.210 9.520 ;
        RECT -90.490 9.040 -89.290 9.520 ;
        RECT -80.570 9.040 -79.370 9.520 ;
        RECT -70.650 9.040 -69.450 9.520 ;
        RECT -60.730 9.040 -59.530 9.520 ;
        RECT -50.810 9.040 -49.610 9.520 ;
        RECT -40.890 9.040 -39.690 9.520 ;
        RECT -30.970 9.040 -29.770 9.520 ;
        RECT -21.050 9.040 -19.850 9.520 ;
        RECT -11.130 9.040 -9.930 9.520 ;
        RECT -1.210 9.040 -0.010 9.520 ;
        RECT 8.710 9.040 9.910 9.520 ;
        RECT 18.630 9.040 19.830 9.520 ;
        RECT -283.930 6.320 -282.730 6.800 ;
        RECT -274.010 6.320 -272.810 6.800 ;
        RECT -264.090 6.320 -262.890 6.800 ;
        RECT -254.170 6.320 -252.970 6.800 ;
        RECT -244.250 6.320 -243.050 6.800 ;
        RECT -234.330 6.320 -233.130 6.800 ;
        RECT -224.410 6.320 -223.210 6.800 ;
        RECT -214.490 6.320 -213.290 6.800 ;
        RECT -204.570 6.320 -203.370 6.800 ;
        RECT -194.650 6.320 -193.450 6.800 ;
        RECT -184.730 6.320 -183.530 6.800 ;
        RECT -174.810 6.320 -173.610 6.800 ;
        RECT -164.890 6.320 -163.690 6.800 ;
        RECT -154.970 6.320 -153.770 6.800 ;
        RECT -145.050 6.320 -143.850 6.800 ;
        RECT -135.130 6.320 -133.930 6.800 ;
        RECT -125.210 6.320 -124.010 6.800 ;
        RECT -115.290 6.320 -114.090 6.800 ;
        RECT -105.370 6.320 -104.170 6.800 ;
        RECT -95.450 6.320 -94.250 6.800 ;
        RECT -85.530 6.320 -84.330 6.800 ;
        RECT -75.610 6.320 -74.410 6.800 ;
        RECT -65.690 6.320 -64.490 6.800 ;
        RECT -55.770 6.320 -54.570 6.800 ;
        RECT -45.850 6.320 -44.650 6.800 ;
        RECT -35.930 6.320 -34.730 6.800 ;
        RECT -26.010 6.320 -24.810 6.800 ;
        RECT -16.090 6.320 -14.890 6.800 ;
        RECT -6.170 6.320 -4.970 6.800 ;
        RECT 3.750 6.320 4.950 6.800 ;
        RECT 13.670 6.320 14.870 6.800 ;
        RECT 23.590 6.320 24.420 6.800 ;
        RECT -289.000 4.750 -287.580 5.160 ;
        RECT -279.080 4.750 -277.660 5.160 ;
        RECT -269.160 4.750 -267.740 5.160 ;
        RECT -259.240 4.750 -257.820 5.160 ;
        RECT -249.320 4.750 -247.900 5.160 ;
        RECT -239.400 4.750 -237.980 5.160 ;
        RECT -229.480 4.750 -228.060 5.160 ;
        RECT -219.560 4.750 -218.140 5.160 ;
        RECT -209.640 4.750 -208.220 5.160 ;
        RECT -199.720 4.750 -198.300 5.160 ;
        RECT -189.800 4.750 -188.380 5.160 ;
        RECT -179.880 4.750 -178.460 5.160 ;
        RECT -169.960 4.750 -168.540 5.160 ;
        RECT -160.040 4.750 -158.620 5.160 ;
        RECT -150.120 4.750 -148.700 5.160 ;
        RECT -140.200 4.750 -138.780 5.160 ;
        RECT -130.280 4.750 -128.860 5.160 ;
        RECT -120.360 4.750 -118.940 5.160 ;
        RECT -110.440 4.750 -109.020 5.160 ;
        RECT -100.520 4.750 -99.100 5.160 ;
        RECT -90.600 4.750 -89.180 5.160 ;
        RECT -80.680 4.750 -79.260 5.160 ;
        RECT -70.760 4.750 -69.340 5.160 ;
        RECT -60.840 4.750 -59.420 5.160 ;
        RECT -50.920 4.750 -49.500 5.160 ;
        RECT -41.000 4.750 -39.580 5.160 ;
        RECT -31.080 4.750 -29.660 5.160 ;
        RECT -21.160 4.750 -19.740 5.160 ;
        RECT -11.240 4.750 -9.820 5.160 ;
        RECT -1.320 4.750 0.100 5.160 ;
        RECT 8.600 4.750 10.020 5.160 ;
        RECT 18.520 4.750 19.940 5.160 ;
        RECT -283.680 -78.270 -282.260 -77.860 ;
        RECT -273.760 -78.270 -272.340 -77.860 ;
        RECT -263.840 -78.270 -262.420 -77.860 ;
        RECT -253.920 -78.270 -252.500 -77.860 ;
        RECT -244.000 -78.270 -242.580 -77.860 ;
        RECT -234.080 -78.270 -232.660 -77.860 ;
        RECT -224.160 -78.270 -222.740 -77.860 ;
        RECT -214.240 -78.270 -212.820 -77.860 ;
        RECT -204.320 -78.270 -202.900 -77.860 ;
        RECT -194.400 -78.270 -192.980 -77.860 ;
        RECT -184.480 -78.270 -183.060 -77.860 ;
        RECT -174.560 -78.270 -173.140 -77.860 ;
        RECT -164.640 -78.270 -163.220 -77.860 ;
        RECT -154.720 -78.270 -153.300 -77.860 ;
        RECT -144.800 -78.270 -143.380 -77.860 ;
        RECT -134.880 -78.270 -133.460 -77.860 ;
        RECT -124.960 -78.270 -123.540 -77.860 ;
        RECT -115.040 -78.270 -113.620 -77.860 ;
        RECT -105.120 -78.270 -103.700 -77.860 ;
        RECT -95.200 -78.270 -93.780 -77.860 ;
        RECT -85.280 -78.270 -83.860 -77.860 ;
        RECT -75.360 -78.270 -73.940 -77.860 ;
        RECT -65.440 -78.270 -64.020 -77.860 ;
        RECT -55.520 -78.270 -54.100 -77.860 ;
        RECT -45.600 -78.270 -44.180 -77.860 ;
        RECT -35.680 -78.270 -34.260 -77.860 ;
        RECT -25.760 -78.270 -24.340 -77.860 ;
        RECT -15.840 -78.270 -14.420 -77.860 ;
        RECT -5.920 -78.270 -4.500 -77.860 ;
        RECT 4.000 -78.270 5.420 -77.860 ;
        RECT 13.920 -78.270 15.340 -77.860 ;
        RECT 23.840 -78.270 24.780 -77.860 ;
        RECT -273.760 -78.640 -272.350 -78.270 ;
        RECT -288.530 -79.910 -287.330 -79.430 ;
        RECT -278.610 -79.910 -277.410 -79.430 ;
        RECT -268.690 -79.910 -267.490 -79.430 ;
        RECT -258.770 -79.910 -257.570 -79.430 ;
        RECT -248.850 -79.910 -247.650 -79.430 ;
        RECT -238.930 -79.910 -237.730 -79.430 ;
        RECT -229.010 -79.910 -227.810 -79.430 ;
        RECT -219.090 -79.910 -217.890 -79.430 ;
        RECT -209.170 -79.910 -207.970 -79.430 ;
        RECT -199.250 -79.910 -198.050 -79.430 ;
        RECT -189.330 -79.910 -188.130 -79.430 ;
        RECT -179.410 -79.910 -178.210 -79.430 ;
        RECT -169.490 -79.910 -168.290 -79.430 ;
        RECT -159.570 -79.910 -158.370 -79.430 ;
        RECT -149.650 -79.910 -148.450 -79.430 ;
        RECT -139.730 -79.910 -138.530 -79.430 ;
        RECT -129.810 -79.910 -128.610 -79.430 ;
        RECT -119.890 -79.910 -118.690 -79.430 ;
        RECT -109.970 -79.910 -108.770 -79.430 ;
        RECT -100.050 -79.910 -98.850 -79.430 ;
        RECT -90.130 -79.910 -88.930 -79.430 ;
        RECT -80.210 -79.910 -79.010 -79.430 ;
        RECT -70.290 -79.910 -69.090 -79.430 ;
        RECT -60.370 -79.910 -59.170 -79.430 ;
        RECT -50.450 -79.910 -49.250 -79.430 ;
        RECT -40.530 -79.910 -39.330 -79.430 ;
        RECT -30.610 -79.910 -29.410 -79.430 ;
        RECT -20.690 -79.910 -19.490 -79.430 ;
        RECT -10.770 -79.910 -9.570 -79.430 ;
        RECT -0.850 -79.910 0.350 -79.430 ;
        RECT 9.070 -79.910 10.270 -79.430 ;
        RECT 18.990 -79.910 20.190 -79.430 ;
        RECT -283.570 -82.630 -282.370 -82.150 ;
        RECT -273.650 -82.630 -272.450 -82.150 ;
        RECT -263.730 -82.630 -262.530 -82.150 ;
        RECT -253.810 -82.630 -252.610 -82.150 ;
        RECT -243.890 -82.630 -242.690 -82.150 ;
        RECT -233.970 -82.630 -232.770 -82.150 ;
        RECT -224.050 -82.630 -222.850 -82.150 ;
        RECT -214.130 -82.630 -212.930 -82.150 ;
        RECT -204.210 -82.630 -203.010 -82.150 ;
        RECT -194.290 -82.630 -193.090 -82.150 ;
        RECT -184.370 -82.630 -183.170 -82.150 ;
        RECT -174.450 -82.630 -173.250 -82.150 ;
        RECT -164.530 -82.630 -163.330 -82.150 ;
        RECT -154.610 -82.630 -153.410 -82.150 ;
        RECT -144.690 -82.630 -143.490 -82.150 ;
        RECT -134.770 -82.630 -133.570 -82.150 ;
        RECT -124.850 -82.630 -123.650 -82.150 ;
        RECT -114.930 -82.630 -113.730 -82.150 ;
        RECT -105.010 -82.630 -103.810 -82.150 ;
        RECT -95.090 -82.630 -93.890 -82.150 ;
        RECT -85.170 -82.630 -83.970 -82.150 ;
        RECT -75.250 -82.630 -74.050 -82.150 ;
        RECT -65.330 -82.630 -64.130 -82.150 ;
        RECT -55.410 -82.630 -54.210 -82.150 ;
        RECT -45.490 -82.630 -44.290 -82.150 ;
        RECT -35.570 -82.630 -34.370 -82.150 ;
        RECT -25.650 -82.630 -24.450 -82.150 ;
        RECT -15.730 -82.630 -14.530 -82.150 ;
        RECT -5.810 -82.630 -4.610 -82.150 ;
        RECT 4.110 -82.630 5.310 -82.150 ;
        RECT 14.030 -82.630 15.230 -82.150 ;
        RECT 23.950 -82.630 24.780 -82.150 ;
        RECT -288.640 -84.200 -287.220 -83.790 ;
        RECT -278.720 -84.200 -277.300 -83.790 ;
        RECT -268.800 -84.200 -267.380 -83.790 ;
        RECT -258.880 -84.200 -257.460 -83.790 ;
        RECT -248.960 -84.200 -247.540 -83.790 ;
        RECT -239.040 -84.200 -237.620 -83.790 ;
        RECT -229.120 -84.200 -227.700 -83.790 ;
        RECT -219.200 -84.200 -217.780 -83.790 ;
        RECT -209.280 -84.200 -207.860 -83.790 ;
        RECT -199.360 -84.200 -197.940 -83.790 ;
        RECT -189.440 -84.200 -188.020 -83.790 ;
        RECT -179.520 -84.200 -178.100 -83.790 ;
        RECT -169.600 -84.200 -168.180 -83.790 ;
        RECT -159.680 -84.200 -158.260 -83.790 ;
        RECT -149.760 -84.200 -148.340 -83.790 ;
        RECT -139.840 -84.200 -138.420 -83.790 ;
        RECT -129.920 -84.200 -128.500 -83.790 ;
        RECT -120.000 -84.200 -118.580 -83.790 ;
        RECT -110.080 -84.200 -108.660 -83.790 ;
        RECT -100.160 -84.200 -98.740 -83.790 ;
        RECT -90.240 -84.200 -88.820 -83.790 ;
        RECT -80.320 -84.200 -78.900 -83.790 ;
        RECT -70.400 -84.200 -68.980 -83.790 ;
        RECT -60.480 -84.200 -59.060 -83.790 ;
        RECT -50.560 -84.200 -49.140 -83.790 ;
        RECT -40.640 -84.200 -39.220 -83.790 ;
        RECT -30.720 -84.200 -29.300 -83.790 ;
        RECT -20.800 -84.200 -19.380 -83.790 ;
        RECT -10.880 -84.200 -9.460 -83.790 ;
        RECT -0.960 -84.200 0.460 -83.790 ;
        RECT 8.960 -84.200 10.380 -83.790 ;
        RECT 18.880 -84.200 20.300 -83.790 ;
        RECT -285.440 -172.850 -284.020 -172.440 ;
        RECT -275.520 -172.850 -274.100 -172.440 ;
        RECT -265.600 -172.850 -264.180 -172.440 ;
        RECT -255.680 -172.850 -254.260 -172.440 ;
        RECT -245.760 -172.850 -244.340 -172.440 ;
        RECT -235.840 -172.850 -234.420 -172.440 ;
        RECT -225.920 -172.850 -224.500 -172.440 ;
        RECT -216.000 -172.850 -214.580 -172.440 ;
        RECT -206.080 -172.850 -204.660 -172.440 ;
        RECT -196.160 -172.850 -194.740 -172.440 ;
        RECT -186.240 -172.850 -184.820 -172.440 ;
        RECT -176.320 -172.850 -174.900 -172.440 ;
        RECT -166.400 -172.850 -164.980 -172.440 ;
        RECT -156.480 -172.850 -155.060 -172.440 ;
        RECT -146.560 -172.850 -145.140 -172.440 ;
        RECT -136.640 -172.850 -135.220 -172.440 ;
        RECT -126.720 -172.850 -125.300 -172.440 ;
        RECT -116.800 -172.850 -115.380 -172.440 ;
        RECT -106.880 -172.850 -105.460 -172.440 ;
        RECT -96.960 -172.850 -95.540 -172.440 ;
        RECT -87.040 -172.850 -85.620 -172.440 ;
        RECT -77.120 -172.850 -75.700 -172.440 ;
        RECT -67.200 -172.850 -65.780 -172.440 ;
        RECT -57.280 -172.850 -55.860 -172.440 ;
        RECT -47.360 -172.850 -45.940 -172.440 ;
        RECT -37.440 -172.850 -36.020 -172.440 ;
        RECT -27.520 -172.850 -26.100 -172.440 ;
        RECT -17.600 -172.850 -16.180 -172.440 ;
        RECT -7.680 -172.850 -6.260 -172.440 ;
        RECT 2.240 -172.850 3.660 -172.440 ;
        RECT 12.160 -172.850 13.580 -172.440 ;
        RECT 22.080 -172.850 23.020 -172.440 ;
        RECT -275.520 -173.220 -274.110 -172.850 ;
        RECT -290.290 -174.490 -289.090 -174.010 ;
        RECT -280.370 -174.490 -279.170 -174.010 ;
        RECT -270.450 -174.490 -269.250 -174.010 ;
        RECT -260.530 -174.490 -259.330 -174.010 ;
        RECT -250.610 -174.490 -249.410 -174.010 ;
        RECT -240.690 -174.490 -239.490 -174.010 ;
        RECT -230.770 -174.490 -229.570 -174.010 ;
        RECT -220.850 -174.490 -219.650 -174.010 ;
        RECT -210.930 -174.490 -209.730 -174.010 ;
        RECT -201.010 -174.490 -199.810 -174.010 ;
        RECT -191.090 -174.490 -189.890 -174.010 ;
        RECT -181.170 -174.490 -179.970 -174.010 ;
        RECT -171.250 -174.490 -170.050 -174.010 ;
        RECT -161.330 -174.490 -160.130 -174.010 ;
        RECT -151.410 -174.490 -150.210 -174.010 ;
        RECT -141.490 -174.490 -140.290 -174.010 ;
        RECT -131.570 -174.490 -130.370 -174.010 ;
        RECT -121.650 -174.490 -120.450 -174.010 ;
        RECT -111.730 -174.490 -110.530 -174.010 ;
        RECT -101.810 -174.490 -100.610 -174.010 ;
        RECT -91.890 -174.490 -90.690 -174.010 ;
        RECT -81.970 -174.490 -80.770 -174.010 ;
        RECT -72.050 -174.490 -70.850 -174.010 ;
        RECT -62.130 -174.490 -60.930 -174.010 ;
        RECT -52.210 -174.490 -51.010 -174.010 ;
        RECT -42.290 -174.490 -41.090 -174.010 ;
        RECT -32.370 -174.490 -31.170 -174.010 ;
        RECT -22.450 -174.490 -21.250 -174.010 ;
        RECT -12.530 -174.490 -11.330 -174.010 ;
        RECT -2.610 -174.490 -1.410 -174.010 ;
        RECT 7.310 -174.490 8.510 -174.010 ;
        RECT 17.230 -174.490 18.430 -174.010 ;
        RECT -285.330 -177.210 -284.130 -176.730 ;
        RECT -275.410 -177.210 -274.210 -176.730 ;
        RECT -265.490 -177.210 -264.290 -176.730 ;
        RECT -255.570 -177.210 -254.370 -176.730 ;
        RECT -245.650 -177.210 -244.450 -176.730 ;
        RECT -235.730 -177.210 -234.530 -176.730 ;
        RECT -225.810 -177.210 -224.610 -176.730 ;
        RECT -215.890 -177.210 -214.690 -176.730 ;
        RECT -205.970 -177.210 -204.770 -176.730 ;
        RECT -196.050 -177.210 -194.850 -176.730 ;
        RECT -186.130 -177.210 -184.930 -176.730 ;
        RECT -176.210 -177.210 -175.010 -176.730 ;
        RECT -166.290 -177.210 -165.090 -176.730 ;
        RECT -156.370 -177.210 -155.170 -176.730 ;
        RECT -146.450 -177.210 -145.250 -176.730 ;
        RECT -136.530 -177.210 -135.330 -176.730 ;
        RECT -126.610 -177.210 -125.410 -176.730 ;
        RECT -116.690 -177.210 -115.490 -176.730 ;
        RECT -106.770 -177.210 -105.570 -176.730 ;
        RECT -96.850 -177.210 -95.650 -176.730 ;
        RECT -86.930 -177.210 -85.730 -176.730 ;
        RECT -77.010 -177.210 -75.810 -176.730 ;
        RECT -67.090 -177.210 -65.890 -176.730 ;
        RECT -57.170 -177.210 -55.970 -176.730 ;
        RECT -47.250 -177.210 -46.050 -176.730 ;
        RECT -37.330 -177.210 -36.130 -176.730 ;
        RECT -27.410 -177.210 -26.210 -176.730 ;
        RECT -17.490 -177.210 -16.290 -176.730 ;
        RECT -7.570 -177.210 -6.370 -176.730 ;
        RECT 2.350 -177.210 3.550 -176.730 ;
        RECT 12.270 -177.210 13.470 -176.730 ;
        RECT 22.190 -177.210 23.020 -176.730 ;
        RECT -290.400 -178.780 -288.980 -178.370 ;
        RECT -280.480 -178.780 -279.060 -178.370 ;
        RECT -270.560 -178.780 -269.140 -178.370 ;
        RECT -260.640 -178.780 -259.220 -178.370 ;
        RECT -250.720 -178.780 -249.300 -178.370 ;
        RECT -240.800 -178.780 -239.380 -178.370 ;
        RECT -230.880 -178.780 -229.460 -178.370 ;
        RECT -220.960 -178.780 -219.540 -178.370 ;
        RECT -211.040 -178.780 -209.620 -178.370 ;
        RECT -201.120 -178.780 -199.700 -178.370 ;
        RECT -191.200 -178.780 -189.780 -178.370 ;
        RECT -181.280 -178.780 -179.860 -178.370 ;
        RECT -171.360 -178.780 -169.940 -178.370 ;
        RECT -161.440 -178.780 -160.020 -178.370 ;
        RECT -151.520 -178.780 -150.100 -178.370 ;
        RECT -141.600 -178.780 -140.180 -178.370 ;
        RECT -131.680 -178.780 -130.260 -178.370 ;
        RECT -121.760 -178.780 -120.340 -178.370 ;
        RECT -111.840 -178.780 -110.420 -178.370 ;
        RECT -101.920 -178.780 -100.500 -178.370 ;
        RECT -92.000 -178.780 -90.580 -178.370 ;
        RECT -82.080 -178.780 -80.660 -178.370 ;
        RECT -72.160 -178.780 -70.740 -178.370 ;
        RECT -62.240 -178.780 -60.820 -178.370 ;
        RECT -52.320 -178.780 -50.900 -178.370 ;
        RECT -42.400 -178.780 -40.980 -178.370 ;
        RECT -32.480 -178.780 -31.060 -178.370 ;
        RECT -22.560 -178.780 -21.140 -178.370 ;
        RECT -12.640 -178.780 -11.220 -178.370 ;
        RECT -2.720 -178.780 -1.300 -178.370 ;
        RECT 7.200 -178.780 8.620 -178.370 ;
        RECT 17.120 -178.780 18.540 -178.370 ;
      LAYER via2 ;
        RECT -281.920 94.770 -281.630 95.050 ;
        RECT -280.990 94.760 -280.700 95.040 ;
        RECT -272.000 94.770 -271.710 95.050 ;
        RECT -271.070 94.760 -270.780 95.040 ;
        RECT -262.080 94.770 -261.790 95.050 ;
        RECT -261.150 94.760 -260.860 95.040 ;
        RECT -252.160 94.770 -251.870 95.050 ;
        RECT -251.230 94.760 -250.940 95.040 ;
        RECT -242.240 94.770 -241.950 95.050 ;
        RECT -241.310 94.760 -241.020 95.040 ;
        RECT -232.320 94.770 -232.030 95.050 ;
        RECT -231.390 94.760 -231.100 95.040 ;
        RECT -222.400 94.770 -222.110 95.050 ;
        RECT -221.470 94.760 -221.180 95.040 ;
        RECT -212.480 94.770 -212.190 95.050 ;
        RECT -211.550 94.760 -211.260 95.040 ;
        RECT -202.560 94.770 -202.270 95.050 ;
        RECT -201.630 94.760 -201.340 95.040 ;
        RECT -192.640 94.770 -192.350 95.050 ;
        RECT -191.710 94.760 -191.420 95.040 ;
        RECT -182.720 94.770 -182.430 95.050 ;
        RECT -181.790 94.760 -181.500 95.040 ;
        RECT -172.800 94.770 -172.510 95.050 ;
        RECT -171.870 94.760 -171.580 95.040 ;
        RECT -162.880 94.770 -162.590 95.050 ;
        RECT -161.950 94.760 -161.660 95.040 ;
        RECT -152.960 94.770 -152.670 95.050 ;
        RECT -152.030 94.760 -151.740 95.040 ;
        RECT -143.040 94.770 -142.750 95.050 ;
        RECT -142.110 94.760 -141.820 95.040 ;
        RECT -133.120 94.770 -132.830 95.050 ;
        RECT -132.190 94.760 -131.900 95.040 ;
        RECT -123.200 94.770 -122.910 95.050 ;
        RECT -122.270 94.760 -121.980 95.040 ;
        RECT -113.280 94.770 -112.990 95.050 ;
        RECT -112.350 94.760 -112.060 95.040 ;
        RECT -103.360 94.770 -103.070 95.050 ;
        RECT -102.430 94.760 -102.140 95.040 ;
        RECT -93.440 94.770 -93.150 95.050 ;
        RECT -92.510 94.760 -92.220 95.040 ;
        RECT -83.520 94.770 -83.230 95.050 ;
        RECT -82.590 94.760 -82.300 95.040 ;
        RECT -73.600 94.770 -73.310 95.050 ;
        RECT -72.670 94.760 -72.380 95.040 ;
        RECT -63.680 94.770 -63.390 95.050 ;
        RECT -62.750 94.760 -62.460 95.040 ;
        RECT -53.760 94.770 -53.470 95.050 ;
        RECT -52.830 94.760 -52.540 95.040 ;
        RECT -43.840 94.770 -43.550 95.050 ;
        RECT -42.910 94.760 -42.620 95.040 ;
        RECT -33.920 94.770 -33.630 95.050 ;
        RECT -32.990 94.760 -32.700 95.040 ;
        RECT -24.000 94.770 -23.710 95.050 ;
        RECT -23.070 94.760 -22.780 95.040 ;
        RECT -14.080 94.770 -13.790 95.050 ;
        RECT -13.150 94.760 -12.860 95.040 ;
        RECT -4.160 94.770 -3.870 95.050 ;
        RECT -3.230 94.760 -2.940 95.040 ;
        RECT 5.760 94.770 6.050 95.050 ;
        RECT 6.690 94.760 6.980 95.040 ;
        RECT 15.680 94.770 15.970 95.050 ;
        RECT 16.610 94.760 16.900 95.040 ;
        RECT 25.600 94.770 25.890 95.050 ;
        RECT -286.580 93.280 -286.290 93.560 ;
        RECT -276.660 93.280 -276.370 93.560 ;
        RECT -266.740 93.280 -266.450 93.560 ;
        RECT -256.820 93.280 -256.530 93.560 ;
        RECT -246.900 93.280 -246.610 93.560 ;
        RECT -236.980 93.280 -236.690 93.560 ;
        RECT -227.060 93.280 -226.770 93.560 ;
        RECT -217.140 93.280 -216.850 93.560 ;
        RECT -207.220 93.280 -206.930 93.560 ;
        RECT -197.300 93.280 -197.010 93.560 ;
        RECT -187.380 93.280 -187.090 93.560 ;
        RECT -177.460 93.280 -177.170 93.560 ;
        RECT -167.540 93.280 -167.250 93.560 ;
        RECT -157.620 93.280 -157.330 93.560 ;
        RECT -147.700 93.280 -147.410 93.560 ;
        RECT -137.780 93.280 -137.490 93.560 ;
        RECT -127.860 93.280 -127.570 93.560 ;
        RECT -117.940 93.280 -117.650 93.560 ;
        RECT -108.020 93.280 -107.730 93.560 ;
        RECT -98.100 93.280 -97.810 93.560 ;
        RECT -88.180 93.280 -87.890 93.560 ;
        RECT -78.260 93.280 -77.970 93.560 ;
        RECT -68.340 93.280 -68.050 93.560 ;
        RECT -58.420 93.280 -58.130 93.560 ;
        RECT -48.500 93.280 -48.210 93.560 ;
        RECT -38.580 93.280 -38.290 93.560 ;
        RECT -28.660 93.280 -28.370 93.560 ;
        RECT -18.740 93.280 -18.450 93.560 ;
        RECT -8.820 93.280 -8.530 93.560 ;
        RECT 1.100 93.280 1.390 93.560 ;
        RECT 11.020 93.280 11.310 93.560 ;
        RECT 20.940 93.280 21.230 93.560 ;
        RECT -281.540 90.420 -281.250 90.700 ;
        RECT -271.620 90.420 -271.330 90.700 ;
        RECT -261.700 90.420 -261.410 90.700 ;
        RECT -251.780 90.420 -251.490 90.700 ;
        RECT -241.860 90.420 -241.570 90.700 ;
        RECT -231.940 90.420 -231.650 90.700 ;
        RECT -222.020 90.420 -221.730 90.700 ;
        RECT -212.100 90.420 -211.810 90.700 ;
        RECT -202.180 90.420 -201.890 90.700 ;
        RECT -192.260 90.420 -191.970 90.700 ;
        RECT -182.340 90.420 -182.050 90.700 ;
        RECT -172.420 90.420 -172.130 90.700 ;
        RECT -162.500 90.420 -162.210 90.700 ;
        RECT -152.580 90.420 -152.290 90.700 ;
        RECT -142.660 90.420 -142.370 90.700 ;
        RECT -132.740 90.420 -132.450 90.700 ;
        RECT -122.820 90.420 -122.530 90.700 ;
        RECT -112.900 90.420 -112.610 90.700 ;
        RECT -102.980 90.420 -102.690 90.700 ;
        RECT -93.060 90.420 -92.770 90.700 ;
        RECT -83.140 90.420 -82.850 90.700 ;
        RECT -73.220 90.420 -72.930 90.700 ;
        RECT -63.300 90.420 -63.010 90.700 ;
        RECT -53.380 90.420 -53.090 90.700 ;
        RECT -43.460 90.420 -43.170 90.700 ;
        RECT -33.540 90.420 -33.250 90.700 ;
        RECT -23.620 90.420 -23.330 90.700 ;
        RECT -13.700 90.420 -13.410 90.700 ;
        RECT -3.780 90.420 -3.490 90.700 ;
        RECT 6.140 90.420 6.430 90.700 ;
        RECT 16.060 90.420 16.350 90.700 ;
        RECT 25.980 90.420 26.270 90.700 ;
        RECT -286.880 88.880 -286.590 89.160 ;
        RECT -285.950 88.880 -285.660 89.160 ;
        RECT -276.960 88.880 -276.670 89.160 ;
        RECT -276.030 88.880 -275.740 89.160 ;
        RECT -267.040 88.880 -266.750 89.160 ;
        RECT -266.110 88.880 -265.820 89.160 ;
        RECT -257.120 88.880 -256.830 89.160 ;
        RECT -256.190 88.880 -255.900 89.160 ;
        RECT -247.200 88.880 -246.910 89.160 ;
        RECT -246.270 88.880 -245.980 89.160 ;
        RECT -237.280 88.880 -236.990 89.160 ;
        RECT -236.350 88.880 -236.060 89.160 ;
        RECT -227.360 88.880 -227.070 89.160 ;
        RECT -226.430 88.880 -226.140 89.160 ;
        RECT -217.440 88.880 -217.150 89.160 ;
        RECT -216.510 88.880 -216.220 89.160 ;
        RECT -207.520 88.880 -207.230 89.160 ;
        RECT -206.590 88.880 -206.300 89.160 ;
        RECT -197.600 88.880 -197.310 89.160 ;
        RECT -196.670 88.880 -196.380 89.160 ;
        RECT -187.680 88.880 -187.390 89.160 ;
        RECT -186.750 88.880 -186.460 89.160 ;
        RECT -177.760 88.880 -177.470 89.160 ;
        RECT -176.830 88.880 -176.540 89.160 ;
        RECT -167.840 88.880 -167.550 89.160 ;
        RECT -166.910 88.880 -166.620 89.160 ;
        RECT -157.920 88.880 -157.630 89.160 ;
        RECT -156.990 88.880 -156.700 89.160 ;
        RECT -148.000 88.880 -147.710 89.160 ;
        RECT -147.070 88.880 -146.780 89.160 ;
        RECT -138.080 88.880 -137.790 89.160 ;
        RECT -137.150 88.880 -136.860 89.160 ;
        RECT -128.160 88.880 -127.870 89.160 ;
        RECT -127.230 88.880 -126.940 89.160 ;
        RECT -118.240 88.880 -117.950 89.160 ;
        RECT -117.310 88.880 -117.020 89.160 ;
        RECT -108.320 88.880 -108.030 89.160 ;
        RECT -107.390 88.880 -107.100 89.160 ;
        RECT -98.400 88.880 -98.110 89.160 ;
        RECT -97.470 88.880 -97.180 89.160 ;
        RECT -88.480 88.880 -88.190 89.160 ;
        RECT -87.550 88.880 -87.260 89.160 ;
        RECT -78.560 88.880 -78.270 89.160 ;
        RECT -77.630 88.880 -77.340 89.160 ;
        RECT -68.640 88.880 -68.350 89.160 ;
        RECT -67.710 88.880 -67.420 89.160 ;
        RECT -58.720 88.880 -58.430 89.160 ;
        RECT -57.790 88.880 -57.500 89.160 ;
        RECT -48.800 88.880 -48.510 89.160 ;
        RECT -47.870 88.880 -47.580 89.160 ;
        RECT -38.880 88.880 -38.590 89.160 ;
        RECT -37.950 88.880 -37.660 89.160 ;
        RECT -28.960 88.880 -28.670 89.160 ;
        RECT -28.030 88.880 -27.740 89.160 ;
        RECT -19.040 88.880 -18.750 89.160 ;
        RECT -18.110 88.880 -17.820 89.160 ;
        RECT -9.120 88.880 -8.830 89.160 ;
        RECT -8.190 88.880 -7.900 89.160 ;
        RECT 0.800 88.880 1.090 89.160 ;
        RECT 1.730 88.880 2.020 89.160 ;
        RECT 10.720 88.880 11.010 89.160 ;
        RECT 11.650 88.880 11.940 89.160 ;
        RECT 20.640 88.880 20.930 89.160 ;
        RECT 21.570 88.880 21.860 89.160 ;
        RECT -283.940 10.720 -283.650 11.000 ;
        RECT -283.010 10.710 -282.720 10.990 ;
        RECT -274.020 10.720 -273.730 11.000 ;
        RECT -273.090 10.710 -272.800 10.990 ;
        RECT -264.100 10.720 -263.810 11.000 ;
        RECT -263.170 10.710 -262.880 10.990 ;
        RECT -254.180 10.720 -253.890 11.000 ;
        RECT -253.250 10.710 -252.960 10.990 ;
        RECT -244.260 10.720 -243.970 11.000 ;
        RECT -243.330 10.710 -243.040 10.990 ;
        RECT -234.340 10.720 -234.050 11.000 ;
        RECT -233.410 10.710 -233.120 10.990 ;
        RECT -224.420 10.720 -224.130 11.000 ;
        RECT -223.490 10.710 -223.200 10.990 ;
        RECT -214.500 10.720 -214.210 11.000 ;
        RECT -213.570 10.710 -213.280 10.990 ;
        RECT -204.580 10.720 -204.290 11.000 ;
        RECT -203.650 10.710 -203.360 10.990 ;
        RECT -194.660 10.720 -194.370 11.000 ;
        RECT -193.730 10.710 -193.440 10.990 ;
        RECT -184.740 10.720 -184.450 11.000 ;
        RECT -183.810 10.710 -183.520 10.990 ;
        RECT -174.820 10.720 -174.530 11.000 ;
        RECT -173.890 10.710 -173.600 10.990 ;
        RECT -164.900 10.720 -164.610 11.000 ;
        RECT -163.970 10.710 -163.680 10.990 ;
        RECT -154.980 10.720 -154.690 11.000 ;
        RECT -154.050 10.710 -153.760 10.990 ;
        RECT -145.060 10.720 -144.770 11.000 ;
        RECT -144.130 10.710 -143.840 10.990 ;
        RECT -135.140 10.720 -134.850 11.000 ;
        RECT -134.210 10.710 -133.920 10.990 ;
        RECT -125.220 10.720 -124.930 11.000 ;
        RECT -124.290 10.710 -124.000 10.990 ;
        RECT -115.300 10.720 -115.010 11.000 ;
        RECT -114.370 10.710 -114.080 10.990 ;
        RECT -105.380 10.720 -105.090 11.000 ;
        RECT -104.450 10.710 -104.160 10.990 ;
        RECT -95.460 10.720 -95.170 11.000 ;
        RECT -94.530 10.710 -94.240 10.990 ;
        RECT -85.540 10.720 -85.250 11.000 ;
        RECT -84.610 10.710 -84.320 10.990 ;
        RECT -75.620 10.720 -75.330 11.000 ;
        RECT -74.690 10.710 -74.400 10.990 ;
        RECT -65.700 10.720 -65.410 11.000 ;
        RECT -64.770 10.710 -64.480 10.990 ;
        RECT -55.780 10.720 -55.490 11.000 ;
        RECT -54.850 10.710 -54.560 10.990 ;
        RECT -45.860 10.720 -45.570 11.000 ;
        RECT -44.930 10.710 -44.640 10.990 ;
        RECT -35.940 10.720 -35.650 11.000 ;
        RECT -35.010 10.710 -34.720 10.990 ;
        RECT -26.020 10.720 -25.730 11.000 ;
        RECT -25.090 10.710 -24.800 10.990 ;
        RECT -16.100 10.720 -15.810 11.000 ;
        RECT -15.170 10.710 -14.880 10.990 ;
        RECT -6.180 10.720 -5.890 11.000 ;
        RECT -5.250 10.710 -4.960 10.990 ;
        RECT 3.740 10.720 4.030 11.000 ;
        RECT 4.670 10.710 4.960 10.990 ;
        RECT 13.660 10.720 13.950 11.000 ;
        RECT 14.590 10.710 14.880 10.990 ;
        RECT 23.580 10.720 23.870 11.000 ;
        RECT -288.600 9.230 -288.310 9.510 ;
        RECT -278.680 9.230 -278.390 9.510 ;
        RECT -268.760 9.230 -268.470 9.510 ;
        RECT -258.840 9.230 -258.550 9.510 ;
        RECT -248.920 9.230 -248.630 9.510 ;
        RECT -239.000 9.230 -238.710 9.510 ;
        RECT -229.080 9.230 -228.790 9.510 ;
        RECT -219.160 9.230 -218.870 9.510 ;
        RECT -209.240 9.230 -208.950 9.510 ;
        RECT -199.320 9.230 -199.030 9.510 ;
        RECT -189.400 9.230 -189.110 9.510 ;
        RECT -179.480 9.230 -179.190 9.510 ;
        RECT -169.560 9.230 -169.270 9.510 ;
        RECT -159.640 9.230 -159.350 9.510 ;
        RECT -149.720 9.230 -149.430 9.510 ;
        RECT -139.800 9.230 -139.510 9.510 ;
        RECT -129.880 9.230 -129.590 9.510 ;
        RECT -119.960 9.230 -119.670 9.510 ;
        RECT -110.040 9.230 -109.750 9.510 ;
        RECT -100.120 9.230 -99.830 9.510 ;
        RECT -90.200 9.230 -89.910 9.510 ;
        RECT -80.280 9.230 -79.990 9.510 ;
        RECT -70.360 9.230 -70.070 9.510 ;
        RECT -60.440 9.230 -60.150 9.510 ;
        RECT -50.520 9.230 -50.230 9.510 ;
        RECT -40.600 9.230 -40.310 9.510 ;
        RECT -30.680 9.230 -30.390 9.510 ;
        RECT -20.760 9.230 -20.470 9.510 ;
        RECT -10.840 9.230 -10.550 9.510 ;
        RECT -0.920 9.230 -0.630 9.510 ;
        RECT 9.000 9.230 9.290 9.510 ;
        RECT 18.920 9.230 19.210 9.510 ;
        RECT -283.560 6.370 -283.270 6.650 ;
        RECT -273.640 6.370 -273.350 6.650 ;
        RECT -263.720 6.370 -263.430 6.650 ;
        RECT -253.800 6.370 -253.510 6.650 ;
        RECT -243.880 6.370 -243.590 6.650 ;
        RECT -233.960 6.370 -233.670 6.650 ;
        RECT -224.040 6.370 -223.750 6.650 ;
        RECT -214.120 6.370 -213.830 6.650 ;
        RECT -204.200 6.370 -203.910 6.650 ;
        RECT -194.280 6.370 -193.990 6.650 ;
        RECT -184.360 6.370 -184.070 6.650 ;
        RECT -174.440 6.370 -174.150 6.650 ;
        RECT -164.520 6.370 -164.230 6.650 ;
        RECT -154.600 6.370 -154.310 6.650 ;
        RECT -144.680 6.370 -144.390 6.650 ;
        RECT -134.760 6.370 -134.470 6.650 ;
        RECT -124.840 6.370 -124.550 6.650 ;
        RECT -114.920 6.370 -114.630 6.650 ;
        RECT -105.000 6.370 -104.710 6.650 ;
        RECT -95.080 6.370 -94.790 6.650 ;
        RECT -85.160 6.370 -84.870 6.650 ;
        RECT -75.240 6.370 -74.950 6.650 ;
        RECT -65.320 6.370 -65.030 6.650 ;
        RECT -55.400 6.370 -55.110 6.650 ;
        RECT -45.480 6.370 -45.190 6.650 ;
        RECT -35.560 6.370 -35.270 6.650 ;
        RECT -25.640 6.370 -25.350 6.650 ;
        RECT -15.720 6.370 -15.430 6.650 ;
        RECT -5.800 6.370 -5.510 6.650 ;
        RECT 4.120 6.370 4.410 6.650 ;
        RECT 14.040 6.370 14.330 6.650 ;
        RECT 23.960 6.370 24.250 6.650 ;
        RECT -288.900 4.830 -288.610 5.110 ;
        RECT -287.970 4.830 -287.680 5.110 ;
        RECT -278.980 4.830 -278.690 5.110 ;
        RECT -278.050 4.830 -277.760 5.110 ;
        RECT -269.060 4.830 -268.770 5.110 ;
        RECT -268.130 4.830 -267.840 5.110 ;
        RECT -259.140 4.830 -258.850 5.110 ;
        RECT -258.210 4.830 -257.920 5.110 ;
        RECT -249.220 4.830 -248.930 5.110 ;
        RECT -248.290 4.830 -248.000 5.110 ;
        RECT -239.300 4.830 -239.010 5.110 ;
        RECT -238.370 4.830 -238.080 5.110 ;
        RECT -229.380 4.830 -229.090 5.110 ;
        RECT -228.450 4.830 -228.160 5.110 ;
        RECT -219.460 4.830 -219.170 5.110 ;
        RECT -218.530 4.830 -218.240 5.110 ;
        RECT -209.540 4.830 -209.250 5.110 ;
        RECT -208.610 4.830 -208.320 5.110 ;
        RECT -199.620 4.830 -199.330 5.110 ;
        RECT -198.690 4.830 -198.400 5.110 ;
        RECT -189.700 4.830 -189.410 5.110 ;
        RECT -188.770 4.830 -188.480 5.110 ;
        RECT -179.780 4.830 -179.490 5.110 ;
        RECT -178.850 4.830 -178.560 5.110 ;
        RECT -169.860 4.830 -169.570 5.110 ;
        RECT -168.930 4.830 -168.640 5.110 ;
        RECT -159.940 4.830 -159.650 5.110 ;
        RECT -159.010 4.830 -158.720 5.110 ;
        RECT -150.020 4.830 -149.730 5.110 ;
        RECT -149.090 4.830 -148.800 5.110 ;
        RECT -140.100 4.830 -139.810 5.110 ;
        RECT -139.170 4.830 -138.880 5.110 ;
        RECT -130.180 4.830 -129.890 5.110 ;
        RECT -129.250 4.830 -128.960 5.110 ;
        RECT -120.260 4.830 -119.970 5.110 ;
        RECT -119.330 4.830 -119.040 5.110 ;
        RECT -110.340 4.830 -110.050 5.110 ;
        RECT -109.410 4.830 -109.120 5.110 ;
        RECT -100.420 4.830 -100.130 5.110 ;
        RECT -99.490 4.830 -99.200 5.110 ;
        RECT -90.500 4.830 -90.210 5.110 ;
        RECT -89.570 4.830 -89.280 5.110 ;
        RECT -80.580 4.830 -80.290 5.110 ;
        RECT -79.650 4.830 -79.360 5.110 ;
        RECT -70.660 4.830 -70.370 5.110 ;
        RECT -69.730 4.830 -69.440 5.110 ;
        RECT -60.740 4.830 -60.450 5.110 ;
        RECT -59.810 4.830 -59.520 5.110 ;
        RECT -50.820 4.830 -50.530 5.110 ;
        RECT -49.890 4.830 -49.600 5.110 ;
        RECT -40.900 4.830 -40.610 5.110 ;
        RECT -39.970 4.830 -39.680 5.110 ;
        RECT -30.980 4.830 -30.690 5.110 ;
        RECT -30.050 4.830 -29.760 5.110 ;
        RECT -21.060 4.830 -20.770 5.110 ;
        RECT -20.130 4.830 -19.840 5.110 ;
        RECT -11.140 4.830 -10.850 5.110 ;
        RECT -10.210 4.830 -9.920 5.110 ;
        RECT -1.220 4.830 -0.930 5.110 ;
        RECT -0.290 4.830 0.000 5.110 ;
        RECT 8.700 4.830 8.990 5.110 ;
        RECT 9.630 4.830 9.920 5.110 ;
        RECT 18.620 4.830 18.910 5.110 ;
        RECT 19.550 4.830 19.840 5.110 ;
        RECT -283.580 -78.230 -283.290 -77.950 ;
        RECT -282.650 -78.240 -282.360 -77.960 ;
        RECT -273.660 -78.230 -273.370 -77.950 ;
        RECT -272.730 -78.240 -272.440 -77.960 ;
        RECT -263.740 -78.230 -263.450 -77.950 ;
        RECT -262.810 -78.240 -262.520 -77.960 ;
        RECT -253.820 -78.230 -253.530 -77.950 ;
        RECT -252.890 -78.240 -252.600 -77.960 ;
        RECT -243.900 -78.230 -243.610 -77.950 ;
        RECT -242.970 -78.240 -242.680 -77.960 ;
        RECT -233.980 -78.230 -233.690 -77.950 ;
        RECT -233.050 -78.240 -232.760 -77.960 ;
        RECT -224.060 -78.230 -223.770 -77.950 ;
        RECT -223.130 -78.240 -222.840 -77.960 ;
        RECT -214.140 -78.230 -213.850 -77.950 ;
        RECT -213.210 -78.240 -212.920 -77.960 ;
        RECT -204.220 -78.230 -203.930 -77.950 ;
        RECT -203.290 -78.240 -203.000 -77.960 ;
        RECT -194.300 -78.230 -194.010 -77.950 ;
        RECT -193.370 -78.240 -193.080 -77.960 ;
        RECT -184.380 -78.230 -184.090 -77.950 ;
        RECT -183.450 -78.240 -183.160 -77.960 ;
        RECT -174.460 -78.230 -174.170 -77.950 ;
        RECT -173.530 -78.240 -173.240 -77.960 ;
        RECT -164.540 -78.230 -164.250 -77.950 ;
        RECT -163.610 -78.240 -163.320 -77.960 ;
        RECT -154.620 -78.230 -154.330 -77.950 ;
        RECT -153.690 -78.240 -153.400 -77.960 ;
        RECT -144.700 -78.230 -144.410 -77.950 ;
        RECT -143.770 -78.240 -143.480 -77.960 ;
        RECT -134.780 -78.230 -134.490 -77.950 ;
        RECT -133.850 -78.240 -133.560 -77.960 ;
        RECT -124.860 -78.230 -124.570 -77.950 ;
        RECT -123.930 -78.240 -123.640 -77.960 ;
        RECT -114.940 -78.230 -114.650 -77.950 ;
        RECT -114.010 -78.240 -113.720 -77.960 ;
        RECT -105.020 -78.230 -104.730 -77.950 ;
        RECT -104.090 -78.240 -103.800 -77.960 ;
        RECT -95.100 -78.230 -94.810 -77.950 ;
        RECT -94.170 -78.240 -93.880 -77.960 ;
        RECT -85.180 -78.230 -84.890 -77.950 ;
        RECT -84.250 -78.240 -83.960 -77.960 ;
        RECT -75.260 -78.230 -74.970 -77.950 ;
        RECT -74.330 -78.240 -74.040 -77.960 ;
        RECT -65.340 -78.230 -65.050 -77.950 ;
        RECT -64.410 -78.240 -64.120 -77.960 ;
        RECT -55.420 -78.230 -55.130 -77.950 ;
        RECT -54.490 -78.240 -54.200 -77.960 ;
        RECT -45.500 -78.230 -45.210 -77.950 ;
        RECT -44.570 -78.240 -44.280 -77.960 ;
        RECT -35.580 -78.230 -35.290 -77.950 ;
        RECT -34.650 -78.240 -34.360 -77.960 ;
        RECT -25.660 -78.230 -25.370 -77.950 ;
        RECT -24.730 -78.240 -24.440 -77.960 ;
        RECT -15.740 -78.230 -15.450 -77.950 ;
        RECT -14.810 -78.240 -14.520 -77.960 ;
        RECT -5.820 -78.230 -5.530 -77.950 ;
        RECT -4.890 -78.240 -4.600 -77.960 ;
        RECT 4.100 -78.230 4.390 -77.950 ;
        RECT 5.030 -78.240 5.320 -77.960 ;
        RECT 14.020 -78.230 14.310 -77.950 ;
        RECT 14.950 -78.240 15.240 -77.960 ;
        RECT 23.940 -78.230 24.230 -77.950 ;
        RECT -288.240 -79.720 -287.950 -79.440 ;
        RECT -278.320 -79.720 -278.030 -79.440 ;
        RECT -268.400 -79.720 -268.110 -79.440 ;
        RECT -258.480 -79.720 -258.190 -79.440 ;
        RECT -248.560 -79.720 -248.270 -79.440 ;
        RECT -238.640 -79.720 -238.350 -79.440 ;
        RECT -228.720 -79.720 -228.430 -79.440 ;
        RECT -218.800 -79.720 -218.510 -79.440 ;
        RECT -208.880 -79.720 -208.590 -79.440 ;
        RECT -198.960 -79.720 -198.670 -79.440 ;
        RECT -189.040 -79.720 -188.750 -79.440 ;
        RECT -179.120 -79.720 -178.830 -79.440 ;
        RECT -169.200 -79.720 -168.910 -79.440 ;
        RECT -159.280 -79.720 -158.990 -79.440 ;
        RECT -149.360 -79.720 -149.070 -79.440 ;
        RECT -139.440 -79.720 -139.150 -79.440 ;
        RECT -129.520 -79.720 -129.230 -79.440 ;
        RECT -119.600 -79.720 -119.310 -79.440 ;
        RECT -109.680 -79.720 -109.390 -79.440 ;
        RECT -99.760 -79.720 -99.470 -79.440 ;
        RECT -89.840 -79.720 -89.550 -79.440 ;
        RECT -79.920 -79.720 -79.630 -79.440 ;
        RECT -70.000 -79.720 -69.710 -79.440 ;
        RECT -60.080 -79.720 -59.790 -79.440 ;
        RECT -50.160 -79.720 -49.870 -79.440 ;
        RECT -40.240 -79.720 -39.950 -79.440 ;
        RECT -30.320 -79.720 -30.030 -79.440 ;
        RECT -20.400 -79.720 -20.110 -79.440 ;
        RECT -10.480 -79.720 -10.190 -79.440 ;
        RECT -0.560 -79.720 -0.270 -79.440 ;
        RECT 9.360 -79.720 9.650 -79.440 ;
        RECT 19.280 -79.720 19.570 -79.440 ;
        RECT -283.200 -82.580 -282.910 -82.300 ;
        RECT -273.280 -82.580 -272.990 -82.300 ;
        RECT -263.360 -82.580 -263.070 -82.300 ;
        RECT -253.440 -82.580 -253.150 -82.300 ;
        RECT -243.520 -82.580 -243.230 -82.300 ;
        RECT -233.600 -82.580 -233.310 -82.300 ;
        RECT -223.680 -82.580 -223.390 -82.300 ;
        RECT -213.760 -82.580 -213.470 -82.300 ;
        RECT -203.840 -82.580 -203.550 -82.300 ;
        RECT -193.920 -82.580 -193.630 -82.300 ;
        RECT -184.000 -82.580 -183.710 -82.300 ;
        RECT -174.080 -82.580 -173.790 -82.300 ;
        RECT -164.160 -82.580 -163.870 -82.300 ;
        RECT -154.240 -82.580 -153.950 -82.300 ;
        RECT -144.320 -82.580 -144.030 -82.300 ;
        RECT -134.400 -82.580 -134.110 -82.300 ;
        RECT -124.480 -82.580 -124.190 -82.300 ;
        RECT -114.560 -82.580 -114.270 -82.300 ;
        RECT -104.640 -82.580 -104.350 -82.300 ;
        RECT -94.720 -82.580 -94.430 -82.300 ;
        RECT -84.800 -82.580 -84.510 -82.300 ;
        RECT -74.880 -82.580 -74.590 -82.300 ;
        RECT -64.960 -82.580 -64.670 -82.300 ;
        RECT -55.040 -82.580 -54.750 -82.300 ;
        RECT -45.120 -82.580 -44.830 -82.300 ;
        RECT -35.200 -82.580 -34.910 -82.300 ;
        RECT -25.280 -82.580 -24.990 -82.300 ;
        RECT -15.360 -82.580 -15.070 -82.300 ;
        RECT -5.440 -82.580 -5.150 -82.300 ;
        RECT 4.480 -82.580 4.770 -82.300 ;
        RECT 14.400 -82.580 14.690 -82.300 ;
        RECT 24.320 -82.580 24.610 -82.300 ;
        RECT -288.540 -84.120 -288.250 -83.840 ;
        RECT -287.610 -84.120 -287.320 -83.840 ;
        RECT -278.620 -84.120 -278.330 -83.840 ;
        RECT -277.690 -84.120 -277.400 -83.840 ;
        RECT -268.700 -84.120 -268.410 -83.840 ;
        RECT -267.770 -84.120 -267.480 -83.840 ;
        RECT -258.780 -84.120 -258.490 -83.840 ;
        RECT -257.850 -84.120 -257.560 -83.840 ;
        RECT -248.860 -84.120 -248.570 -83.840 ;
        RECT -247.930 -84.120 -247.640 -83.840 ;
        RECT -238.940 -84.120 -238.650 -83.840 ;
        RECT -238.010 -84.120 -237.720 -83.840 ;
        RECT -229.020 -84.120 -228.730 -83.840 ;
        RECT -228.090 -84.120 -227.800 -83.840 ;
        RECT -219.100 -84.120 -218.810 -83.840 ;
        RECT -218.170 -84.120 -217.880 -83.840 ;
        RECT -209.180 -84.120 -208.890 -83.840 ;
        RECT -208.250 -84.120 -207.960 -83.840 ;
        RECT -199.260 -84.120 -198.970 -83.840 ;
        RECT -198.330 -84.120 -198.040 -83.840 ;
        RECT -189.340 -84.120 -189.050 -83.840 ;
        RECT -188.410 -84.120 -188.120 -83.840 ;
        RECT -179.420 -84.120 -179.130 -83.840 ;
        RECT -178.490 -84.120 -178.200 -83.840 ;
        RECT -169.500 -84.120 -169.210 -83.840 ;
        RECT -168.570 -84.120 -168.280 -83.840 ;
        RECT -159.580 -84.120 -159.290 -83.840 ;
        RECT -158.650 -84.120 -158.360 -83.840 ;
        RECT -149.660 -84.120 -149.370 -83.840 ;
        RECT -148.730 -84.120 -148.440 -83.840 ;
        RECT -139.740 -84.120 -139.450 -83.840 ;
        RECT -138.810 -84.120 -138.520 -83.840 ;
        RECT -129.820 -84.120 -129.530 -83.840 ;
        RECT -128.890 -84.120 -128.600 -83.840 ;
        RECT -119.900 -84.120 -119.610 -83.840 ;
        RECT -118.970 -84.120 -118.680 -83.840 ;
        RECT -109.980 -84.120 -109.690 -83.840 ;
        RECT -109.050 -84.120 -108.760 -83.840 ;
        RECT -100.060 -84.120 -99.770 -83.840 ;
        RECT -99.130 -84.120 -98.840 -83.840 ;
        RECT -90.140 -84.120 -89.850 -83.840 ;
        RECT -89.210 -84.120 -88.920 -83.840 ;
        RECT -80.220 -84.120 -79.930 -83.840 ;
        RECT -79.290 -84.120 -79.000 -83.840 ;
        RECT -70.300 -84.120 -70.010 -83.840 ;
        RECT -69.370 -84.120 -69.080 -83.840 ;
        RECT -60.380 -84.120 -60.090 -83.840 ;
        RECT -59.450 -84.120 -59.160 -83.840 ;
        RECT -50.460 -84.120 -50.170 -83.840 ;
        RECT -49.530 -84.120 -49.240 -83.840 ;
        RECT -40.540 -84.120 -40.250 -83.840 ;
        RECT -39.610 -84.120 -39.320 -83.840 ;
        RECT -30.620 -84.120 -30.330 -83.840 ;
        RECT -29.690 -84.120 -29.400 -83.840 ;
        RECT -20.700 -84.120 -20.410 -83.840 ;
        RECT -19.770 -84.120 -19.480 -83.840 ;
        RECT -10.780 -84.120 -10.490 -83.840 ;
        RECT -9.850 -84.120 -9.560 -83.840 ;
        RECT -0.860 -84.120 -0.570 -83.840 ;
        RECT 0.070 -84.120 0.360 -83.840 ;
        RECT 9.060 -84.120 9.350 -83.840 ;
        RECT 9.990 -84.120 10.280 -83.840 ;
        RECT 18.980 -84.120 19.270 -83.840 ;
        RECT 19.910 -84.120 20.200 -83.840 ;
        RECT -285.340 -172.810 -285.050 -172.530 ;
        RECT -284.410 -172.820 -284.120 -172.540 ;
        RECT -275.420 -172.810 -275.130 -172.530 ;
        RECT -274.490 -172.820 -274.200 -172.540 ;
        RECT -265.500 -172.810 -265.210 -172.530 ;
        RECT -264.570 -172.820 -264.280 -172.540 ;
        RECT -255.580 -172.810 -255.290 -172.530 ;
        RECT -254.650 -172.820 -254.360 -172.540 ;
        RECT -245.660 -172.810 -245.370 -172.530 ;
        RECT -244.730 -172.820 -244.440 -172.540 ;
        RECT -235.740 -172.810 -235.450 -172.530 ;
        RECT -234.810 -172.820 -234.520 -172.540 ;
        RECT -225.820 -172.810 -225.530 -172.530 ;
        RECT -224.890 -172.820 -224.600 -172.540 ;
        RECT -215.900 -172.810 -215.610 -172.530 ;
        RECT -214.970 -172.820 -214.680 -172.540 ;
        RECT -205.980 -172.810 -205.690 -172.530 ;
        RECT -205.050 -172.820 -204.760 -172.540 ;
        RECT -196.060 -172.810 -195.770 -172.530 ;
        RECT -195.130 -172.820 -194.840 -172.540 ;
        RECT -186.140 -172.810 -185.850 -172.530 ;
        RECT -185.210 -172.820 -184.920 -172.540 ;
        RECT -176.220 -172.810 -175.930 -172.530 ;
        RECT -175.290 -172.820 -175.000 -172.540 ;
        RECT -166.300 -172.810 -166.010 -172.530 ;
        RECT -165.370 -172.820 -165.080 -172.540 ;
        RECT -156.380 -172.810 -156.090 -172.530 ;
        RECT -155.450 -172.820 -155.160 -172.540 ;
        RECT -146.460 -172.810 -146.170 -172.530 ;
        RECT -145.530 -172.820 -145.240 -172.540 ;
        RECT -136.540 -172.810 -136.250 -172.530 ;
        RECT -135.610 -172.820 -135.320 -172.540 ;
        RECT -126.620 -172.810 -126.330 -172.530 ;
        RECT -125.690 -172.820 -125.400 -172.540 ;
        RECT -116.700 -172.810 -116.410 -172.530 ;
        RECT -115.770 -172.820 -115.480 -172.540 ;
        RECT -106.780 -172.810 -106.490 -172.530 ;
        RECT -105.850 -172.820 -105.560 -172.540 ;
        RECT -96.860 -172.810 -96.570 -172.530 ;
        RECT -95.930 -172.820 -95.640 -172.540 ;
        RECT -86.940 -172.810 -86.650 -172.530 ;
        RECT -86.010 -172.820 -85.720 -172.540 ;
        RECT -77.020 -172.810 -76.730 -172.530 ;
        RECT -76.090 -172.820 -75.800 -172.540 ;
        RECT -67.100 -172.810 -66.810 -172.530 ;
        RECT -66.170 -172.820 -65.880 -172.540 ;
        RECT -57.180 -172.810 -56.890 -172.530 ;
        RECT -56.250 -172.820 -55.960 -172.540 ;
        RECT -47.260 -172.810 -46.970 -172.530 ;
        RECT -46.330 -172.820 -46.040 -172.540 ;
        RECT -37.340 -172.810 -37.050 -172.530 ;
        RECT -36.410 -172.820 -36.120 -172.540 ;
        RECT -27.420 -172.810 -27.130 -172.530 ;
        RECT -26.490 -172.820 -26.200 -172.540 ;
        RECT -17.500 -172.810 -17.210 -172.530 ;
        RECT -16.570 -172.820 -16.280 -172.540 ;
        RECT -7.580 -172.810 -7.290 -172.530 ;
        RECT -6.650 -172.820 -6.360 -172.540 ;
        RECT 2.340 -172.810 2.630 -172.530 ;
        RECT 3.270 -172.820 3.560 -172.540 ;
        RECT 12.260 -172.810 12.550 -172.530 ;
        RECT 13.190 -172.820 13.480 -172.540 ;
        RECT 22.180 -172.810 22.470 -172.530 ;
        RECT -290.000 -174.300 -289.710 -174.020 ;
        RECT -280.080 -174.300 -279.790 -174.020 ;
        RECT -270.160 -174.300 -269.870 -174.020 ;
        RECT -260.240 -174.300 -259.950 -174.020 ;
        RECT -250.320 -174.300 -250.030 -174.020 ;
        RECT -240.400 -174.300 -240.110 -174.020 ;
        RECT -230.480 -174.300 -230.190 -174.020 ;
        RECT -220.560 -174.300 -220.270 -174.020 ;
        RECT -210.640 -174.300 -210.350 -174.020 ;
        RECT -200.720 -174.300 -200.430 -174.020 ;
        RECT -190.800 -174.300 -190.510 -174.020 ;
        RECT -180.880 -174.300 -180.590 -174.020 ;
        RECT -170.960 -174.300 -170.670 -174.020 ;
        RECT -161.040 -174.300 -160.750 -174.020 ;
        RECT -151.120 -174.300 -150.830 -174.020 ;
        RECT -141.200 -174.300 -140.910 -174.020 ;
        RECT -131.280 -174.300 -130.990 -174.020 ;
        RECT -121.360 -174.300 -121.070 -174.020 ;
        RECT -111.440 -174.300 -111.150 -174.020 ;
        RECT -101.520 -174.300 -101.230 -174.020 ;
        RECT -91.600 -174.300 -91.310 -174.020 ;
        RECT -81.680 -174.300 -81.390 -174.020 ;
        RECT -71.760 -174.300 -71.470 -174.020 ;
        RECT -61.840 -174.300 -61.550 -174.020 ;
        RECT -51.920 -174.300 -51.630 -174.020 ;
        RECT -42.000 -174.300 -41.710 -174.020 ;
        RECT -32.080 -174.300 -31.790 -174.020 ;
        RECT -22.160 -174.300 -21.870 -174.020 ;
        RECT -12.240 -174.300 -11.950 -174.020 ;
        RECT -2.320 -174.300 -2.030 -174.020 ;
        RECT 7.600 -174.300 7.890 -174.020 ;
        RECT 17.520 -174.300 17.810 -174.020 ;
        RECT -284.960 -177.160 -284.670 -176.880 ;
        RECT -275.040 -177.160 -274.750 -176.880 ;
        RECT -265.120 -177.160 -264.830 -176.880 ;
        RECT -255.200 -177.160 -254.910 -176.880 ;
        RECT -245.280 -177.160 -244.990 -176.880 ;
        RECT -235.360 -177.160 -235.070 -176.880 ;
        RECT -225.440 -177.160 -225.150 -176.880 ;
        RECT -215.520 -177.160 -215.230 -176.880 ;
        RECT -205.600 -177.160 -205.310 -176.880 ;
        RECT -195.680 -177.160 -195.390 -176.880 ;
        RECT -185.760 -177.160 -185.470 -176.880 ;
        RECT -175.840 -177.160 -175.550 -176.880 ;
        RECT -165.920 -177.160 -165.630 -176.880 ;
        RECT -156.000 -177.160 -155.710 -176.880 ;
        RECT -146.080 -177.160 -145.790 -176.880 ;
        RECT -136.160 -177.160 -135.870 -176.880 ;
        RECT -126.240 -177.160 -125.950 -176.880 ;
        RECT -116.320 -177.160 -116.030 -176.880 ;
        RECT -106.400 -177.160 -106.110 -176.880 ;
        RECT -96.480 -177.160 -96.190 -176.880 ;
        RECT -86.560 -177.160 -86.270 -176.880 ;
        RECT -76.640 -177.160 -76.350 -176.880 ;
        RECT -66.720 -177.160 -66.430 -176.880 ;
        RECT -56.800 -177.160 -56.510 -176.880 ;
        RECT -46.880 -177.160 -46.590 -176.880 ;
        RECT -36.960 -177.160 -36.670 -176.880 ;
        RECT -27.040 -177.160 -26.750 -176.880 ;
        RECT -17.120 -177.160 -16.830 -176.880 ;
        RECT -7.200 -177.160 -6.910 -176.880 ;
        RECT 2.720 -177.160 3.010 -176.880 ;
        RECT 12.640 -177.160 12.930 -176.880 ;
        RECT 22.560 -177.160 22.850 -176.880 ;
        RECT -290.300 -178.700 -290.010 -178.420 ;
        RECT -289.370 -178.700 -289.080 -178.420 ;
        RECT -280.380 -178.700 -280.090 -178.420 ;
        RECT -279.450 -178.700 -279.160 -178.420 ;
        RECT -270.460 -178.700 -270.170 -178.420 ;
        RECT -269.530 -178.700 -269.240 -178.420 ;
        RECT -260.540 -178.700 -260.250 -178.420 ;
        RECT -259.610 -178.700 -259.320 -178.420 ;
        RECT -250.620 -178.700 -250.330 -178.420 ;
        RECT -249.690 -178.700 -249.400 -178.420 ;
        RECT -240.700 -178.700 -240.410 -178.420 ;
        RECT -239.770 -178.700 -239.480 -178.420 ;
        RECT -230.780 -178.700 -230.490 -178.420 ;
        RECT -229.850 -178.700 -229.560 -178.420 ;
        RECT -220.860 -178.700 -220.570 -178.420 ;
        RECT -219.930 -178.700 -219.640 -178.420 ;
        RECT -210.940 -178.700 -210.650 -178.420 ;
        RECT -210.010 -178.700 -209.720 -178.420 ;
        RECT -201.020 -178.700 -200.730 -178.420 ;
        RECT -200.090 -178.700 -199.800 -178.420 ;
        RECT -191.100 -178.700 -190.810 -178.420 ;
        RECT -190.170 -178.700 -189.880 -178.420 ;
        RECT -181.180 -178.700 -180.890 -178.420 ;
        RECT -180.250 -178.700 -179.960 -178.420 ;
        RECT -171.260 -178.700 -170.970 -178.420 ;
        RECT -170.330 -178.700 -170.040 -178.420 ;
        RECT -161.340 -178.700 -161.050 -178.420 ;
        RECT -160.410 -178.700 -160.120 -178.420 ;
        RECT -151.420 -178.700 -151.130 -178.420 ;
        RECT -150.490 -178.700 -150.200 -178.420 ;
        RECT -141.500 -178.700 -141.210 -178.420 ;
        RECT -140.570 -178.700 -140.280 -178.420 ;
        RECT -131.580 -178.700 -131.290 -178.420 ;
        RECT -130.650 -178.700 -130.360 -178.420 ;
        RECT -121.660 -178.700 -121.370 -178.420 ;
        RECT -120.730 -178.700 -120.440 -178.420 ;
        RECT -111.740 -178.700 -111.450 -178.420 ;
        RECT -110.810 -178.700 -110.520 -178.420 ;
        RECT -101.820 -178.700 -101.530 -178.420 ;
        RECT -100.890 -178.700 -100.600 -178.420 ;
        RECT -91.900 -178.700 -91.610 -178.420 ;
        RECT -90.970 -178.700 -90.680 -178.420 ;
        RECT -81.980 -178.700 -81.690 -178.420 ;
        RECT -81.050 -178.700 -80.760 -178.420 ;
        RECT -72.060 -178.700 -71.770 -178.420 ;
        RECT -71.130 -178.700 -70.840 -178.420 ;
        RECT -62.140 -178.700 -61.850 -178.420 ;
        RECT -61.210 -178.700 -60.920 -178.420 ;
        RECT -52.220 -178.700 -51.930 -178.420 ;
        RECT -51.290 -178.700 -51.000 -178.420 ;
        RECT -42.300 -178.700 -42.010 -178.420 ;
        RECT -41.370 -178.700 -41.080 -178.420 ;
        RECT -32.380 -178.700 -32.090 -178.420 ;
        RECT -31.450 -178.700 -31.160 -178.420 ;
        RECT -22.460 -178.700 -22.170 -178.420 ;
        RECT -21.530 -178.700 -21.240 -178.420 ;
        RECT -12.540 -178.700 -12.250 -178.420 ;
        RECT -11.610 -178.700 -11.320 -178.420 ;
        RECT -2.620 -178.700 -2.330 -178.420 ;
        RECT -1.690 -178.700 -1.400 -178.420 ;
        RECT 7.300 -178.700 7.590 -178.420 ;
        RECT 8.230 -178.700 8.520 -178.420 ;
        RECT 17.220 -178.700 17.510 -178.420 ;
        RECT 18.150 -178.700 18.440 -178.420 ;
      LAYER met3 ;
        RECT -298.750 109.690 -293.660 109.870 ;
        RECT 29.330 109.690 34.420 109.750 ;
        RECT -298.750 100.060 34.420 109.690 ;
        RECT -298.750 82.780 -293.660 100.060 ;
        RECT -291.620 82.780 -290.850 100.060 ;
        RECT -286.660 89.210 -285.890 100.060 ;
        RECT -281.700 95.140 -280.930 100.060 ;
        RECT -282.020 94.730 -280.600 95.140 ;
        RECT -281.700 90.850 -280.930 94.730 ;
        RECT -281.910 90.370 -280.710 90.850 ;
        RECT -286.980 88.800 -285.560 89.210 ;
        RECT -286.660 82.780 -285.890 88.800 ;
        RECT -281.700 82.780 -280.930 90.370 ;
        RECT -276.760 89.210 -275.990 100.060 ;
        RECT -271.780 95.230 -271.010 100.060 ;
        RECT -271.780 95.140 -271.000 95.230 ;
        RECT -272.100 94.730 -270.680 95.140 ;
        RECT -271.780 92.780 -271.000 94.730 ;
        RECT -271.820 90.850 -271.000 92.780 ;
        RECT -271.990 90.370 -270.790 90.850 ;
        RECT -277.060 88.800 -275.640 89.210 ;
        RECT -271.820 88.880 -271.000 90.370 ;
        RECT -266.810 89.210 -266.040 100.060 ;
        RECT -261.820 95.140 -261.050 100.060 ;
        RECT -262.180 94.730 -260.760 95.140 ;
        RECT -261.820 90.850 -261.050 94.730 ;
        RECT -262.070 90.370 -260.870 90.850 ;
        RECT -276.760 82.780 -275.990 88.800 ;
        RECT -271.830 85.270 -271.000 88.880 ;
        RECT -267.140 88.800 -265.720 89.210 ;
        RECT -271.830 82.780 -271.010 85.270 ;
        RECT -266.810 82.780 -266.040 88.800 ;
        RECT -261.820 82.780 -261.050 90.370 ;
        RECT -256.920 89.210 -256.150 100.060 ;
        RECT -251.930 95.140 -251.160 100.060 ;
        RECT -252.260 94.730 -250.840 95.140 ;
        RECT -251.930 90.850 -251.160 94.730 ;
        RECT -252.150 90.370 -250.950 90.850 ;
        RECT -257.220 88.800 -255.800 89.210 ;
        RECT -256.920 82.780 -256.150 88.800 ;
        RECT -251.930 82.780 -251.160 90.370 ;
        RECT -246.990 89.210 -246.220 100.060 ;
        RECT -242.020 95.140 -241.250 100.060 ;
        RECT -242.340 94.730 -240.920 95.140 ;
        RECT -242.020 90.850 -241.250 94.730 ;
        RECT -242.230 90.370 -241.030 90.850 ;
        RECT -247.300 88.800 -245.880 89.210 ;
        RECT -246.990 82.780 -246.220 88.800 ;
        RECT -242.020 82.780 -241.250 90.370 ;
        RECT -237.080 89.210 -236.310 100.060 ;
        RECT -232.120 95.140 -231.350 100.060 ;
        RECT -232.420 94.730 -231.000 95.140 ;
        RECT -232.120 90.850 -231.350 94.730 ;
        RECT -232.310 90.370 -231.110 90.850 ;
        RECT -237.380 88.800 -235.960 89.210 ;
        RECT -237.080 82.780 -236.310 88.800 ;
        RECT -232.120 82.780 -231.350 90.370 ;
        RECT -227.150 89.210 -226.380 100.060 ;
        RECT -222.180 95.140 -221.410 100.060 ;
        RECT -222.500 94.730 -221.080 95.140 ;
        RECT -222.180 90.850 -221.410 94.730 ;
        RECT -222.390 90.370 -221.190 90.850 ;
        RECT -227.460 88.800 -226.040 89.210 ;
        RECT -227.150 82.780 -226.380 88.800 ;
        RECT -222.180 82.780 -221.410 90.370 ;
        RECT -217.200 89.210 -216.430 100.060 ;
        RECT -212.240 95.140 -211.470 100.060 ;
        RECT -212.580 94.730 -211.160 95.140 ;
        RECT -212.240 90.850 -211.470 94.730 ;
        RECT -212.470 90.370 -211.270 90.850 ;
        RECT -217.540 88.800 -216.120 89.210 ;
        RECT -217.200 82.780 -216.430 88.800 ;
        RECT -212.240 82.780 -211.470 90.370 ;
        RECT -207.290 89.210 -206.520 100.060 ;
        RECT -202.350 95.140 -201.580 100.060 ;
        RECT -202.660 94.730 -201.240 95.140 ;
        RECT -202.350 90.850 -201.580 94.730 ;
        RECT -202.550 90.370 -201.350 90.850 ;
        RECT -207.620 88.800 -206.200 89.210 ;
        RECT -207.290 82.780 -206.520 88.800 ;
        RECT -202.350 82.780 -201.580 90.370 ;
        RECT -197.420 89.210 -196.650 100.060 ;
        RECT -192.420 95.140 -191.650 100.060 ;
        RECT -192.740 94.730 -191.320 95.140 ;
        RECT -192.420 90.850 -191.650 94.730 ;
        RECT -192.630 90.370 -191.430 90.850 ;
        RECT -197.700 88.800 -196.280 89.210 ;
        RECT -197.420 82.780 -196.650 88.800 ;
        RECT -192.420 82.780 -191.650 90.370 ;
        RECT -187.460 89.210 -186.690 100.060 ;
        RECT -182.510 95.140 -181.740 100.060 ;
        RECT -182.820 94.730 -181.400 95.140 ;
        RECT -182.510 90.850 -181.740 94.730 ;
        RECT -182.710 90.370 -181.510 90.850 ;
        RECT -187.780 88.800 -186.360 89.210 ;
        RECT -187.460 82.780 -186.690 88.800 ;
        RECT -182.510 82.780 -181.740 90.370 ;
        RECT -177.550 89.210 -176.780 100.060 ;
        RECT -172.560 95.140 -171.790 100.060 ;
        RECT -172.900 94.730 -171.480 95.140 ;
        RECT -172.560 90.850 -171.790 94.730 ;
        RECT -172.790 90.370 -171.590 90.850 ;
        RECT -177.860 88.800 -176.440 89.210 ;
        RECT -177.550 82.780 -176.780 88.800 ;
        RECT -172.560 82.780 -171.790 90.370 ;
        RECT -167.620 89.210 -166.850 100.060 ;
        RECT -162.620 95.140 -161.850 100.060 ;
        RECT -162.980 94.730 -161.560 95.140 ;
        RECT -162.620 90.850 -161.850 94.730 ;
        RECT -162.870 90.370 -161.670 90.850 ;
        RECT -167.940 88.800 -166.520 89.210 ;
        RECT -167.620 82.780 -166.850 88.800 ;
        RECT -162.620 82.780 -161.850 90.370 ;
        RECT -157.710 89.210 -156.940 100.060 ;
        RECT -152.760 95.140 -151.990 100.060 ;
        RECT -153.060 94.730 -151.640 95.140 ;
        RECT -152.760 90.850 -151.990 94.730 ;
        RECT -152.950 90.370 -151.750 90.850 ;
        RECT -158.020 88.800 -156.600 89.210 ;
        RECT -157.710 82.780 -156.940 88.800 ;
        RECT -152.760 82.780 -151.990 90.370 ;
        RECT -147.790 89.210 -147.020 100.060 ;
        RECT -142.830 95.140 -142.060 100.060 ;
        RECT -143.140 94.730 -141.720 95.140 ;
        RECT -142.830 90.850 -142.060 94.730 ;
        RECT -143.030 90.370 -141.830 90.850 ;
        RECT -148.100 88.800 -146.680 89.210 ;
        RECT -147.790 82.780 -147.020 88.800 ;
        RECT -142.830 82.780 -142.060 90.370 ;
        RECT -137.850 89.210 -137.080 100.060 ;
        RECT -132.920 95.140 -132.150 100.060 ;
        RECT -133.220 94.730 -131.800 95.140 ;
        RECT -132.920 90.850 -132.150 94.730 ;
        RECT -133.110 90.370 -131.910 90.850 ;
        RECT -138.180 88.800 -136.760 89.210 ;
        RECT -137.850 82.780 -137.080 88.800 ;
        RECT -132.920 82.780 -132.150 90.370 ;
        RECT -127.940 89.210 -127.170 100.060 ;
        RECT -122.960 95.140 -122.190 100.060 ;
        RECT -123.300 94.730 -121.880 95.140 ;
        RECT -122.960 90.850 -122.190 94.730 ;
        RECT -123.190 90.370 -121.990 90.850 ;
        RECT -128.260 88.800 -126.840 89.210 ;
        RECT -127.940 82.780 -127.170 88.800 ;
        RECT -122.960 82.780 -122.190 90.370 ;
        RECT -118.040 89.210 -117.270 100.060 ;
        RECT -113.080 95.140 -112.310 100.060 ;
        RECT -113.380 94.730 -111.960 95.140 ;
        RECT -113.080 90.850 -112.310 94.730 ;
        RECT -113.270 90.370 -112.070 90.850 ;
        RECT -118.340 88.800 -116.920 89.210 ;
        RECT -118.040 82.780 -117.270 88.800 ;
        RECT -113.080 82.780 -112.310 90.370 ;
        RECT -108.110 89.210 -107.340 100.060 ;
        RECT -103.150 95.140 -102.380 100.060 ;
        RECT -103.460 94.730 -102.040 95.140 ;
        RECT -103.150 90.850 -102.380 94.730 ;
        RECT -103.350 90.370 -102.150 90.850 ;
        RECT -108.420 88.800 -107.000 89.210 ;
        RECT -108.110 82.780 -107.340 88.800 ;
        RECT -103.150 82.780 -102.380 90.370 ;
        RECT -98.160 89.210 -97.390 100.060 ;
        RECT -93.210 95.140 -92.440 100.060 ;
        RECT -93.540 94.730 -92.120 95.140 ;
        RECT -93.210 90.850 -92.440 94.730 ;
        RECT -93.430 90.370 -92.230 90.850 ;
        RECT -98.500 88.800 -97.080 89.210 ;
        RECT -98.160 82.780 -97.390 88.800 ;
        RECT -93.210 82.780 -92.440 90.370 ;
        RECT -88.260 89.210 -87.490 100.060 ;
        RECT -83.270 95.140 -82.500 100.060 ;
        RECT -83.620 94.730 -82.200 95.140 ;
        RECT -83.270 90.850 -82.500 94.730 ;
        RECT -83.510 90.370 -82.310 90.850 ;
        RECT -88.580 88.800 -87.160 89.210 ;
        RECT -88.260 82.780 -87.490 88.800 ;
        RECT -83.270 82.780 -82.500 90.370 ;
        RECT -78.350 89.210 -77.580 100.060 ;
        RECT -73.390 95.140 -72.620 100.060 ;
        RECT -73.700 94.730 -72.280 95.140 ;
        RECT -73.390 90.850 -72.620 94.730 ;
        RECT -73.590 90.370 -72.390 90.850 ;
        RECT -78.660 88.800 -77.240 89.210 ;
        RECT -78.350 82.780 -77.580 88.800 ;
        RECT -73.390 82.780 -72.620 90.370 ;
        RECT -68.410 89.210 -67.640 100.060 ;
        RECT -63.430 95.140 -62.660 100.060 ;
        RECT -63.780 94.730 -62.360 95.140 ;
        RECT -63.430 90.850 -62.660 94.730 ;
        RECT -63.670 90.370 -62.470 90.850 ;
        RECT -68.740 88.800 -67.320 89.210 ;
        RECT -68.410 82.780 -67.640 88.800 ;
        RECT -63.430 82.780 -62.660 90.370 ;
        RECT -58.520 89.210 -57.750 100.060 ;
        RECT -53.520 95.140 -52.750 100.060 ;
        RECT -53.860 94.730 -52.440 95.140 ;
        RECT -53.520 90.850 -52.750 94.730 ;
        RECT -53.750 90.370 -52.550 90.850 ;
        RECT -58.820 88.800 -57.400 89.210 ;
        RECT -58.520 82.780 -57.750 88.800 ;
        RECT -53.520 82.780 -52.750 90.370 ;
        RECT -48.560 89.210 -47.790 100.060 ;
        RECT -43.630 95.140 -42.860 100.060 ;
        RECT -43.940 94.730 -42.520 95.140 ;
        RECT -43.630 90.850 -42.860 94.730 ;
        RECT -43.830 90.370 -42.630 90.850 ;
        RECT -48.900 88.800 -47.480 89.210 ;
        RECT -48.560 82.780 -47.790 88.800 ;
        RECT -43.630 82.780 -42.860 90.370 ;
        RECT -38.680 89.210 -37.910 100.060 ;
        RECT -33.700 95.140 -32.930 100.060 ;
        RECT -34.020 94.730 -32.600 95.140 ;
        RECT -33.700 90.850 -32.930 94.730 ;
        RECT -33.910 90.370 -32.710 90.850 ;
        RECT -38.980 88.800 -37.560 89.210 ;
        RECT -38.680 82.780 -37.910 88.800 ;
        RECT -33.700 82.780 -32.930 90.370 ;
        RECT -28.750 89.210 -27.980 100.060 ;
        RECT -23.800 95.140 -23.030 100.060 ;
        RECT -24.100 94.730 -22.680 95.140 ;
        RECT -23.800 90.850 -23.030 94.730 ;
        RECT -23.990 90.370 -22.790 90.850 ;
        RECT -29.060 88.800 -27.640 89.210 ;
        RECT -28.750 82.780 -27.980 88.800 ;
        RECT -23.800 82.780 -23.030 90.370 ;
        RECT -18.820 89.210 -18.050 100.060 ;
        RECT -13.870 95.140 -13.100 100.060 ;
        RECT -14.180 94.730 -12.760 95.140 ;
        RECT -13.870 90.850 -13.100 94.730 ;
        RECT -14.070 90.370 -12.870 90.850 ;
        RECT -19.140 88.800 -17.720 89.210 ;
        RECT -18.820 82.780 -18.050 88.800 ;
        RECT -13.870 82.780 -13.100 90.370 ;
        RECT -8.920 89.210 -8.150 100.060 ;
        RECT -3.940 95.140 -3.170 100.060 ;
        RECT -4.260 94.730 -2.840 95.140 ;
        RECT -3.940 90.850 -3.170 94.730 ;
        RECT -4.150 90.370 -2.950 90.850 ;
        RECT -9.220 88.800 -7.800 89.210 ;
        RECT -8.920 82.780 -8.150 88.800 ;
        RECT -3.940 82.780 -3.170 90.370 ;
        RECT 1.010 89.210 1.780 100.060 ;
        RECT 5.940 95.140 6.710 100.060 ;
        RECT 5.660 94.730 7.080 95.140 ;
        RECT 5.940 90.850 6.710 94.730 ;
        RECT 5.770 90.370 6.970 90.850 ;
        RECT 0.700 88.800 2.120 89.210 ;
        RECT 1.010 82.780 1.780 88.800 ;
        RECT 5.940 82.780 6.710 90.370 ;
        RECT 10.940 89.210 11.710 100.060 ;
        RECT 15.890 95.140 16.660 100.060 ;
        RECT 15.580 94.730 17.000 95.140 ;
        RECT 15.890 90.850 16.660 94.730 ;
        RECT 15.690 90.370 16.890 90.850 ;
        RECT 10.620 88.800 12.040 89.210 ;
        RECT 10.940 82.780 11.710 88.800 ;
        RECT 15.890 82.780 16.660 90.370 ;
        RECT 20.870 89.210 21.640 100.060 ;
        RECT 25.880 95.140 26.650 100.060 ;
        RECT 25.500 94.730 26.650 95.140 ;
        RECT 25.880 90.850 26.650 94.730 ;
        RECT 25.610 90.370 26.440 90.850 ;
        RECT 20.540 88.800 21.960 89.210 ;
        RECT 20.870 82.780 21.640 88.800 ;
        RECT 25.880 82.780 26.650 90.370 ;
        RECT 29.330 83.200 34.420 100.060 ;
        RECT 27.700 82.780 164.350 83.200 ;
        RECT -298.750 78.340 164.350 82.780 ;
        RECT -317.240 78.330 164.350 78.340 ;
        RECT -335.510 73.570 164.350 78.330 ;
        RECT -335.510 73.150 34.420 73.570 ;
        RECT -335.510 73.140 -293.660 73.150 ;
        RECT -335.510 73.120 -298.380 73.140 ;
        RECT -335.510 73.110 -316.650 73.120 ;
        RECT -300.770 25.640 -295.680 25.820 ;
        RECT -196.490 25.640 -159.330 73.150 ;
        RECT 29.330 73.020 34.420 73.150 ;
        RECT 27.310 25.640 32.400 25.700 ;
        RECT -300.770 16.010 32.400 25.640 ;
        RECT -300.770 -1.270 -295.680 16.010 ;
        RECT -293.640 -1.270 -292.870 16.010 ;
        RECT -288.680 5.160 -287.910 16.010 ;
        RECT -283.720 11.090 -282.950 16.010 ;
        RECT -284.040 10.680 -282.620 11.090 ;
        RECT -283.720 6.800 -282.950 10.680 ;
        RECT -283.930 6.320 -282.730 6.800 ;
        RECT -289.000 4.750 -287.580 5.160 ;
        RECT -288.680 -1.270 -287.910 4.750 ;
        RECT -283.720 -1.270 -282.950 6.320 ;
        RECT -278.780 5.160 -278.010 16.010 ;
        RECT -273.800 11.180 -273.030 16.010 ;
        RECT -273.800 11.090 -273.020 11.180 ;
        RECT -274.120 10.680 -272.700 11.090 ;
        RECT -273.800 8.730 -273.020 10.680 ;
        RECT -273.840 6.800 -273.020 8.730 ;
        RECT -274.010 6.320 -272.810 6.800 ;
        RECT -279.080 4.750 -277.660 5.160 ;
        RECT -273.840 4.830 -273.020 6.320 ;
        RECT -268.830 5.160 -268.060 16.010 ;
        RECT -263.840 11.090 -263.070 16.010 ;
        RECT -264.200 10.680 -262.780 11.090 ;
        RECT -263.840 6.800 -263.070 10.680 ;
        RECT -264.090 6.320 -262.890 6.800 ;
        RECT -278.780 -1.270 -278.010 4.750 ;
        RECT -273.850 1.220 -273.020 4.830 ;
        RECT -269.160 4.750 -267.740 5.160 ;
        RECT -273.850 -1.270 -273.030 1.220 ;
        RECT -268.830 -1.270 -268.060 4.750 ;
        RECT -263.840 -1.270 -263.070 6.320 ;
        RECT -258.940 5.160 -258.170 16.010 ;
        RECT -253.950 11.090 -253.180 16.010 ;
        RECT -254.280 10.680 -252.860 11.090 ;
        RECT -253.950 6.800 -253.180 10.680 ;
        RECT -254.170 6.320 -252.970 6.800 ;
        RECT -259.240 4.750 -257.820 5.160 ;
        RECT -258.940 -1.270 -258.170 4.750 ;
        RECT -253.950 -1.270 -253.180 6.320 ;
        RECT -249.010 5.160 -248.240 16.010 ;
        RECT -244.040 11.090 -243.270 16.010 ;
        RECT -244.360 10.680 -242.940 11.090 ;
        RECT -244.040 6.800 -243.270 10.680 ;
        RECT -244.250 6.320 -243.050 6.800 ;
        RECT -249.320 4.750 -247.900 5.160 ;
        RECT -249.010 -1.270 -248.240 4.750 ;
        RECT -244.040 -1.270 -243.270 6.320 ;
        RECT -239.100 5.160 -238.330 16.010 ;
        RECT -234.140 11.090 -233.370 16.010 ;
        RECT -234.440 10.680 -233.020 11.090 ;
        RECT -234.140 6.800 -233.370 10.680 ;
        RECT -234.330 6.320 -233.130 6.800 ;
        RECT -239.400 4.750 -237.980 5.160 ;
        RECT -239.100 -1.270 -238.330 4.750 ;
        RECT -234.140 -1.270 -233.370 6.320 ;
        RECT -229.170 5.160 -228.400 16.010 ;
        RECT -224.200 11.090 -223.430 16.010 ;
        RECT -224.520 10.680 -223.100 11.090 ;
        RECT -224.200 6.800 -223.430 10.680 ;
        RECT -224.410 6.320 -223.210 6.800 ;
        RECT -229.480 4.750 -228.060 5.160 ;
        RECT -229.170 -1.270 -228.400 4.750 ;
        RECT -224.200 -1.270 -223.430 6.320 ;
        RECT -219.220 5.160 -218.450 16.010 ;
        RECT -214.260 11.090 -213.490 16.010 ;
        RECT -214.600 10.680 -213.180 11.090 ;
        RECT -214.260 6.800 -213.490 10.680 ;
        RECT -214.490 6.320 -213.290 6.800 ;
        RECT -219.560 4.750 -218.140 5.160 ;
        RECT -219.220 -1.270 -218.450 4.750 ;
        RECT -214.260 -1.270 -213.490 6.320 ;
        RECT -209.310 5.160 -208.540 16.010 ;
        RECT -204.370 11.090 -203.600 16.010 ;
        RECT -204.680 10.680 -203.260 11.090 ;
        RECT -204.370 6.800 -203.600 10.680 ;
        RECT -204.570 6.320 -203.370 6.800 ;
        RECT -209.640 4.750 -208.220 5.160 ;
        RECT -209.310 -1.270 -208.540 4.750 ;
        RECT -204.370 -1.270 -203.600 6.320 ;
        RECT -199.440 5.160 -198.670 16.010 ;
        RECT -194.440 11.090 -193.670 16.010 ;
        RECT -194.760 10.680 -193.340 11.090 ;
        RECT -194.440 6.800 -193.670 10.680 ;
        RECT -194.650 6.320 -193.450 6.800 ;
        RECT -199.720 4.750 -198.300 5.160 ;
        RECT -199.440 -1.270 -198.670 4.750 ;
        RECT -194.440 -1.270 -193.670 6.320 ;
        RECT -189.480 5.160 -188.710 16.010 ;
        RECT -184.530 11.090 -183.760 16.010 ;
        RECT -184.840 10.680 -183.420 11.090 ;
        RECT -184.530 6.800 -183.760 10.680 ;
        RECT -184.730 6.320 -183.530 6.800 ;
        RECT -189.800 4.750 -188.380 5.160 ;
        RECT -189.480 -1.270 -188.710 4.750 ;
        RECT -184.530 -1.270 -183.760 6.320 ;
        RECT -179.570 5.160 -178.800 16.010 ;
        RECT -174.580 11.090 -173.810 16.010 ;
        RECT -174.920 10.680 -173.500 11.090 ;
        RECT -174.580 6.800 -173.810 10.680 ;
        RECT -174.810 6.320 -173.610 6.800 ;
        RECT -179.880 4.750 -178.460 5.160 ;
        RECT -179.570 -1.270 -178.800 4.750 ;
        RECT -174.580 -1.270 -173.810 6.320 ;
        RECT -169.640 5.160 -168.870 16.010 ;
        RECT -164.640 11.090 -163.870 16.010 ;
        RECT -165.000 10.680 -163.580 11.090 ;
        RECT -164.640 6.800 -163.870 10.680 ;
        RECT -164.890 6.320 -163.690 6.800 ;
        RECT -169.960 4.750 -168.540 5.160 ;
        RECT -169.640 -1.270 -168.870 4.750 ;
        RECT -164.640 -1.270 -163.870 6.320 ;
        RECT -159.730 5.160 -158.960 16.010 ;
        RECT -154.780 11.090 -154.010 16.010 ;
        RECT -155.080 10.680 -153.660 11.090 ;
        RECT -154.780 6.800 -154.010 10.680 ;
        RECT -154.970 6.320 -153.770 6.800 ;
        RECT -160.040 4.750 -158.620 5.160 ;
        RECT -159.730 -1.270 -158.960 4.750 ;
        RECT -154.780 -1.270 -154.010 6.320 ;
        RECT -149.810 5.160 -149.040 16.010 ;
        RECT -144.850 11.090 -144.080 16.010 ;
        RECT -145.160 10.680 -143.740 11.090 ;
        RECT -144.850 6.800 -144.080 10.680 ;
        RECT -145.050 6.320 -143.850 6.800 ;
        RECT -150.120 4.750 -148.700 5.160 ;
        RECT -149.810 -1.270 -149.040 4.750 ;
        RECT -144.850 -1.270 -144.080 6.320 ;
        RECT -139.870 5.160 -139.100 16.010 ;
        RECT -134.940 11.090 -134.170 16.010 ;
        RECT -135.240 10.680 -133.820 11.090 ;
        RECT -134.940 6.800 -134.170 10.680 ;
        RECT -135.130 6.320 -133.930 6.800 ;
        RECT -140.200 4.750 -138.780 5.160 ;
        RECT -139.870 -1.270 -139.100 4.750 ;
        RECT -134.940 -1.270 -134.170 6.320 ;
        RECT -129.960 5.160 -129.190 16.010 ;
        RECT -124.980 11.090 -124.210 16.010 ;
        RECT -125.320 10.680 -123.900 11.090 ;
        RECT -124.980 6.800 -124.210 10.680 ;
        RECT -125.210 6.320 -124.010 6.800 ;
        RECT -130.280 4.750 -128.860 5.160 ;
        RECT -129.960 -1.270 -129.190 4.750 ;
        RECT -124.980 -1.270 -124.210 6.320 ;
        RECT -120.060 5.160 -119.290 16.010 ;
        RECT -115.100 11.090 -114.330 16.010 ;
        RECT -115.400 10.680 -113.980 11.090 ;
        RECT -115.100 6.800 -114.330 10.680 ;
        RECT -115.290 6.320 -114.090 6.800 ;
        RECT -120.360 4.750 -118.940 5.160 ;
        RECT -120.060 -1.270 -119.290 4.750 ;
        RECT -115.100 -1.270 -114.330 6.320 ;
        RECT -110.130 5.160 -109.360 16.010 ;
        RECT -105.170 11.090 -104.400 16.010 ;
        RECT -105.480 10.680 -104.060 11.090 ;
        RECT -105.170 6.800 -104.400 10.680 ;
        RECT -105.370 6.320 -104.170 6.800 ;
        RECT -110.440 4.750 -109.020 5.160 ;
        RECT -110.130 -1.270 -109.360 4.750 ;
        RECT -105.170 -1.270 -104.400 6.320 ;
        RECT -100.180 5.160 -99.410 16.010 ;
        RECT -95.230 11.090 -94.460 16.010 ;
        RECT -95.560 10.680 -94.140 11.090 ;
        RECT -95.230 6.800 -94.460 10.680 ;
        RECT -95.450 6.320 -94.250 6.800 ;
        RECT -100.520 4.750 -99.100 5.160 ;
        RECT -100.180 -1.270 -99.410 4.750 ;
        RECT -95.230 -1.270 -94.460 6.320 ;
        RECT -90.280 5.160 -89.510 16.010 ;
        RECT -85.290 11.090 -84.520 16.010 ;
        RECT -85.640 10.680 -84.220 11.090 ;
        RECT -85.290 6.800 -84.520 10.680 ;
        RECT -85.530 6.320 -84.330 6.800 ;
        RECT -90.600 4.750 -89.180 5.160 ;
        RECT -90.280 -1.270 -89.510 4.750 ;
        RECT -85.290 -1.270 -84.520 6.320 ;
        RECT -80.370 5.160 -79.600 16.010 ;
        RECT -75.410 11.090 -74.640 16.010 ;
        RECT -75.720 10.680 -74.300 11.090 ;
        RECT -75.410 6.800 -74.640 10.680 ;
        RECT -75.610 6.320 -74.410 6.800 ;
        RECT -80.680 4.750 -79.260 5.160 ;
        RECT -80.370 -1.270 -79.600 4.750 ;
        RECT -75.410 -1.270 -74.640 6.320 ;
        RECT -70.430 5.160 -69.660 16.010 ;
        RECT -65.450 11.090 -64.680 16.010 ;
        RECT -65.800 10.680 -64.380 11.090 ;
        RECT -65.450 6.800 -64.680 10.680 ;
        RECT -65.690 6.320 -64.490 6.800 ;
        RECT -70.760 4.750 -69.340 5.160 ;
        RECT -70.430 -1.270 -69.660 4.750 ;
        RECT -65.450 -1.270 -64.680 6.320 ;
        RECT -60.540 5.160 -59.770 16.010 ;
        RECT -55.540 11.090 -54.770 16.010 ;
        RECT -55.880 10.680 -54.460 11.090 ;
        RECT -55.540 6.800 -54.770 10.680 ;
        RECT -55.770 6.320 -54.570 6.800 ;
        RECT -60.840 4.750 -59.420 5.160 ;
        RECT -60.540 -1.270 -59.770 4.750 ;
        RECT -55.540 -1.270 -54.770 6.320 ;
        RECT -50.580 5.160 -49.810 16.010 ;
        RECT -45.650 11.090 -44.880 16.010 ;
        RECT -45.960 10.680 -44.540 11.090 ;
        RECT -45.650 6.800 -44.880 10.680 ;
        RECT -45.850 6.320 -44.650 6.800 ;
        RECT -50.920 4.750 -49.500 5.160 ;
        RECT -50.580 -1.270 -49.810 4.750 ;
        RECT -45.650 -1.270 -44.880 6.320 ;
        RECT -40.700 5.160 -39.930 16.010 ;
        RECT -35.720 11.090 -34.950 16.010 ;
        RECT -36.040 10.680 -34.620 11.090 ;
        RECT -35.720 6.800 -34.950 10.680 ;
        RECT -35.930 6.320 -34.730 6.800 ;
        RECT -41.000 4.750 -39.580 5.160 ;
        RECT -40.700 -1.270 -39.930 4.750 ;
        RECT -35.720 -1.270 -34.950 6.320 ;
        RECT -30.770 5.160 -30.000 16.010 ;
        RECT -25.820 11.090 -25.050 16.010 ;
        RECT -26.120 10.680 -24.700 11.090 ;
        RECT -25.820 6.800 -25.050 10.680 ;
        RECT -26.010 6.320 -24.810 6.800 ;
        RECT -31.080 4.750 -29.660 5.160 ;
        RECT -30.770 -1.270 -30.000 4.750 ;
        RECT -25.820 -1.270 -25.050 6.320 ;
        RECT -20.840 5.160 -20.070 16.010 ;
        RECT -15.890 11.090 -15.120 16.010 ;
        RECT -16.200 10.680 -14.780 11.090 ;
        RECT -15.890 6.800 -15.120 10.680 ;
        RECT -16.090 6.320 -14.890 6.800 ;
        RECT -21.160 4.750 -19.740 5.160 ;
        RECT -20.840 -1.270 -20.070 4.750 ;
        RECT -15.890 -1.270 -15.120 6.320 ;
        RECT -10.940 5.160 -10.170 16.010 ;
        RECT -5.960 11.090 -5.190 16.010 ;
        RECT -6.280 10.680 -4.860 11.090 ;
        RECT -5.960 6.800 -5.190 10.680 ;
        RECT -6.170 6.320 -4.970 6.800 ;
        RECT -11.240 4.750 -9.820 5.160 ;
        RECT -10.940 -1.270 -10.170 4.750 ;
        RECT -5.960 -1.270 -5.190 6.320 ;
        RECT -1.010 5.160 -0.240 16.010 ;
        RECT 3.920 11.090 4.690 16.010 ;
        RECT 3.640 10.680 5.060 11.090 ;
        RECT 3.920 6.800 4.690 10.680 ;
        RECT 3.750 6.320 4.950 6.800 ;
        RECT -1.320 4.750 0.100 5.160 ;
        RECT -1.010 -1.270 -0.240 4.750 ;
        RECT 3.920 -1.270 4.690 6.320 ;
        RECT 8.920 5.160 9.690 16.010 ;
        RECT 13.870 11.090 14.640 16.010 ;
        RECT 13.560 10.680 14.980 11.090 ;
        RECT 13.870 6.800 14.640 10.680 ;
        RECT 13.670 6.320 14.870 6.800 ;
        RECT 8.600 4.750 10.020 5.160 ;
        RECT 8.920 -1.270 9.690 4.750 ;
        RECT 13.870 -1.270 14.640 6.320 ;
        RECT 18.850 5.160 19.620 16.010 ;
        RECT 23.860 11.090 24.630 16.010 ;
        RECT 23.480 10.680 24.630 11.090 ;
        RECT 23.860 6.800 24.630 10.680 ;
        RECT 23.590 6.320 24.420 6.800 ;
        RECT 18.520 4.750 19.940 5.160 ;
        RECT 18.850 -1.270 19.620 4.750 ;
        RECT 23.860 -1.270 24.630 6.320 ;
        RECT 27.310 -0.850 32.400 16.010 ;
        RECT 134.170 -0.850 160.570 73.570 ;
        RECT 25.680 -1.270 162.330 -0.850 ;
        RECT -300.770 -5.710 162.330 -1.270 ;
        RECT -319.260 -5.720 162.330 -5.710 ;
        RECT -337.530 -10.480 162.330 -5.720 ;
        RECT -337.530 -10.900 32.400 -10.480 ;
        RECT -337.530 -10.910 -295.680 -10.900 ;
        RECT -337.530 -10.930 -300.400 -10.910 ;
        RECT -337.530 -10.940 -318.670 -10.930 ;
        RECT -300.410 -63.310 -295.320 -63.130 ;
        RECT -57.010 -63.310 -19.850 -10.900 ;
        RECT 27.310 -11.030 32.400 -10.900 ;
        RECT 27.670 -63.310 32.760 -63.250 ;
        RECT -300.410 -72.940 32.760 -63.310 ;
        RECT -300.410 -90.220 -295.320 -72.940 ;
        RECT -293.280 -90.220 -292.510 -72.940 ;
        RECT -288.320 -83.790 -287.550 -72.940 ;
        RECT -283.360 -77.860 -282.590 -72.940 ;
        RECT -283.680 -78.270 -282.260 -77.860 ;
        RECT -283.360 -82.150 -282.590 -78.270 ;
        RECT -283.570 -82.630 -282.370 -82.150 ;
        RECT -288.640 -84.200 -287.220 -83.790 ;
        RECT -288.320 -90.220 -287.550 -84.200 ;
        RECT -283.360 -90.220 -282.590 -82.630 ;
        RECT -278.420 -83.790 -277.650 -72.940 ;
        RECT -273.440 -77.770 -272.670 -72.940 ;
        RECT -273.440 -77.860 -272.660 -77.770 ;
        RECT -273.760 -78.270 -272.340 -77.860 ;
        RECT -273.440 -80.220 -272.660 -78.270 ;
        RECT -273.480 -82.150 -272.660 -80.220 ;
        RECT -273.650 -82.630 -272.450 -82.150 ;
        RECT -278.720 -84.200 -277.300 -83.790 ;
        RECT -273.480 -84.120 -272.660 -82.630 ;
        RECT -268.470 -83.790 -267.700 -72.940 ;
        RECT -263.480 -77.860 -262.710 -72.940 ;
        RECT -263.840 -78.270 -262.420 -77.860 ;
        RECT -263.480 -82.150 -262.710 -78.270 ;
        RECT -263.730 -82.630 -262.530 -82.150 ;
        RECT -278.420 -90.220 -277.650 -84.200 ;
        RECT -273.490 -87.730 -272.660 -84.120 ;
        RECT -268.800 -84.200 -267.380 -83.790 ;
        RECT -273.490 -90.220 -272.670 -87.730 ;
        RECT -268.470 -90.220 -267.700 -84.200 ;
        RECT -263.480 -90.220 -262.710 -82.630 ;
        RECT -258.580 -83.790 -257.810 -72.940 ;
        RECT -253.590 -77.860 -252.820 -72.940 ;
        RECT -253.920 -78.270 -252.500 -77.860 ;
        RECT -253.590 -82.150 -252.820 -78.270 ;
        RECT -253.810 -82.630 -252.610 -82.150 ;
        RECT -258.880 -84.200 -257.460 -83.790 ;
        RECT -258.580 -90.220 -257.810 -84.200 ;
        RECT -253.590 -90.220 -252.820 -82.630 ;
        RECT -248.650 -83.790 -247.880 -72.940 ;
        RECT -243.680 -77.860 -242.910 -72.940 ;
        RECT -244.000 -78.270 -242.580 -77.860 ;
        RECT -243.680 -82.150 -242.910 -78.270 ;
        RECT -243.890 -82.630 -242.690 -82.150 ;
        RECT -248.960 -84.200 -247.540 -83.790 ;
        RECT -248.650 -90.220 -247.880 -84.200 ;
        RECT -243.680 -90.220 -242.910 -82.630 ;
        RECT -238.740 -83.790 -237.970 -72.940 ;
        RECT -233.780 -77.860 -233.010 -72.940 ;
        RECT -234.080 -78.270 -232.660 -77.860 ;
        RECT -233.780 -82.150 -233.010 -78.270 ;
        RECT -233.970 -82.630 -232.770 -82.150 ;
        RECT -239.040 -84.200 -237.620 -83.790 ;
        RECT -238.740 -90.220 -237.970 -84.200 ;
        RECT -233.780 -90.220 -233.010 -82.630 ;
        RECT -228.810 -83.790 -228.040 -72.940 ;
        RECT -223.840 -77.860 -223.070 -72.940 ;
        RECT -224.160 -78.270 -222.740 -77.860 ;
        RECT -223.840 -82.150 -223.070 -78.270 ;
        RECT -224.050 -82.630 -222.850 -82.150 ;
        RECT -229.120 -84.200 -227.700 -83.790 ;
        RECT -228.810 -90.220 -228.040 -84.200 ;
        RECT -223.840 -90.220 -223.070 -82.630 ;
        RECT -218.860 -83.790 -218.090 -72.940 ;
        RECT -213.900 -77.860 -213.130 -72.940 ;
        RECT -214.240 -78.270 -212.820 -77.860 ;
        RECT -213.900 -82.150 -213.130 -78.270 ;
        RECT -214.130 -82.630 -212.930 -82.150 ;
        RECT -219.200 -84.200 -217.780 -83.790 ;
        RECT -218.860 -90.220 -218.090 -84.200 ;
        RECT -213.900 -90.220 -213.130 -82.630 ;
        RECT -208.950 -83.790 -208.180 -72.940 ;
        RECT -204.010 -77.860 -203.240 -72.940 ;
        RECT -204.320 -78.270 -202.900 -77.860 ;
        RECT -204.010 -82.150 -203.240 -78.270 ;
        RECT -204.210 -82.630 -203.010 -82.150 ;
        RECT -209.280 -84.200 -207.860 -83.790 ;
        RECT -208.950 -90.220 -208.180 -84.200 ;
        RECT -204.010 -90.220 -203.240 -82.630 ;
        RECT -199.080 -83.790 -198.310 -72.940 ;
        RECT -194.080 -77.860 -193.310 -72.940 ;
        RECT -194.400 -78.270 -192.980 -77.860 ;
        RECT -194.080 -82.150 -193.310 -78.270 ;
        RECT -194.290 -82.630 -193.090 -82.150 ;
        RECT -199.360 -84.200 -197.940 -83.790 ;
        RECT -199.080 -90.220 -198.310 -84.200 ;
        RECT -194.080 -90.220 -193.310 -82.630 ;
        RECT -189.120 -83.790 -188.350 -72.940 ;
        RECT -184.170 -77.860 -183.400 -72.940 ;
        RECT -184.480 -78.270 -183.060 -77.860 ;
        RECT -184.170 -82.150 -183.400 -78.270 ;
        RECT -184.370 -82.630 -183.170 -82.150 ;
        RECT -189.440 -84.200 -188.020 -83.790 ;
        RECT -189.120 -90.220 -188.350 -84.200 ;
        RECT -184.170 -90.220 -183.400 -82.630 ;
        RECT -179.210 -83.790 -178.440 -72.940 ;
        RECT -174.220 -77.860 -173.450 -72.940 ;
        RECT -174.560 -78.270 -173.140 -77.860 ;
        RECT -174.220 -82.150 -173.450 -78.270 ;
        RECT -174.450 -82.630 -173.250 -82.150 ;
        RECT -179.520 -84.200 -178.100 -83.790 ;
        RECT -179.210 -90.220 -178.440 -84.200 ;
        RECT -174.220 -90.220 -173.450 -82.630 ;
        RECT -169.280 -83.790 -168.510 -72.940 ;
        RECT -164.280 -77.860 -163.510 -72.940 ;
        RECT -164.640 -78.270 -163.220 -77.860 ;
        RECT -164.280 -82.150 -163.510 -78.270 ;
        RECT -164.530 -82.630 -163.330 -82.150 ;
        RECT -169.600 -84.200 -168.180 -83.790 ;
        RECT -169.280 -90.220 -168.510 -84.200 ;
        RECT -164.280 -90.220 -163.510 -82.630 ;
        RECT -159.370 -83.790 -158.600 -72.940 ;
        RECT -154.420 -77.860 -153.650 -72.940 ;
        RECT -154.720 -78.270 -153.300 -77.860 ;
        RECT -154.420 -82.150 -153.650 -78.270 ;
        RECT -154.610 -82.630 -153.410 -82.150 ;
        RECT -159.680 -84.200 -158.260 -83.790 ;
        RECT -159.370 -90.220 -158.600 -84.200 ;
        RECT -154.420 -90.220 -153.650 -82.630 ;
        RECT -149.450 -83.790 -148.680 -72.940 ;
        RECT -144.490 -77.860 -143.720 -72.940 ;
        RECT -144.800 -78.270 -143.380 -77.860 ;
        RECT -144.490 -82.150 -143.720 -78.270 ;
        RECT -144.690 -82.630 -143.490 -82.150 ;
        RECT -149.760 -84.200 -148.340 -83.790 ;
        RECT -149.450 -90.220 -148.680 -84.200 ;
        RECT -144.490 -90.220 -143.720 -82.630 ;
        RECT -139.510 -83.790 -138.740 -72.940 ;
        RECT -134.580 -77.860 -133.810 -72.940 ;
        RECT -134.880 -78.270 -133.460 -77.860 ;
        RECT -134.580 -82.150 -133.810 -78.270 ;
        RECT -134.770 -82.630 -133.570 -82.150 ;
        RECT -139.840 -84.200 -138.420 -83.790 ;
        RECT -139.510 -90.220 -138.740 -84.200 ;
        RECT -134.580 -90.220 -133.810 -82.630 ;
        RECT -129.600 -83.790 -128.830 -72.940 ;
        RECT -124.620 -77.860 -123.850 -72.940 ;
        RECT -124.960 -78.270 -123.540 -77.860 ;
        RECT -124.620 -82.150 -123.850 -78.270 ;
        RECT -124.850 -82.630 -123.650 -82.150 ;
        RECT -129.920 -84.200 -128.500 -83.790 ;
        RECT -129.600 -90.220 -128.830 -84.200 ;
        RECT -124.620 -90.220 -123.850 -82.630 ;
        RECT -119.700 -83.790 -118.930 -72.940 ;
        RECT -114.740 -77.860 -113.970 -72.940 ;
        RECT -115.040 -78.270 -113.620 -77.860 ;
        RECT -114.740 -82.150 -113.970 -78.270 ;
        RECT -114.930 -82.630 -113.730 -82.150 ;
        RECT -120.000 -84.200 -118.580 -83.790 ;
        RECT -119.700 -90.220 -118.930 -84.200 ;
        RECT -114.740 -90.220 -113.970 -82.630 ;
        RECT -109.770 -83.790 -109.000 -72.940 ;
        RECT -104.810 -77.860 -104.040 -72.940 ;
        RECT -105.120 -78.270 -103.700 -77.860 ;
        RECT -104.810 -82.150 -104.040 -78.270 ;
        RECT -105.010 -82.630 -103.810 -82.150 ;
        RECT -110.080 -84.200 -108.660 -83.790 ;
        RECT -109.770 -90.220 -109.000 -84.200 ;
        RECT -104.810 -90.220 -104.040 -82.630 ;
        RECT -99.820 -83.790 -99.050 -72.940 ;
        RECT -94.870 -77.860 -94.100 -72.940 ;
        RECT -95.200 -78.270 -93.780 -77.860 ;
        RECT -94.870 -82.150 -94.100 -78.270 ;
        RECT -95.090 -82.630 -93.890 -82.150 ;
        RECT -100.160 -84.200 -98.740 -83.790 ;
        RECT -99.820 -90.220 -99.050 -84.200 ;
        RECT -94.870 -90.220 -94.100 -82.630 ;
        RECT -89.920 -83.790 -89.150 -72.940 ;
        RECT -84.930 -77.860 -84.160 -72.940 ;
        RECT -85.280 -78.270 -83.860 -77.860 ;
        RECT -84.930 -82.150 -84.160 -78.270 ;
        RECT -85.170 -82.630 -83.970 -82.150 ;
        RECT -90.240 -84.200 -88.820 -83.790 ;
        RECT -89.920 -90.220 -89.150 -84.200 ;
        RECT -84.930 -90.220 -84.160 -82.630 ;
        RECT -80.010 -83.790 -79.240 -72.940 ;
        RECT -75.050 -77.860 -74.280 -72.940 ;
        RECT -75.360 -78.270 -73.940 -77.860 ;
        RECT -75.050 -82.150 -74.280 -78.270 ;
        RECT -75.250 -82.630 -74.050 -82.150 ;
        RECT -80.320 -84.200 -78.900 -83.790 ;
        RECT -80.010 -90.220 -79.240 -84.200 ;
        RECT -75.050 -90.220 -74.280 -82.630 ;
        RECT -70.070 -83.790 -69.300 -72.940 ;
        RECT -65.090 -77.860 -64.320 -72.940 ;
        RECT -65.440 -78.270 -64.020 -77.860 ;
        RECT -65.090 -82.150 -64.320 -78.270 ;
        RECT -65.330 -82.630 -64.130 -82.150 ;
        RECT -70.400 -84.200 -68.980 -83.790 ;
        RECT -70.070 -90.220 -69.300 -84.200 ;
        RECT -65.090 -90.220 -64.320 -82.630 ;
        RECT -60.180 -83.790 -59.410 -72.940 ;
        RECT -55.180 -77.860 -54.410 -72.940 ;
        RECT -55.520 -78.270 -54.100 -77.860 ;
        RECT -55.180 -82.150 -54.410 -78.270 ;
        RECT -55.410 -82.630 -54.210 -82.150 ;
        RECT -60.480 -84.200 -59.060 -83.790 ;
        RECT -60.180 -90.220 -59.410 -84.200 ;
        RECT -55.180 -90.220 -54.410 -82.630 ;
        RECT -50.220 -83.790 -49.450 -72.940 ;
        RECT -45.290 -77.860 -44.520 -72.940 ;
        RECT -45.600 -78.270 -44.180 -77.860 ;
        RECT -45.290 -82.150 -44.520 -78.270 ;
        RECT -45.490 -82.630 -44.290 -82.150 ;
        RECT -50.560 -84.200 -49.140 -83.790 ;
        RECT -50.220 -90.220 -49.450 -84.200 ;
        RECT -45.290 -90.220 -44.520 -82.630 ;
        RECT -40.340 -83.790 -39.570 -72.940 ;
        RECT -35.360 -77.860 -34.590 -72.940 ;
        RECT -35.680 -78.270 -34.260 -77.860 ;
        RECT -35.360 -82.150 -34.590 -78.270 ;
        RECT -35.570 -82.630 -34.370 -82.150 ;
        RECT -40.640 -84.200 -39.220 -83.790 ;
        RECT -40.340 -90.220 -39.570 -84.200 ;
        RECT -35.360 -90.220 -34.590 -82.630 ;
        RECT -30.410 -83.790 -29.640 -72.940 ;
        RECT -25.460 -77.860 -24.690 -72.940 ;
        RECT -25.760 -78.270 -24.340 -77.860 ;
        RECT -25.460 -82.150 -24.690 -78.270 ;
        RECT -25.650 -82.630 -24.450 -82.150 ;
        RECT -30.720 -84.200 -29.300 -83.790 ;
        RECT -30.410 -90.220 -29.640 -84.200 ;
        RECT -25.460 -90.220 -24.690 -82.630 ;
        RECT -20.480 -83.790 -19.710 -72.940 ;
        RECT -15.530 -77.860 -14.760 -72.940 ;
        RECT -15.840 -78.270 -14.420 -77.860 ;
        RECT -15.530 -82.150 -14.760 -78.270 ;
        RECT -15.730 -82.630 -14.530 -82.150 ;
        RECT -20.800 -84.200 -19.380 -83.790 ;
        RECT -20.480 -90.220 -19.710 -84.200 ;
        RECT -15.530 -90.220 -14.760 -82.630 ;
        RECT -10.580 -83.790 -9.810 -72.940 ;
        RECT -5.600 -77.860 -4.830 -72.940 ;
        RECT -5.920 -78.270 -4.500 -77.860 ;
        RECT -5.600 -82.150 -4.830 -78.270 ;
        RECT -5.810 -82.630 -4.610 -82.150 ;
        RECT -10.880 -84.200 -9.460 -83.790 ;
        RECT -10.580 -90.220 -9.810 -84.200 ;
        RECT -5.600 -90.220 -4.830 -82.630 ;
        RECT -0.650 -83.790 0.120 -72.940 ;
        RECT 4.280 -77.860 5.050 -72.940 ;
        RECT 4.000 -78.270 5.420 -77.860 ;
        RECT 4.280 -82.150 5.050 -78.270 ;
        RECT 4.110 -82.630 5.310 -82.150 ;
        RECT -0.960 -84.200 0.460 -83.790 ;
        RECT -0.650 -90.220 0.120 -84.200 ;
        RECT 4.280 -90.220 5.050 -82.630 ;
        RECT 9.280 -83.790 10.050 -72.940 ;
        RECT 14.230 -77.860 15.000 -72.940 ;
        RECT 13.920 -78.270 15.340 -77.860 ;
        RECT 14.230 -82.150 15.000 -78.270 ;
        RECT 14.030 -82.630 15.230 -82.150 ;
        RECT 8.960 -84.200 10.380 -83.790 ;
        RECT 9.280 -90.220 10.050 -84.200 ;
        RECT 14.230 -90.220 15.000 -82.630 ;
        RECT 19.210 -83.790 19.980 -72.940 ;
        RECT 24.220 -77.860 24.990 -72.940 ;
        RECT 23.840 -78.270 24.990 -77.860 ;
        RECT 24.220 -82.150 24.990 -78.270 ;
        RECT 23.950 -82.630 24.780 -82.150 ;
        RECT 18.880 -84.200 20.300 -83.790 ;
        RECT 19.210 -90.220 19.980 -84.200 ;
        RECT 24.220 -90.220 24.990 -82.630 ;
        RECT 27.670 -89.800 32.760 -72.940 ;
        RECT 134.170 -89.800 160.570 -10.480 ;
        RECT 26.040 -90.220 162.690 -89.800 ;
        RECT -300.410 -94.660 162.690 -90.220 ;
        RECT -318.900 -94.670 162.690 -94.660 ;
        RECT -337.170 -99.430 162.690 -94.670 ;
        RECT -337.170 -99.850 32.760 -99.430 ;
        RECT -337.170 -99.860 -295.320 -99.850 ;
        RECT -337.170 -99.880 -300.040 -99.860 ;
        RECT -337.170 -99.890 -318.310 -99.880 ;
        RECT -302.170 -157.890 -297.080 -157.710 ;
        RECT -206.330 -157.890 -169.170 -99.850 ;
        RECT 27.670 -99.980 32.760 -99.850 ;
        RECT 25.910 -157.890 31.000 -157.830 ;
        RECT -302.170 -167.520 31.000 -157.890 ;
        RECT -302.170 -184.800 -297.080 -167.520 ;
        RECT -295.040 -184.800 -294.270 -167.520 ;
        RECT -290.080 -178.370 -289.310 -167.520 ;
        RECT -285.120 -172.440 -284.350 -167.520 ;
        RECT -285.440 -172.850 -284.020 -172.440 ;
        RECT -285.120 -176.730 -284.350 -172.850 ;
        RECT -285.330 -177.210 -284.130 -176.730 ;
        RECT -290.400 -178.780 -288.980 -178.370 ;
        RECT -290.080 -184.800 -289.310 -178.780 ;
        RECT -285.120 -184.800 -284.350 -177.210 ;
        RECT -280.180 -178.370 -279.410 -167.520 ;
        RECT -275.200 -172.350 -274.430 -167.520 ;
        RECT -275.200 -172.440 -274.420 -172.350 ;
        RECT -275.520 -172.850 -274.100 -172.440 ;
        RECT -275.200 -174.800 -274.420 -172.850 ;
        RECT -275.240 -176.730 -274.420 -174.800 ;
        RECT -275.410 -177.210 -274.210 -176.730 ;
        RECT -280.480 -178.780 -279.060 -178.370 ;
        RECT -275.240 -178.700 -274.420 -177.210 ;
        RECT -270.230 -178.370 -269.460 -167.520 ;
        RECT -265.240 -172.440 -264.470 -167.520 ;
        RECT -265.600 -172.850 -264.180 -172.440 ;
        RECT -265.240 -176.730 -264.470 -172.850 ;
        RECT -265.490 -177.210 -264.290 -176.730 ;
        RECT -280.180 -184.800 -279.410 -178.780 ;
        RECT -275.250 -182.310 -274.420 -178.700 ;
        RECT -270.560 -178.780 -269.140 -178.370 ;
        RECT -275.250 -184.800 -274.430 -182.310 ;
        RECT -270.230 -184.800 -269.460 -178.780 ;
        RECT -265.240 -184.800 -264.470 -177.210 ;
        RECT -260.340 -178.370 -259.570 -167.520 ;
        RECT -255.350 -172.440 -254.580 -167.520 ;
        RECT -255.680 -172.850 -254.260 -172.440 ;
        RECT -255.350 -176.730 -254.580 -172.850 ;
        RECT -255.570 -177.210 -254.370 -176.730 ;
        RECT -260.640 -178.780 -259.220 -178.370 ;
        RECT -260.340 -184.800 -259.570 -178.780 ;
        RECT -255.350 -184.800 -254.580 -177.210 ;
        RECT -250.410 -178.370 -249.640 -167.520 ;
        RECT -245.440 -172.440 -244.670 -167.520 ;
        RECT -245.760 -172.850 -244.340 -172.440 ;
        RECT -245.440 -176.730 -244.670 -172.850 ;
        RECT -245.650 -177.210 -244.450 -176.730 ;
        RECT -250.720 -178.780 -249.300 -178.370 ;
        RECT -250.410 -184.800 -249.640 -178.780 ;
        RECT -245.440 -184.800 -244.670 -177.210 ;
        RECT -240.500 -178.370 -239.730 -167.520 ;
        RECT -235.540 -172.440 -234.770 -167.520 ;
        RECT -235.840 -172.850 -234.420 -172.440 ;
        RECT -235.540 -176.730 -234.770 -172.850 ;
        RECT -235.730 -177.210 -234.530 -176.730 ;
        RECT -240.800 -178.780 -239.380 -178.370 ;
        RECT -240.500 -184.800 -239.730 -178.780 ;
        RECT -235.540 -184.800 -234.770 -177.210 ;
        RECT -230.570 -178.370 -229.800 -167.520 ;
        RECT -225.600 -172.440 -224.830 -167.520 ;
        RECT -225.920 -172.850 -224.500 -172.440 ;
        RECT -225.600 -176.730 -224.830 -172.850 ;
        RECT -225.810 -177.210 -224.610 -176.730 ;
        RECT -230.880 -178.780 -229.460 -178.370 ;
        RECT -230.570 -184.800 -229.800 -178.780 ;
        RECT -225.600 -184.800 -224.830 -177.210 ;
        RECT -220.620 -178.370 -219.850 -167.520 ;
        RECT -215.660 -172.440 -214.890 -167.520 ;
        RECT -216.000 -172.850 -214.580 -172.440 ;
        RECT -215.660 -176.730 -214.890 -172.850 ;
        RECT -215.890 -177.210 -214.690 -176.730 ;
        RECT -220.960 -178.780 -219.540 -178.370 ;
        RECT -220.620 -184.800 -219.850 -178.780 ;
        RECT -215.660 -184.800 -214.890 -177.210 ;
        RECT -210.710 -178.370 -209.940 -167.520 ;
        RECT -205.770 -172.440 -205.000 -167.520 ;
        RECT -206.080 -172.850 -204.660 -172.440 ;
        RECT -205.770 -176.730 -205.000 -172.850 ;
        RECT -205.970 -177.210 -204.770 -176.730 ;
        RECT -211.040 -178.780 -209.620 -178.370 ;
        RECT -210.710 -184.800 -209.940 -178.780 ;
        RECT -205.770 -184.800 -205.000 -177.210 ;
        RECT -200.840 -178.370 -200.070 -167.520 ;
        RECT -195.840 -172.440 -195.070 -167.520 ;
        RECT -196.160 -172.850 -194.740 -172.440 ;
        RECT -195.840 -176.730 -195.070 -172.850 ;
        RECT -196.050 -177.210 -194.850 -176.730 ;
        RECT -201.120 -178.780 -199.700 -178.370 ;
        RECT -200.840 -184.800 -200.070 -178.780 ;
        RECT -195.840 -184.800 -195.070 -177.210 ;
        RECT -190.880 -178.370 -190.110 -167.520 ;
        RECT -185.930 -172.440 -185.160 -167.520 ;
        RECT -186.240 -172.850 -184.820 -172.440 ;
        RECT -185.930 -176.730 -185.160 -172.850 ;
        RECT -186.130 -177.210 -184.930 -176.730 ;
        RECT -191.200 -178.780 -189.780 -178.370 ;
        RECT -190.880 -184.800 -190.110 -178.780 ;
        RECT -185.930 -184.800 -185.160 -177.210 ;
        RECT -180.970 -178.370 -180.200 -167.520 ;
        RECT -175.980 -172.440 -175.210 -167.520 ;
        RECT -176.320 -172.850 -174.900 -172.440 ;
        RECT -175.980 -176.730 -175.210 -172.850 ;
        RECT -176.210 -177.210 -175.010 -176.730 ;
        RECT -181.280 -178.780 -179.860 -178.370 ;
        RECT -180.970 -184.800 -180.200 -178.780 ;
        RECT -175.980 -184.800 -175.210 -177.210 ;
        RECT -171.040 -178.370 -170.270 -167.520 ;
        RECT -166.040 -172.440 -165.270 -167.520 ;
        RECT -166.400 -172.850 -164.980 -172.440 ;
        RECT -166.040 -176.730 -165.270 -172.850 ;
        RECT -166.290 -177.210 -165.090 -176.730 ;
        RECT -171.360 -178.780 -169.940 -178.370 ;
        RECT -171.040 -184.800 -170.270 -178.780 ;
        RECT -166.040 -184.800 -165.270 -177.210 ;
        RECT -161.130 -178.370 -160.360 -167.520 ;
        RECT -156.180 -172.440 -155.410 -167.520 ;
        RECT -156.480 -172.850 -155.060 -172.440 ;
        RECT -156.180 -176.730 -155.410 -172.850 ;
        RECT -156.370 -177.210 -155.170 -176.730 ;
        RECT -161.440 -178.780 -160.020 -178.370 ;
        RECT -161.130 -184.800 -160.360 -178.780 ;
        RECT -156.180 -184.800 -155.410 -177.210 ;
        RECT -151.210 -178.370 -150.440 -167.520 ;
        RECT -146.250 -172.440 -145.480 -167.520 ;
        RECT -146.560 -172.850 -145.140 -172.440 ;
        RECT -146.250 -176.730 -145.480 -172.850 ;
        RECT -146.450 -177.210 -145.250 -176.730 ;
        RECT -151.520 -178.780 -150.100 -178.370 ;
        RECT -151.210 -184.800 -150.440 -178.780 ;
        RECT -146.250 -184.800 -145.480 -177.210 ;
        RECT -141.270 -178.370 -140.500 -167.520 ;
        RECT -136.340 -172.440 -135.570 -167.520 ;
        RECT -136.640 -172.850 -135.220 -172.440 ;
        RECT -136.340 -176.730 -135.570 -172.850 ;
        RECT -136.530 -177.210 -135.330 -176.730 ;
        RECT -141.600 -178.780 -140.180 -178.370 ;
        RECT -141.270 -184.800 -140.500 -178.780 ;
        RECT -136.340 -184.800 -135.570 -177.210 ;
        RECT -131.360 -178.370 -130.590 -167.520 ;
        RECT -126.380 -172.440 -125.610 -167.520 ;
        RECT -126.720 -172.850 -125.300 -172.440 ;
        RECT -126.380 -176.730 -125.610 -172.850 ;
        RECT -126.610 -177.210 -125.410 -176.730 ;
        RECT -131.680 -178.780 -130.260 -178.370 ;
        RECT -131.360 -184.800 -130.590 -178.780 ;
        RECT -126.380 -184.800 -125.610 -177.210 ;
        RECT -121.460 -178.370 -120.690 -167.520 ;
        RECT -116.500 -172.440 -115.730 -167.520 ;
        RECT -116.800 -172.850 -115.380 -172.440 ;
        RECT -116.500 -176.730 -115.730 -172.850 ;
        RECT -116.690 -177.210 -115.490 -176.730 ;
        RECT -121.760 -178.780 -120.340 -178.370 ;
        RECT -121.460 -184.800 -120.690 -178.780 ;
        RECT -116.500 -184.800 -115.730 -177.210 ;
        RECT -111.530 -178.370 -110.760 -167.520 ;
        RECT -106.570 -172.440 -105.800 -167.520 ;
        RECT -106.880 -172.850 -105.460 -172.440 ;
        RECT -106.570 -176.730 -105.800 -172.850 ;
        RECT -106.770 -177.210 -105.570 -176.730 ;
        RECT -111.840 -178.780 -110.420 -178.370 ;
        RECT -111.530 -184.800 -110.760 -178.780 ;
        RECT -106.570 -184.800 -105.800 -177.210 ;
        RECT -101.580 -178.370 -100.810 -167.520 ;
        RECT -96.630 -172.440 -95.860 -167.520 ;
        RECT -96.960 -172.850 -95.540 -172.440 ;
        RECT -96.630 -176.730 -95.860 -172.850 ;
        RECT -96.850 -177.210 -95.650 -176.730 ;
        RECT -101.920 -178.780 -100.500 -178.370 ;
        RECT -101.580 -184.800 -100.810 -178.780 ;
        RECT -96.630 -184.800 -95.860 -177.210 ;
        RECT -91.680 -178.370 -90.910 -167.520 ;
        RECT -86.690 -172.440 -85.920 -167.520 ;
        RECT -87.040 -172.850 -85.620 -172.440 ;
        RECT -86.690 -176.730 -85.920 -172.850 ;
        RECT -86.930 -177.210 -85.730 -176.730 ;
        RECT -92.000 -178.780 -90.580 -178.370 ;
        RECT -91.680 -184.800 -90.910 -178.780 ;
        RECT -86.690 -184.800 -85.920 -177.210 ;
        RECT -81.770 -178.370 -81.000 -167.520 ;
        RECT -76.810 -172.440 -76.040 -167.520 ;
        RECT -77.120 -172.850 -75.700 -172.440 ;
        RECT -76.810 -176.730 -76.040 -172.850 ;
        RECT -77.010 -177.210 -75.810 -176.730 ;
        RECT -82.080 -178.780 -80.660 -178.370 ;
        RECT -81.770 -184.800 -81.000 -178.780 ;
        RECT -76.810 -184.800 -76.040 -177.210 ;
        RECT -71.830 -178.370 -71.060 -167.520 ;
        RECT -66.850 -172.440 -66.080 -167.520 ;
        RECT -67.200 -172.850 -65.780 -172.440 ;
        RECT -66.850 -176.730 -66.080 -172.850 ;
        RECT -67.090 -177.210 -65.890 -176.730 ;
        RECT -72.160 -178.780 -70.740 -178.370 ;
        RECT -71.830 -184.800 -71.060 -178.780 ;
        RECT -66.850 -184.800 -66.080 -177.210 ;
        RECT -61.940 -178.370 -61.170 -167.520 ;
        RECT -56.940 -172.440 -56.170 -167.520 ;
        RECT -57.280 -172.850 -55.860 -172.440 ;
        RECT -56.940 -176.730 -56.170 -172.850 ;
        RECT -57.170 -177.210 -55.970 -176.730 ;
        RECT -62.240 -178.780 -60.820 -178.370 ;
        RECT -61.940 -184.800 -61.170 -178.780 ;
        RECT -56.940 -184.800 -56.170 -177.210 ;
        RECT -51.980 -178.370 -51.210 -167.520 ;
        RECT -47.050 -172.440 -46.280 -167.520 ;
        RECT -47.360 -172.850 -45.940 -172.440 ;
        RECT -47.050 -176.730 -46.280 -172.850 ;
        RECT -47.250 -177.210 -46.050 -176.730 ;
        RECT -52.320 -178.780 -50.900 -178.370 ;
        RECT -51.980 -184.800 -51.210 -178.780 ;
        RECT -47.050 -184.800 -46.280 -177.210 ;
        RECT -42.100 -178.370 -41.330 -167.520 ;
        RECT -37.120 -172.440 -36.350 -167.520 ;
        RECT -37.440 -172.850 -36.020 -172.440 ;
        RECT -37.120 -176.730 -36.350 -172.850 ;
        RECT -37.330 -177.210 -36.130 -176.730 ;
        RECT -42.400 -178.780 -40.980 -178.370 ;
        RECT -42.100 -184.800 -41.330 -178.780 ;
        RECT -37.120 -184.800 -36.350 -177.210 ;
        RECT -32.170 -178.370 -31.400 -167.520 ;
        RECT -27.220 -172.440 -26.450 -167.520 ;
        RECT -27.520 -172.850 -26.100 -172.440 ;
        RECT -27.220 -176.730 -26.450 -172.850 ;
        RECT -27.410 -177.210 -26.210 -176.730 ;
        RECT -32.480 -178.780 -31.060 -178.370 ;
        RECT -32.170 -184.800 -31.400 -178.780 ;
        RECT -27.220 -184.800 -26.450 -177.210 ;
        RECT -22.240 -178.370 -21.470 -167.520 ;
        RECT -17.290 -172.440 -16.520 -167.520 ;
        RECT -17.600 -172.850 -16.180 -172.440 ;
        RECT -17.290 -176.730 -16.520 -172.850 ;
        RECT -17.490 -177.210 -16.290 -176.730 ;
        RECT -22.560 -178.780 -21.140 -178.370 ;
        RECT -22.240 -184.800 -21.470 -178.780 ;
        RECT -17.290 -184.800 -16.520 -177.210 ;
        RECT -12.340 -178.370 -11.570 -167.520 ;
        RECT -7.360 -172.440 -6.590 -167.520 ;
        RECT -7.680 -172.850 -6.260 -172.440 ;
        RECT -7.360 -176.730 -6.590 -172.850 ;
        RECT -7.570 -177.210 -6.370 -176.730 ;
        RECT -12.640 -178.780 -11.220 -178.370 ;
        RECT -12.340 -184.800 -11.570 -178.780 ;
        RECT -7.360 -184.800 -6.590 -177.210 ;
        RECT -2.410 -178.370 -1.640 -167.520 ;
        RECT 2.520 -172.440 3.290 -167.520 ;
        RECT 2.240 -172.850 3.660 -172.440 ;
        RECT 2.520 -176.730 3.290 -172.850 ;
        RECT 2.350 -177.210 3.550 -176.730 ;
        RECT -2.720 -178.780 -1.300 -178.370 ;
        RECT -2.410 -184.800 -1.640 -178.780 ;
        RECT 2.520 -184.800 3.290 -177.210 ;
        RECT 7.520 -178.370 8.290 -167.520 ;
        RECT 12.470 -172.440 13.240 -167.520 ;
        RECT 12.160 -172.850 13.580 -172.440 ;
        RECT 12.470 -176.730 13.240 -172.850 ;
        RECT 12.270 -177.210 13.470 -176.730 ;
        RECT 7.200 -178.780 8.620 -178.370 ;
        RECT 7.520 -184.800 8.290 -178.780 ;
        RECT 12.470 -184.800 13.240 -177.210 ;
        RECT 17.450 -178.370 18.220 -167.520 ;
        RECT 22.460 -172.440 23.230 -167.520 ;
        RECT 22.080 -172.850 23.230 -172.440 ;
        RECT 22.460 -176.730 23.230 -172.850 ;
        RECT 22.190 -177.210 23.020 -176.730 ;
        RECT 17.120 -178.780 18.540 -178.370 ;
        RECT 17.450 -184.800 18.220 -178.780 ;
        RECT 22.460 -184.800 23.230 -177.210 ;
        RECT 25.910 -184.380 31.000 -167.520 ;
        RECT 134.170 -184.380 160.570 -99.430 ;
        RECT 24.280 -184.800 160.930 -184.380 ;
        RECT -302.170 -189.240 160.930 -184.800 ;
        RECT -320.660 -189.250 160.930 -189.240 ;
        RECT -338.930 -194.010 160.930 -189.250 ;
        RECT -338.930 -194.430 31.000 -194.010 ;
        RECT -338.930 -194.440 -297.080 -194.430 ;
        RECT -338.930 -194.460 -301.800 -194.440 ;
        RECT -338.930 -194.470 -320.070 -194.460 ;
        RECT 25.910 -194.560 31.000 -194.430 ;
      LAYER via3 ;
        RECT -182.080 47.160 -172.340 57.620 ;
        RECT 143.900 49.220 151.510 56.120 ;
        RECT 143.990 40.090 151.600 46.990 ;
        RECT -42.060 -43.240 -32.320 -32.780 ;
        RECT 143.800 -35.490 151.410 -28.590 ;
        RECT 143.800 -44.910 151.410 -38.010 ;
        RECT -193.810 -132.560 -184.070 -122.100 ;
        RECT 143.620 -132.630 151.230 -125.730 ;
        RECT 143.590 -141.430 151.200 -134.530 ;
      LAYER met4 ;
        RECT -185.350 42.890 -124.840 61.310 ;
        RECT 140.410 39.640 156.210 57.390 ;
        RECT -45.270 -47.490 -29.510 -29.220 ;
        RECT 139.810 -45.690 155.570 -27.420 ;
        RECT -196.870 -136.790 -181.110 -118.520 ;
        RECT 139.810 -142.200 155.570 -123.930 ;
    END
  END vccd1
  OBS
      LAYER nwell ;
        RECT -290.950 95.095 -289.345 95.330 ;
        RECT -291.650 93.570 -289.345 95.095 ;
        RECT -291.650 93.510 -290.810 93.570 ;
      LAYER pwell ;
        RECT -290.860 93.225 -290.690 93.415 ;
        RECT 25.670 93.225 25.840 93.415 ;
        RECT -290.975 93.220 -289.625 93.225 ;
        RECT -291.440 93.140 -289.625 93.220 ;
        RECT -291.445 92.355 -289.625 93.140 ;
        RECT -291.440 92.350 -289.625 92.355 ;
        RECT -290.975 92.315 -289.625 92.350 ;
        RECT 24.605 93.220 25.955 93.225 ;
        RECT 24.605 93.140 26.420 93.220 ;
        RECT 24.605 92.355 26.425 93.140 ;
        RECT 24.605 92.320 26.420 92.355 ;
        RECT 24.605 92.315 25.955 92.320 ;
      LAYER nwell ;
        RECT -291.650 90.420 -289.430 92.025 ;
      LAYER pwell ;
        RECT -289.355 90.025 -288.575 90.175 ;
        RECT -289.545 90.020 -288.575 90.025 ;
        RECT -290.140 90.015 -288.575 90.020 ;
        RECT -290.145 89.230 -288.575 90.015 ;
        RECT -289.355 88.805 -288.575 89.230 ;
        RECT 23.555 90.025 24.335 90.175 ;
        RECT 23.555 90.020 24.525 90.025 ;
        RECT 23.555 88.810 25.130 90.020 ;
        RECT 23.555 88.805 24.335 88.810 ;
      LAYER nwell ;
        RECT -292.970 11.045 -291.365 11.280 ;
        RECT -293.670 9.520 -291.365 11.045 ;
        RECT -293.670 9.460 -292.830 9.520 ;
      LAYER pwell ;
        RECT -292.880 9.175 -292.710 9.365 ;
        RECT 23.650 9.175 23.820 9.365 ;
        RECT -292.995 9.170 -291.645 9.175 ;
        RECT -293.460 9.090 -291.645 9.170 ;
        RECT -293.465 8.305 -291.645 9.090 ;
        RECT -293.460 8.300 -291.645 8.305 ;
        RECT -292.995 8.265 -291.645 8.300 ;
        RECT 22.585 9.170 23.935 9.175 ;
        RECT 22.585 9.090 24.400 9.170 ;
        RECT 22.585 8.305 24.405 9.090 ;
        RECT 22.585 8.270 24.400 8.305 ;
        RECT 22.585 8.265 23.935 8.270 ;
      LAYER nwell ;
        RECT -293.670 6.370 -291.450 7.975 ;
      LAYER pwell ;
        RECT -291.375 5.975 -290.595 6.125 ;
        RECT -291.565 5.970 -290.595 5.975 ;
        RECT -292.160 5.965 -290.595 5.970 ;
        RECT -292.165 5.180 -290.595 5.965 ;
        RECT -291.375 4.755 -290.595 5.180 ;
        RECT 21.535 5.975 22.315 6.125 ;
        RECT 21.535 5.970 22.505 5.975 ;
        RECT 21.535 4.760 23.110 5.970 ;
        RECT 21.535 4.755 22.315 4.760 ;
      LAYER nwell ;
        RECT -292.610 -77.905 -291.005 -77.670 ;
        RECT -293.310 -79.430 -291.005 -77.905 ;
        RECT -293.310 -79.490 -292.470 -79.430 ;
      LAYER pwell ;
        RECT -292.520 -79.775 -292.350 -79.585 ;
        RECT 24.010 -79.775 24.180 -79.585 ;
        RECT -292.635 -79.780 -291.285 -79.775 ;
        RECT -293.100 -79.860 -291.285 -79.780 ;
        RECT -293.105 -80.645 -291.285 -79.860 ;
        RECT -293.100 -80.650 -291.285 -80.645 ;
        RECT -292.635 -80.685 -291.285 -80.650 ;
        RECT 22.945 -79.780 24.295 -79.775 ;
        RECT 22.945 -79.860 24.760 -79.780 ;
        RECT 22.945 -80.645 24.765 -79.860 ;
        RECT 22.945 -80.680 24.760 -80.645 ;
        RECT 22.945 -80.685 24.295 -80.680 ;
      LAYER nwell ;
        RECT -293.310 -82.580 -291.090 -80.975 ;
      LAYER pwell ;
        RECT -291.015 -82.975 -290.235 -82.825 ;
        RECT -291.205 -82.980 -290.235 -82.975 ;
        RECT -291.800 -82.985 -290.235 -82.980 ;
        RECT -291.805 -83.770 -290.235 -82.985 ;
        RECT -291.015 -84.195 -290.235 -83.770 ;
        RECT 21.895 -82.975 22.675 -82.825 ;
        RECT 21.895 -82.980 22.865 -82.975 ;
        RECT 21.895 -84.190 23.470 -82.980 ;
        RECT 21.895 -84.195 22.675 -84.190 ;
      LAYER nwell ;
        RECT -294.370 -172.485 -292.765 -172.250 ;
        RECT -295.070 -174.010 -292.765 -172.485 ;
        RECT -295.070 -174.070 -294.230 -174.010 ;
      LAYER pwell ;
        RECT -294.280 -174.355 -294.110 -174.165 ;
        RECT 22.250 -174.355 22.420 -174.165 ;
        RECT -294.395 -174.360 -293.045 -174.355 ;
        RECT -294.860 -174.440 -293.045 -174.360 ;
        RECT -294.865 -175.225 -293.045 -174.440 ;
        RECT -294.860 -175.230 -293.045 -175.225 ;
        RECT -294.395 -175.265 -293.045 -175.230 ;
        RECT 21.185 -174.360 22.535 -174.355 ;
        RECT 21.185 -174.440 23.000 -174.360 ;
        RECT 21.185 -175.225 23.005 -174.440 ;
        RECT 21.185 -175.260 23.000 -175.225 ;
        RECT 21.185 -175.265 22.535 -175.260 ;
      LAYER nwell ;
        RECT -295.070 -177.160 -292.850 -175.555 ;
      LAYER pwell ;
        RECT -292.775 -177.555 -291.995 -177.405 ;
        RECT -292.965 -177.560 -291.995 -177.555 ;
        RECT -293.560 -177.565 -291.995 -177.560 ;
        RECT -293.565 -178.350 -291.995 -177.565 ;
        RECT -292.775 -178.775 -291.995 -178.350 ;
        RECT 20.135 -177.555 20.915 -177.405 ;
        RECT 20.135 -177.560 21.105 -177.555 ;
        RECT 20.135 -178.770 21.710 -177.560 ;
        RECT 20.135 -178.775 20.915 -178.770 ;
      LAYER li1 ;
        RECT -290.845 94.990 -290.675 95.140 ;
        RECT -291.460 94.820 -290.675 94.990 ;
        RECT -291.375 93.655 -291.085 94.820 ;
        RECT -290.845 94.615 -290.675 94.820 ;
        RECT -290.505 94.875 -288.295 95.055 ;
        RECT -290.505 94.785 -289.600 94.875 ;
        RECT -288.800 94.795 -288.295 94.875 ;
        RECT -280.585 94.875 -278.375 95.055 ;
        RECT -280.585 94.785 -279.680 94.875 ;
        RECT -278.880 94.795 -278.375 94.875 ;
        RECT -270.665 94.875 -268.455 95.055 ;
        RECT -270.665 94.785 -269.760 94.875 ;
        RECT -268.960 94.795 -268.455 94.875 ;
        RECT -260.745 94.875 -258.535 95.055 ;
        RECT -260.745 94.785 -259.840 94.875 ;
        RECT -259.040 94.795 -258.535 94.875 ;
        RECT -250.825 94.875 -248.615 95.055 ;
        RECT -250.825 94.785 -249.920 94.875 ;
        RECT -249.120 94.795 -248.615 94.875 ;
        RECT -240.905 94.875 -238.695 95.055 ;
        RECT -240.905 94.785 -240.000 94.875 ;
        RECT -239.200 94.795 -238.695 94.875 ;
        RECT -230.985 94.875 -228.775 95.055 ;
        RECT -230.985 94.785 -230.080 94.875 ;
        RECT -229.280 94.795 -228.775 94.875 ;
        RECT -221.065 94.875 -218.855 95.055 ;
        RECT -221.065 94.785 -220.160 94.875 ;
        RECT -219.360 94.795 -218.855 94.875 ;
        RECT -211.145 94.875 -208.935 95.055 ;
        RECT -211.145 94.785 -210.240 94.875 ;
        RECT -209.440 94.795 -208.935 94.875 ;
        RECT -201.225 94.875 -199.015 95.055 ;
        RECT -201.225 94.785 -200.320 94.875 ;
        RECT -199.520 94.795 -199.015 94.875 ;
        RECT -191.305 94.875 -189.095 95.055 ;
        RECT -191.305 94.785 -190.400 94.875 ;
        RECT -189.600 94.795 -189.095 94.875 ;
        RECT -181.385 94.875 -179.175 95.055 ;
        RECT -181.385 94.785 -180.480 94.875 ;
        RECT -179.680 94.795 -179.175 94.875 ;
        RECT -171.465 94.875 -169.255 95.055 ;
        RECT -171.465 94.785 -170.560 94.875 ;
        RECT -169.760 94.795 -169.255 94.875 ;
        RECT -161.545 94.875 -159.335 95.055 ;
        RECT -161.545 94.785 -160.640 94.875 ;
        RECT -159.840 94.795 -159.335 94.875 ;
        RECT -151.625 94.875 -149.415 95.055 ;
        RECT -151.625 94.785 -150.720 94.875 ;
        RECT -149.920 94.795 -149.415 94.875 ;
        RECT -141.705 94.875 -139.495 95.055 ;
        RECT -141.705 94.785 -140.800 94.875 ;
        RECT -140.000 94.795 -139.495 94.875 ;
        RECT -131.785 94.875 -129.575 95.055 ;
        RECT -131.785 94.785 -130.880 94.875 ;
        RECT -130.080 94.795 -129.575 94.875 ;
        RECT -121.865 94.875 -119.655 95.055 ;
        RECT -121.865 94.785 -120.960 94.875 ;
        RECT -120.160 94.795 -119.655 94.875 ;
        RECT -111.945 94.875 -109.735 95.055 ;
        RECT -111.945 94.785 -111.040 94.875 ;
        RECT -110.240 94.795 -109.735 94.875 ;
        RECT -102.025 94.875 -99.815 95.055 ;
        RECT -102.025 94.785 -101.120 94.875 ;
        RECT -100.320 94.795 -99.815 94.875 ;
        RECT -92.105 94.875 -89.895 95.055 ;
        RECT -92.105 94.785 -91.200 94.875 ;
        RECT -90.400 94.795 -89.895 94.875 ;
        RECT -82.185 94.875 -79.975 95.055 ;
        RECT -82.185 94.785 -81.280 94.875 ;
        RECT -80.480 94.795 -79.975 94.875 ;
        RECT -72.265 94.875 -70.055 95.055 ;
        RECT -72.265 94.785 -71.360 94.875 ;
        RECT -70.560 94.795 -70.055 94.875 ;
        RECT -62.345 94.875 -60.135 95.055 ;
        RECT -62.345 94.785 -61.440 94.875 ;
        RECT -60.640 94.795 -60.135 94.875 ;
        RECT -52.425 94.875 -50.215 95.055 ;
        RECT -52.425 94.785 -51.520 94.875 ;
        RECT -50.720 94.795 -50.215 94.875 ;
        RECT -42.505 94.875 -40.295 95.055 ;
        RECT -42.505 94.785 -41.600 94.875 ;
        RECT -40.800 94.795 -40.295 94.875 ;
        RECT -32.585 94.875 -30.375 95.055 ;
        RECT -32.585 94.785 -31.680 94.875 ;
        RECT -30.880 94.795 -30.375 94.875 ;
        RECT -22.665 94.875 -20.455 95.055 ;
        RECT -22.665 94.785 -21.760 94.875 ;
        RECT -20.960 94.795 -20.455 94.875 ;
        RECT -12.745 94.875 -10.535 95.055 ;
        RECT -12.745 94.785 -11.840 94.875 ;
        RECT -11.040 94.795 -10.535 94.875 ;
        RECT -2.825 94.875 -0.615 95.055 ;
        RECT -2.825 94.785 -1.920 94.875 ;
        RECT -1.120 94.795 -0.615 94.875 ;
        RECT 7.095 94.875 9.305 95.055 ;
        RECT 7.095 94.785 8.000 94.875 ;
        RECT 8.800 94.795 9.305 94.875 ;
        RECT 17.015 94.875 19.225 95.055 ;
        RECT 17.015 94.785 17.920 94.875 ;
        RECT 18.720 94.795 19.225 94.875 ;
        RECT -290.845 94.285 -289.915 94.615 ;
        RECT -289.430 94.600 -289.100 94.705 ;
        RECT -283.440 94.600 -283.110 94.705 ;
        RECT -279.510 94.600 -279.180 94.705 ;
        RECT -273.520 94.600 -273.190 94.705 ;
        RECT -269.590 94.600 -269.260 94.705 ;
        RECT -263.600 94.600 -263.270 94.705 ;
        RECT -259.670 94.600 -259.340 94.705 ;
        RECT -253.680 94.600 -253.350 94.705 ;
        RECT -249.750 94.600 -249.420 94.705 ;
        RECT -243.760 94.600 -243.430 94.705 ;
        RECT -239.830 94.600 -239.500 94.705 ;
        RECT -233.840 94.600 -233.510 94.705 ;
        RECT -229.910 94.600 -229.580 94.705 ;
        RECT -223.920 94.600 -223.590 94.705 ;
        RECT -219.990 94.600 -219.660 94.705 ;
        RECT -214.000 94.600 -213.670 94.705 ;
        RECT -210.070 94.600 -209.740 94.705 ;
        RECT -204.080 94.600 -203.750 94.705 ;
        RECT -200.150 94.600 -199.820 94.705 ;
        RECT -194.160 94.600 -193.830 94.705 ;
        RECT -190.230 94.600 -189.900 94.705 ;
        RECT -184.240 94.600 -183.910 94.705 ;
        RECT -180.310 94.600 -179.980 94.705 ;
        RECT -174.320 94.600 -173.990 94.705 ;
        RECT -170.390 94.600 -170.060 94.705 ;
        RECT -164.400 94.600 -164.070 94.705 ;
        RECT -160.470 94.600 -160.140 94.705 ;
        RECT -154.480 94.600 -154.150 94.705 ;
        RECT -150.550 94.600 -150.220 94.705 ;
        RECT -144.560 94.600 -144.230 94.705 ;
        RECT -140.630 94.600 -140.300 94.705 ;
        RECT -134.640 94.600 -134.310 94.705 ;
        RECT -130.710 94.600 -130.380 94.705 ;
        RECT -124.720 94.600 -124.390 94.705 ;
        RECT -120.790 94.600 -120.460 94.705 ;
        RECT -114.800 94.600 -114.470 94.705 ;
        RECT -110.870 94.600 -110.540 94.705 ;
        RECT -104.880 94.600 -104.550 94.705 ;
        RECT -100.950 94.600 -100.620 94.705 ;
        RECT -94.960 94.600 -94.630 94.705 ;
        RECT -91.030 94.600 -90.700 94.705 ;
        RECT -85.040 94.600 -84.710 94.705 ;
        RECT -81.110 94.600 -80.780 94.705 ;
        RECT -75.120 94.600 -74.790 94.705 ;
        RECT -71.190 94.600 -70.860 94.705 ;
        RECT -65.200 94.600 -64.870 94.705 ;
        RECT -61.270 94.600 -60.940 94.705 ;
        RECT -55.280 94.600 -54.950 94.705 ;
        RECT -51.350 94.600 -51.020 94.705 ;
        RECT -45.360 94.600 -45.030 94.705 ;
        RECT -41.430 94.600 -41.100 94.705 ;
        RECT -35.440 94.600 -35.110 94.705 ;
        RECT -31.510 94.600 -31.180 94.705 ;
        RECT -25.520 94.600 -25.190 94.705 ;
        RECT -21.590 94.600 -21.260 94.705 ;
        RECT -15.600 94.600 -15.270 94.705 ;
        RECT -11.670 94.600 -11.340 94.705 ;
        RECT -5.680 94.600 -5.350 94.705 ;
        RECT -1.750 94.600 -1.420 94.705 ;
        RECT 4.240 94.600 4.570 94.705 ;
        RECT 8.170 94.600 8.500 94.705 ;
        RECT 14.160 94.600 14.490 94.705 ;
        RECT 18.090 94.600 18.420 94.705 ;
        RECT 24.080 94.600 24.410 94.705 ;
        RECT -289.745 94.430 -288.675 94.600 ;
        RECT -290.845 93.760 -290.675 94.285 ;
        RECT -289.745 94.105 -289.575 94.430 ;
        RECT -290.505 93.925 -289.575 94.105 ;
        RECT -289.395 93.865 -289.025 94.205 ;
        RECT -288.845 94.105 -288.675 94.430 ;
        RECT -283.865 94.430 -282.795 94.600 ;
        RECT -283.865 94.105 -283.695 94.430 ;
        RECT -288.845 93.935 -288.295 94.105 ;
        RECT -284.245 93.935 -283.695 94.105 ;
        RECT -283.515 93.865 -283.145 94.205 ;
        RECT -282.965 94.105 -282.795 94.430 ;
        RECT -279.825 94.430 -278.755 94.600 ;
        RECT -279.825 94.105 -279.655 94.430 ;
        RECT -282.965 93.925 -282.035 94.105 ;
        RECT -280.585 93.925 -279.655 94.105 ;
        RECT -279.475 93.865 -279.105 94.205 ;
        RECT -278.925 94.105 -278.755 94.430 ;
        RECT -273.945 94.430 -272.875 94.600 ;
        RECT -273.945 94.105 -273.775 94.430 ;
        RECT -278.925 93.935 -278.375 94.105 ;
        RECT -274.325 93.935 -273.775 94.105 ;
        RECT -273.595 93.865 -273.225 94.205 ;
        RECT -273.045 94.105 -272.875 94.430 ;
        RECT -269.905 94.430 -268.835 94.600 ;
        RECT -269.905 94.105 -269.735 94.430 ;
        RECT -273.045 93.925 -272.115 94.105 ;
        RECT -270.665 93.925 -269.735 94.105 ;
        RECT -269.555 93.865 -269.185 94.205 ;
        RECT -269.005 94.105 -268.835 94.430 ;
        RECT -264.025 94.430 -262.955 94.600 ;
        RECT -264.025 94.105 -263.855 94.430 ;
        RECT -269.005 93.935 -268.455 94.105 ;
        RECT -264.405 93.935 -263.855 94.105 ;
        RECT -263.675 93.865 -263.305 94.205 ;
        RECT -263.125 94.105 -262.955 94.430 ;
        RECT -259.985 94.430 -258.915 94.600 ;
        RECT -259.985 94.105 -259.815 94.430 ;
        RECT -263.125 93.925 -262.195 94.105 ;
        RECT -260.745 93.925 -259.815 94.105 ;
        RECT -259.635 93.865 -259.265 94.205 ;
        RECT -259.085 94.105 -258.915 94.430 ;
        RECT -254.105 94.430 -253.035 94.600 ;
        RECT -254.105 94.105 -253.935 94.430 ;
        RECT -259.085 93.935 -258.535 94.105 ;
        RECT -254.485 93.935 -253.935 94.105 ;
        RECT -253.755 93.865 -253.385 94.205 ;
        RECT -253.205 94.105 -253.035 94.430 ;
        RECT -250.065 94.430 -248.995 94.600 ;
        RECT -250.065 94.105 -249.895 94.430 ;
        RECT -253.205 93.925 -252.275 94.105 ;
        RECT -250.825 93.925 -249.895 94.105 ;
        RECT -249.715 93.865 -249.345 94.205 ;
        RECT -249.165 94.105 -248.995 94.430 ;
        RECT -244.185 94.430 -243.115 94.600 ;
        RECT -244.185 94.105 -244.015 94.430 ;
        RECT -249.165 93.935 -248.615 94.105 ;
        RECT -244.565 93.935 -244.015 94.105 ;
        RECT -243.835 93.865 -243.465 94.205 ;
        RECT -243.285 94.105 -243.115 94.430 ;
        RECT -240.145 94.430 -239.075 94.600 ;
        RECT -240.145 94.105 -239.975 94.430 ;
        RECT -243.285 93.925 -242.355 94.105 ;
        RECT -240.905 93.925 -239.975 94.105 ;
        RECT -239.795 93.865 -239.425 94.205 ;
        RECT -239.245 94.105 -239.075 94.430 ;
        RECT -234.265 94.430 -233.195 94.600 ;
        RECT -234.265 94.105 -234.095 94.430 ;
        RECT -239.245 93.935 -238.695 94.105 ;
        RECT -234.645 93.935 -234.095 94.105 ;
        RECT -233.915 93.865 -233.545 94.205 ;
        RECT -233.365 94.105 -233.195 94.430 ;
        RECT -230.225 94.430 -229.155 94.600 ;
        RECT -230.225 94.105 -230.055 94.430 ;
        RECT -233.365 93.925 -232.435 94.105 ;
        RECT -230.985 93.925 -230.055 94.105 ;
        RECT -229.875 93.865 -229.505 94.205 ;
        RECT -229.325 94.105 -229.155 94.430 ;
        RECT -224.345 94.430 -223.275 94.600 ;
        RECT -224.345 94.105 -224.175 94.430 ;
        RECT -229.325 93.935 -228.775 94.105 ;
        RECT -224.725 93.935 -224.175 94.105 ;
        RECT -223.995 93.865 -223.625 94.205 ;
        RECT -223.445 94.105 -223.275 94.430 ;
        RECT -220.305 94.430 -219.235 94.600 ;
        RECT -220.305 94.105 -220.135 94.430 ;
        RECT -223.445 93.925 -222.515 94.105 ;
        RECT -221.065 93.925 -220.135 94.105 ;
        RECT -219.955 93.865 -219.585 94.205 ;
        RECT -219.405 94.105 -219.235 94.430 ;
        RECT -214.425 94.430 -213.355 94.600 ;
        RECT -214.425 94.105 -214.255 94.430 ;
        RECT -219.405 93.935 -218.855 94.105 ;
        RECT -214.805 93.935 -214.255 94.105 ;
        RECT -214.075 93.865 -213.705 94.205 ;
        RECT -213.525 94.105 -213.355 94.430 ;
        RECT -210.385 94.430 -209.315 94.600 ;
        RECT -210.385 94.105 -210.215 94.430 ;
        RECT -213.525 93.925 -212.595 94.105 ;
        RECT -211.145 93.925 -210.215 94.105 ;
        RECT -210.035 93.865 -209.665 94.205 ;
        RECT -209.485 94.105 -209.315 94.430 ;
        RECT -204.505 94.430 -203.435 94.600 ;
        RECT -204.505 94.105 -204.335 94.430 ;
        RECT -209.485 93.935 -208.935 94.105 ;
        RECT -204.885 93.935 -204.335 94.105 ;
        RECT -204.155 93.865 -203.785 94.205 ;
        RECT -203.605 94.105 -203.435 94.430 ;
        RECT -200.465 94.430 -199.395 94.600 ;
        RECT -200.465 94.105 -200.295 94.430 ;
        RECT -203.605 93.925 -202.675 94.105 ;
        RECT -201.225 93.925 -200.295 94.105 ;
        RECT -200.115 93.865 -199.745 94.205 ;
        RECT -199.565 94.105 -199.395 94.430 ;
        RECT -194.585 94.430 -193.515 94.600 ;
        RECT -194.585 94.105 -194.415 94.430 ;
        RECT -199.565 93.935 -199.015 94.105 ;
        RECT -194.965 93.935 -194.415 94.105 ;
        RECT -194.235 93.865 -193.865 94.205 ;
        RECT -193.685 94.105 -193.515 94.430 ;
        RECT -190.545 94.430 -189.475 94.600 ;
        RECT -190.545 94.105 -190.375 94.430 ;
        RECT -193.685 93.925 -192.755 94.105 ;
        RECT -191.305 93.925 -190.375 94.105 ;
        RECT -190.195 93.865 -189.825 94.205 ;
        RECT -189.645 94.105 -189.475 94.430 ;
        RECT -184.665 94.430 -183.595 94.600 ;
        RECT -184.665 94.105 -184.495 94.430 ;
        RECT -189.645 93.935 -189.095 94.105 ;
        RECT -185.045 93.935 -184.495 94.105 ;
        RECT -184.315 93.865 -183.945 94.205 ;
        RECT -183.765 94.105 -183.595 94.430 ;
        RECT -180.625 94.430 -179.555 94.600 ;
        RECT -180.625 94.105 -180.455 94.430 ;
        RECT -183.765 93.925 -182.835 94.105 ;
        RECT -181.385 93.925 -180.455 94.105 ;
        RECT -180.275 93.865 -179.905 94.205 ;
        RECT -179.725 94.105 -179.555 94.430 ;
        RECT -174.745 94.430 -173.675 94.600 ;
        RECT -174.745 94.105 -174.575 94.430 ;
        RECT -179.725 93.935 -179.175 94.105 ;
        RECT -175.125 93.935 -174.575 94.105 ;
        RECT -174.395 93.865 -174.025 94.205 ;
        RECT -173.845 94.105 -173.675 94.430 ;
        RECT -170.705 94.430 -169.635 94.600 ;
        RECT -170.705 94.105 -170.535 94.430 ;
        RECT -173.845 93.925 -172.915 94.105 ;
        RECT -171.465 93.925 -170.535 94.105 ;
        RECT -170.355 93.865 -169.985 94.205 ;
        RECT -169.805 94.105 -169.635 94.430 ;
        RECT -164.825 94.430 -163.755 94.600 ;
        RECT -164.825 94.105 -164.655 94.430 ;
        RECT -169.805 93.935 -169.255 94.105 ;
        RECT -165.205 93.935 -164.655 94.105 ;
        RECT -164.475 93.865 -164.105 94.205 ;
        RECT -163.925 94.105 -163.755 94.430 ;
        RECT -160.785 94.430 -159.715 94.600 ;
        RECT -160.785 94.105 -160.615 94.430 ;
        RECT -163.925 93.925 -162.995 94.105 ;
        RECT -161.545 93.925 -160.615 94.105 ;
        RECT -160.435 93.865 -160.065 94.205 ;
        RECT -159.885 94.105 -159.715 94.430 ;
        RECT -154.905 94.430 -153.835 94.600 ;
        RECT -154.905 94.105 -154.735 94.430 ;
        RECT -159.885 93.935 -159.335 94.105 ;
        RECT -155.285 93.935 -154.735 94.105 ;
        RECT -154.555 93.865 -154.185 94.205 ;
        RECT -154.005 94.105 -153.835 94.430 ;
        RECT -150.865 94.430 -149.795 94.600 ;
        RECT -150.865 94.105 -150.695 94.430 ;
        RECT -154.005 93.925 -153.075 94.105 ;
        RECT -151.625 93.925 -150.695 94.105 ;
        RECT -150.515 93.865 -150.145 94.205 ;
        RECT -149.965 94.105 -149.795 94.430 ;
        RECT -144.985 94.430 -143.915 94.600 ;
        RECT -144.985 94.105 -144.815 94.430 ;
        RECT -149.965 93.935 -149.415 94.105 ;
        RECT -145.365 93.935 -144.815 94.105 ;
        RECT -144.635 93.865 -144.265 94.205 ;
        RECT -144.085 94.105 -143.915 94.430 ;
        RECT -140.945 94.430 -139.875 94.600 ;
        RECT -140.945 94.105 -140.775 94.430 ;
        RECT -144.085 93.925 -143.155 94.105 ;
        RECT -141.705 93.925 -140.775 94.105 ;
        RECT -140.595 93.865 -140.225 94.205 ;
        RECT -140.045 94.105 -139.875 94.430 ;
        RECT -135.065 94.430 -133.995 94.600 ;
        RECT -135.065 94.105 -134.895 94.430 ;
        RECT -140.045 93.935 -139.495 94.105 ;
        RECT -135.445 93.935 -134.895 94.105 ;
        RECT -134.715 93.865 -134.345 94.205 ;
        RECT -134.165 94.105 -133.995 94.430 ;
        RECT -131.025 94.430 -129.955 94.600 ;
        RECT -131.025 94.105 -130.855 94.430 ;
        RECT -134.165 93.925 -133.235 94.105 ;
        RECT -131.785 93.925 -130.855 94.105 ;
        RECT -130.675 93.865 -130.305 94.205 ;
        RECT -130.125 94.105 -129.955 94.430 ;
        RECT -125.145 94.430 -124.075 94.600 ;
        RECT -125.145 94.105 -124.975 94.430 ;
        RECT -130.125 93.935 -129.575 94.105 ;
        RECT -125.525 93.935 -124.975 94.105 ;
        RECT -124.795 93.865 -124.425 94.205 ;
        RECT -124.245 94.105 -124.075 94.430 ;
        RECT -121.105 94.430 -120.035 94.600 ;
        RECT -121.105 94.105 -120.935 94.430 ;
        RECT -124.245 93.925 -123.315 94.105 ;
        RECT -121.865 93.925 -120.935 94.105 ;
        RECT -120.755 93.865 -120.385 94.205 ;
        RECT -120.205 94.105 -120.035 94.430 ;
        RECT -115.225 94.430 -114.155 94.600 ;
        RECT -115.225 94.105 -115.055 94.430 ;
        RECT -120.205 93.935 -119.655 94.105 ;
        RECT -115.605 93.935 -115.055 94.105 ;
        RECT -114.875 93.865 -114.505 94.205 ;
        RECT -114.325 94.105 -114.155 94.430 ;
        RECT -111.185 94.430 -110.115 94.600 ;
        RECT -111.185 94.105 -111.015 94.430 ;
        RECT -114.325 93.925 -113.395 94.105 ;
        RECT -111.945 93.925 -111.015 94.105 ;
        RECT -110.835 93.865 -110.465 94.205 ;
        RECT -110.285 94.105 -110.115 94.430 ;
        RECT -105.305 94.430 -104.235 94.600 ;
        RECT -105.305 94.105 -105.135 94.430 ;
        RECT -110.285 93.935 -109.735 94.105 ;
        RECT -105.685 93.935 -105.135 94.105 ;
        RECT -104.955 93.865 -104.585 94.205 ;
        RECT -104.405 94.105 -104.235 94.430 ;
        RECT -101.265 94.430 -100.195 94.600 ;
        RECT -101.265 94.105 -101.095 94.430 ;
        RECT -104.405 93.925 -103.475 94.105 ;
        RECT -102.025 93.925 -101.095 94.105 ;
        RECT -100.915 93.865 -100.545 94.205 ;
        RECT -100.365 94.105 -100.195 94.430 ;
        RECT -95.385 94.430 -94.315 94.600 ;
        RECT -95.385 94.105 -95.215 94.430 ;
        RECT -100.365 93.935 -99.815 94.105 ;
        RECT -95.765 93.935 -95.215 94.105 ;
        RECT -95.035 93.865 -94.665 94.205 ;
        RECT -94.485 94.105 -94.315 94.430 ;
        RECT -91.345 94.430 -90.275 94.600 ;
        RECT -91.345 94.105 -91.175 94.430 ;
        RECT -94.485 93.925 -93.555 94.105 ;
        RECT -92.105 93.925 -91.175 94.105 ;
        RECT -90.995 93.865 -90.625 94.205 ;
        RECT -90.445 94.105 -90.275 94.430 ;
        RECT -85.465 94.430 -84.395 94.600 ;
        RECT -85.465 94.105 -85.295 94.430 ;
        RECT -90.445 93.935 -89.895 94.105 ;
        RECT -85.845 93.935 -85.295 94.105 ;
        RECT -85.115 93.865 -84.745 94.205 ;
        RECT -84.565 94.105 -84.395 94.430 ;
        RECT -81.425 94.430 -80.355 94.600 ;
        RECT -81.425 94.105 -81.255 94.430 ;
        RECT -84.565 93.925 -83.635 94.105 ;
        RECT -82.185 93.925 -81.255 94.105 ;
        RECT -81.075 93.865 -80.705 94.205 ;
        RECT -80.525 94.105 -80.355 94.430 ;
        RECT -75.545 94.430 -74.475 94.600 ;
        RECT -75.545 94.105 -75.375 94.430 ;
        RECT -80.525 93.935 -79.975 94.105 ;
        RECT -75.925 93.935 -75.375 94.105 ;
        RECT -75.195 93.865 -74.825 94.205 ;
        RECT -74.645 94.105 -74.475 94.430 ;
        RECT -71.505 94.430 -70.435 94.600 ;
        RECT -71.505 94.105 -71.335 94.430 ;
        RECT -74.645 93.925 -73.715 94.105 ;
        RECT -72.265 93.925 -71.335 94.105 ;
        RECT -71.155 93.865 -70.785 94.205 ;
        RECT -70.605 94.105 -70.435 94.430 ;
        RECT -65.625 94.430 -64.555 94.600 ;
        RECT -65.625 94.105 -65.455 94.430 ;
        RECT -70.605 93.935 -70.055 94.105 ;
        RECT -66.005 93.935 -65.455 94.105 ;
        RECT -65.275 93.865 -64.905 94.205 ;
        RECT -64.725 94.105 -64.555 94.430 ;
        RECT -61.585 94.430 -60.515 94.600 ;
        RECT -61.585 94.105 -61.415 94.430 ;
        RECT -64.725 93.925 -63.795 94.105 ;
        RECT -62.345 93.925 -61.415 94.105 ;
        RECT -61.235 93.865 -60.865 94.205 ;
        RECT -60.685 94.105 -60.515 94.430 ;
        RECT -55.705 94.430 -54.635 94.600 ;
        RECT -55.705 94.105 -55.535 94.430 ;
        RECT -60.685 93.935 -60.135 94.105 ;
        RECT -56.085 93.935 -55.535 94.105 ;
        RECT -55.355 93.865 -54.985 94.205 ;
        RECT -54.805 94.105 -54.635 94.430 ;
        RECT -51.665 94.430 -50.595 94.600 ;
        RECT -51.665 94.105 -51.495 94.430 ;
        RECT -54.805 93.925 -53.875 94.105 ;
        RECT -52.425 93.925 -51.495 94.105 ;
        RECT -51.315 93.865 -50.945 94.205 ;
        RECT -50.765 94.105 -50.595 94.430 ;
        RECT -45.785 94.430 -44.715 94.600 ;
        RECT -45.785 94.105 -45.615 94.430 ;
        RECT -50.765 93.935 -50.215 94.105 ;
        RECT -46.165 93.935 -45.615 94.105 ;
        RECT -45.435 93.865 -45.065 94.205 ;
        RECT -44.885 94.105 -44.715 94.430 ;
        RECT -41.745 94.430 -40.675 94.600 ;
        RECT -41.745 94.105 -41.575 94.430 ;
        RECT -44.885 93.925 -43.955 94.105 ;
        RECT -42.505 93.925 -41.575 94.105 ;
        RECT -41.395 93.865 -41.025 94.205 ;
        RECT -40.845 94.105 -40.675 94.430 ;
        RECT -35.865 94.430 -34.795 94.600 ;
        RECT -35.865 94.105 -35.695 94.430 ;
        RECT -40.845 93.935 -40.295 94.105 ;
        RECT -36.245 93.935 -35.695 94.105 ;
        RECT -35.515 93.865 -35.145 94.205 ;
        RECT -34.965 94.105 -34.795 94.430 ;
        RECT -31.825 94.430 -30.755 94.600 ;
        RECT -31.825 94.105 -31.655 94.430 ;
        RECT -34.965 93.925 -34.035 94.105 ;
        RECT -32.585 93.925 -31.655 94.105 ;
        RECT -31.475 93.865 -31.105 94.205 ;
        RECT -30.925 94.105 -30.755 94.430 ;
        RECT -25.945 94.430 -24.875 94.600 ;
        RECT -25.945 94.105 -25.775 94.430 ;
        RECT -30.925 93.935 -30.375 94.105 ;
        RECT -26.325 93.935 -25.775 94.105 ;
        RECT -25.595 93.865 -25.225 94.205 ;
        RECT -25.045 94.105 -24.875 94.430 ;
        RECT -21.905 94.430 -20.835 94.600 ;
        RECT -21.905 94.105 -21.735 94.430 ;
        RECT -25.045 93.925 -24.115 94.105 ;
        RECT -22.665 93.925 -21.735 94.105 ;
        RECT -21.555 93.865 -21.185 94.205 ;
        RECT -21.005 94.105 -20.835 94.430 ;
        RECT -16.025 94.430 -14.955 94.600 ;
        RECT -16.025 94.105 -15.855 94.430 ;
        RECT -21.005 93.935 -20.455 94.105 ;
        RECT -16.405 93.935 -15.855 94.105 ;
        RECT -15.675 93.865 -15.305 94.205 ;
        RECT -15.125 94.105 -14.955 94.430 ;
        RECT -11.985 94.430 -10.915 94.600 ;
        RECT -11.985 94.105 -11.815 94.430 ;
        RECT -15.125 93.925 -14.195 94.105 ;
        RECT -12.745 93.925 -11.815 94.105 ;
        RECT -11.635 93.865 -11.265 94.205 ;
        RECT -11.085 94.105 -10.915 94.430 ;
        RECT -6.105 94.430 -5.035 94.600 ;
        RECT -6.105 94.105 -5.935 94.430 ;
        RECT -11.085 93.935 -10.535 94.105 ;
        RECT -6.485 93.935 -5.935 94.105 ;
        RECT -5.755 93.865 -5.385 94.205 ;
        RECT -5.205 94.105 -5.035 94.430 ;
        RECT -2.065 94.430 -0.995 94.600 ;
        RECT -2.065 94.105 -1.895 94.430 ;
        RECT -5.205 93.925 -4.275 94.105 ;
        RECT -2.825 93.925 -1.895 94.105 ;
        RECT -1.715 93.865 -1.345 94.205 ;
        RECT -1.165 94.105 -0.995 94.430 ;
        RECT 3.815 94.430 4.885 94.600 ;
        RECT 3.815 94.105 3.985 94.430 ;
        RECT -1.165 93.935 -0.615 94.105 ;
        RECT 3.435 93.935 3.985 94.105 ;
        RECT 4.165 93.865 4.535 94.205 ;
        RECT 4.715 94.105 4.885 94.430 ;
        RECT 7.855 94.430 8.925 94.600 ;
        RECT 7.855 94.105 8.025 94.430 ;
        RECT 4.715 93.925 5.645 94.105 ;
        RECT 7.095 93.925 8.025 94.105 ;
        RECT 8.205 93.865 8.575 94.205 ;
        RECT 8.755 94.105 8.925 94.430 ;
        RECT 13.735 94.430 14.805 94.600 ;
        RECT 13.735 94.105 13.905 94.430 ;
        RECT 8.755 93.935 9.305 94.105 ;
        RECT 13.355 93.935 13.905 94.105 ;
        RECT 14.085 93.865 14.455 94.205 ;
        RECT 14.635 94.105 14.805 94.430 ;
        RECT 17.775 94.430 18.845 94.600 ;
        RECT 17.775 94.105 17.945 94.430 ;
        RECT 14.635 93.925 15.565 94.105 ;
        RECT 17.015 93.925 17.945 94.105 ;
        RECT 18.125 93.865 18.495 94.205 ;
        RECT 18.675 94.105 18.845 94.430 ;
        RECT 23.655 94.430 24.725 94.600 ;
        RECT 23.655 94.105 23.825 94.430 ;
        RECT 18.675 93.935 19.225 94.105 ;
        RECT 23.275 93.935 23.825 94.105 ;
        RECT 24.005 93.865 24.375 94.205 ;
        RECT 24.555 94.105 24.725 94.430 ;
        RECT 24.555 93.925 25.485 94.105 ;
        RECT -291.460 93.245 -289.620 93.415 ;
        RECT 24.600 93.245 26.440 93.415 ;
        RECT -291.375 92.520 -291.085 93.245 ;
        RECT -290.915 92.445 -290.605 93.245 ;
        RECT -290.400 92.445 -289.705 93.075 ;
        RECT -291.375 90.695 -291.085 91.860 ;
        RECT -290.400 91.845 -290.230 92.445 ;
        RECT -290.060 92.005 -289.725 92.255 ;
        RECT -287.365 92.095 -287.035 93.075 ;
        RECT -285.505 92.095 -285.175 93.075 ;
        RECT -282.835 92.445 -282.140 93.075 ;
        RECT -290.915 90.695 -290.635 91.835 ;
        RECT -290.465 90.865 -290.135 91.845 ;
        RECT -289.965 90.695 -289.705 91.835 ;
        RECT -287.775 91.685 -287.440 91.935 ;
        RECT -287.270 91.495 -287.100 92.095 ;
        RECT -287.795 90.865 -287.100 91.495 ;
        RECT -285.440 91.495 -285.270 92.095 ;
        RECT -282.815 92.005 -282.480 92.255 ;
        RECT -285.100 91.685 -284.765 91.935 ;
        RECT -282.310 91.845 -282.140 92.445 ;
        RECT -280.480 92.445 -279.785 93.075 ;
        RECT -280.480 91.845 -280.310 92.445 ;
        RECT -280.140 92.005 -279.805 92.255 ;
        RECT -277.445 92.095 -277.115 93.075 ;
        RECT -275.585 92.095 -275.255 93.075 ;
        RECT -272.915 92.445 -272.220 93.075 ;
        RECT -285.440 90.865 -284.745 91.495 ;
        RECT -282.405 90.865 -282.075 91.845 ;
        RECT -280.545 90.865 -280.215 91.845 ;
        RECT -277.855 91.685 -277.520 91.935 ;
        RECT -277.350 91.495 -277.180 92.095 ;
        RECT -277.875 90.865 -277.180 91.495 ;
        RECT -275.520 91.495 -275.350 92.095 ;
        RECT -272.895 92.005 -272.560 92.255 ;
        RECT -275.180 91.685 -274.845 91.935 ;
        RECT -272.390 91.845 -272.220 92.445 ;
        RECT -270.560 92.445 -269.865 93.075 ;
        RECT -270.560 91.845 -270.390 92.445 ;
        RECT -270.220 92.005 -269.885 92.255 ;
        RECT -267.525 92.095 -267.195 93.075 ;
        RECT -265.665 92.095 -265.335 93.075 ;
        RECT -262.995 92.445 -262.300 93.075 ;
        RECT -275.520 90.865 -274.825 91.495 ;
        RECT -272.485 90.865 -272.155 91.845 ;
        RECT -270.625 90.865 -270.295 91.845 ;
        RECT -267.935 91.685 -267.600 91.935 ;
        RECT -267.430 91.495 -267.260 92.095 ;
        RECT -267.955 90.865 -267.260 91.495 ;
        RECT -265.600 91.495 -265.430 92.095 ;
        RECT -262.975 92.005 -262.640 92.255 ;
        RECT -265.260 91.685 -264.925 91.935 ;
        RECT -262.470 91.845 -262.300 92.445 ;
        RECT -260.640 92.445 -259.945 93.075 ;
        RECT -260.640 91.845 -260.470 92.445 ;
        RECT -260.300 92.005 -259.965 92.255 ;
        RECT -257.605 92.095 -257.275 93.075 ;
        RECT -255.745 92.095 -255.415 93.075 ;
        RECT -253.075 92.445 -252.380 93.075 ;
        RECT -265.600 90.865 -264.905 91.495 ;
        RECT -262.565 90.865 -262.235 91.845 ;
        RECT -260.705 90.865 -260.375 91.845 ;
        RECT -258.015 91.685 -257.680 91.935 ;
        RECT -257.510 91.495 -257.340 92.095 ;
        RECT -258.035 90.865 -257.340 91.495 ;
        RECT -255.680 91.495 -255.510 92.095 ;
        RECT -253.055 92.005 -252.720 92.255 ;
        RECT -255.340 91.685 -255.005 91.935 ;
        RECT -252.550 91.845 -252.380 92.445 ;
        RECT -250.720 92.445 -250.025 93.075 ;
        RECT -250.720 91.845 -250.550 92.445 ;
        RECT -250.380 92.005 -250.045 92.255 ;
        RECT -247.685 92.095 -247.355 93.075 ;
        RECT -245.825 92.095 -245.495 93.075 ;
        RECT -243.155 92.445 -242.460 93.075 ;
        RECT -255.680 90.865 -254.985 91.495 ;
        RECT -252.645 90.865 -252.315 91.845 ;
        RECT -250.785 90.865 -250.455 91.845 ;
        RECT -248.095 91.685 -247.760 91.935 ;
        RECT -247.590 91.495 -247.420 92.095 ;
        RECT -248.115 90.865 -247.420 91.495 ;
        RECT -245.760 91.495 -245.590 92.095 ;
        RECT -243.135 92.005 -242.800 92.255 ;
        RECT -245.420 91.685 -245.085 91.935 ;
        RECT -242.630 91.845 -242.460 92.445 ;
        RECT -240.800 92.445 -240.105 93.075 ;
        RECT -240.800 91.845 -240.630 92.445 ;
        RECT -240.460 92.005 -240.125 92.255 ;
        RECT -237.765 92.095 -237.435 93.075 ;
        RECT -235.905 92.095 -235.575 93.075 ;
        RECT -233.235 92.445 -232.540 93.075 ;
        RECT -245.760 90.865 -245.065 91.495 ;
        RECT -242.725 90.865 -242.395 91.845 ;
        RECT -240.865 90.865 -240.535 91.845 ;
        RECT -238.175 91.685 -237.840 91.935 ;
        RECT -237.670 91.495 -237.500 92.095 ;
        RECT -238.195 90.865 -237.500 91.495 ;
        RECT -235.840 91.495 -235.670 92.095 ;
        RECT -233.215 92.005 -232.880 92.255 ;
        RECT -235.500 91.685 -235.165 91.935 ;
        RECT -232.710 91.845 -232.540 92.445 ;
        RECT -230.880 92.445 -230.185 93.075 ;
        RECT -230.880 91.845 -230.710 92.445 ;
        RECT -230.540 92.005 -230.205 92.255 ;
        RECT -227.845 92.095 -227.515 93.075 ;
        RECT -225.985 92.095 -225.655 93.075 ;
        RECT -223.315 92.445 -222.620 93.075 ;
        RECT -235.840 90.865 -235.145 91.495 ;
        RECT -232.805 90.865 -232.475 91.845 ;
        RECT -230.945 90.865 -230.615 91.845 ;
        RECT -228.255 91.685 -227.920 91.935 ;
        RECT -227.750 91.495 -227.580 92.095 ;
        RECT -228.275 90.865 -227.580 91.495 ;
        RECT -225.920 91.495 -225.750 92.095 ;
        RECT -223.295 92.005 -222.960 92.255 ;
        RECT -225.580 91.685 -225.245 91.935 ;
        RECT -222.790 91.845 -222.620 92.445 ;
        RECT -220.960 92.445 -220.265 93.075 ;
        RECT -220.960 91.845 -220.790 92.445 ;
        RECT -220.620 92.005 -220.285 92.255 ;
        RECT -217.925 92.095 -217.595 93.075 ;
        RECT -216.065 92.095 -215.735 93.075 ;
        RECT -213.395 92.445 -212.700 93.075 ;
        RECT -225.920 90.865 -225.225 91.495 ;
        RECT -222.885 90.865 -222.555 91.845 ;
        RECT -221.025 90.865 -220.695 91.845 ;
        RECT -218.335 91.685 -218.000 91.935 ;
        RECT -217.830 91.495 -217.660 92.095 ;
        RECT -218.355 90.865 -217.660 91.495 ;
        RECT -216.000 91.495 -215.830 92.095 ;
        RECT -213.375 92.005 -213.040 92.255 ;
        RECT -215.660 91.685 -215.325 91.935 ;
        RECT -212.870 91.845 -212.700 92.445 ;
        RECT -211.040 92.445 -210.345 93.075 ;
        RECT -211.040 91.845 -210.870 92.445 ;
        RECT -210.700 92.005 -210.365 92.255 ;
        RECT -208.005 92.095 -207.675 93.075 ;
        RECT -206.145 92.095 -205.815 93.075 ;
        RECT -203.475 92.445 -202.780 93.075 ;
        RECT -216.000 90.865 -215.305 91.495 ;
        RECT -212.965 90.865 -212.635 91.845 ;
        RECT -211.105 90.865 -210.775 91.845 ;
        RECT -208.415 91.685 -208.080 91.935 ;
        RECT -207.910 91.495 -207.740 92.095 ;
        RECT -208.435 90.865 -207.740 91.495 ;
        RECT -206.080 91.495 -205.910 92.095 ;
        RECT -203.455 92.005 -203.120 92.255 ;
        RECT -205.740 91.685 -205.405 91.935 ;
        RECT -202.950 91.845 -202.780 92.445 ;
        RECT -201.120 92.445 -200.425 93.075 ;
        RECT -201.120 91.845 -200.950 92.445 ;
        RECT -200.780 92.005 -200.445 92.255 ;
        RECT -198.085 92.095 -197.755 93.075 ;
        RECT -196.225 92.095 -195.895 93.075 ;
        RECT -193.555 92.445 -192.860 93.075 ;
        RECT -206.080 90.865 -205.385 91.495 ;
        RECT -203.045 90.865 -202.715 91.845 ;
        RECT -201.185 90.865 -200.855 91.845 ;
        RECT -198.495 91.685 -198.160 91.935 ;
        RECT -197.990 91.495 -197.820 92.095 ;
        RECT -198.515 90.865 -197.820 91.495 ;
        RECT -196.160 91.495 -195.990 92.095 ;
        RECT -193.535 92.005 -193.200 92.255 ;
        RECT -195.820 91.685 -195.485 91.935 ;
        RECT -193.030 91.845 -192.860 92.445 ;
        RECT -191.200 92.445 -190.505 93.075 ;
        RECT -191.200 91.845 -191.030 92.445 ;
        RECT -190.860 92.005 -190.525 92.255 ;
        RECT -188.165 92.095 -187.835 93.075 ;
        RECT -186.305 92.095 -185.975 93.075 ;
        RECT -183.635 92.445 -182.940 93.075 ;
        RECT -196.160 90.865 -195.465 91.495 ;
        RECT -193.125 90.865 -192.795 91.845 ;
        RECT -191.265 90.865 -190.935 91.845 ;
        RECT -188.575 91.685 -188.240 91.935 ;
        RECT -188.070 91.495 -187.900 92.095 ;
        RECT -188.595 90.865 -187.900 91.495 ;
        RECT -186.240 91.495 -186.070 92.095 ;
        RECT -183.615 92.005 -183.280 92.255 ;
        RECT -185.900 91.685 -185.565 91.935 ;
        RECT -183.110 91.845 -182.940 92.445 ;
        RECT -181.280 92.445 -180.585 93.075 ;
        RECT -181.280 91.845 -181.110 92.445 ;
        RECT -180.940 92.005 -180.605 92.255 ;
        RECT -178.245 92.095 -177.915 93.075 ;
        RECT -176.385 92.095 -176.055 93.075 ;
        RECT -173.715 92.445 -173.020 93.075 ;
        RECT -186.240 90.865 -185.545 91.495 ;
        RECT -183.205 90.865 -182.875 91.845 ;
        RECT -181.345 90.865 -181.015 91.845 ;
        RECT -178.655 91.685 -178.320 91.935 ;
        RECT -178.150 91.495 -177.980 92.095 ;
        RECT -178.675 90.865 -177.980 91.495 ;
        RECT -176.320 91.495 -176.150 92.095 ;
        RECT -173.695 92.005 -173.360 92.255 ;
        RECT -175.980 91.685 -175.645 91.935 ;
        RECT -173.190 91.845 -173.020 92.445 ;
        RECT -171.360 92.445 -170.665 93.075 ;
        RECT -171.360 91.845 -171.190 92.445 ;
        RECT -171.020 92.005 -170.685 92.255 ;
        RECT -168.325 92.095 -167.995 93.075 ;
        RECT -166.465 92.095 -166.135 93.075 ;
        RECT -163.795 92.445 -163.100 93.075 ;
        RECT -176.320 90.865 -175.625 91.495 ;
        RECT -173.285 90.865 -172.955 91.845 ;
        RECT -171.425 90.865 -171.095 91.845 ;
        RECT -168.735 91.685 -168.400 91.935 ;
        RECT -168.230 91.495 -168.060 92.095 ;
        RECT -168.755 90.865 -168.060 91.495 ;
        RECT -166.400 91.495 -166.230 92.095 ;
        RECT -163.775 92.005 -163.440 92.255 ;
        RECT -166.060 91.685 -165.725 91.935 ;
        RECT -163.270 91.845 -163.100 92.445 ;
        RECT -161.440 92.445 -160.745 93.075 ;
        RECT -161.440 91.845 -161.270 92.445 ;
        RECT -161.100 92.005 -160.765 92.255 ;
        RECT -158.405 92.095 -158.075 93.075 ;
        RECT -156.545 92.095 -156.215 93.075 ;
        RECT -153.875 92.445 -153.180 93.075 ;
        RECT -166.400 90.865 -165.705 91.495 ;
        RECT -163.365 90.865 -163.035 91.845 ;
        RECT -161.505 90.865 -161.175 91.845 ;
        RECT -158.815 91.685 -158.480 91.935 ;
        RECT -158.310 91.495 -158.140 92.095 ;
        RECT -158.835 90.865 -158.140 91.495 ;
        RECT -156.480 91.495 -156.310 92.095 ;
        RECT -153.855 92.005 -153.520 92.255 ;
        RECT -156.140 91.685 -155.805 91.935 ;
        RECT -153.350 91.845 -153.180 92.445 ;
        RECT -151.520 92.445 -150.825 93.075 ;
        RECT -151.520 91.845 -151.350 92.445 ;
        RECT -151.180 92.005 -150.845 92.255 ;
        RECT -148.485 92.095 -148.155 93.075 ;
        RECT -146.625 92.095 -146.295 93.075 ;
        RECT -143.955 92.445 -143.260 93.075 ;
        RECT -156.480 90.865 -155.785 91.495 ;
        RECT -153.445 90.865 -153.115 91.845 ;
        RECT -151.585 90.865 -151.255 91.845 ;
        RECT -148.895 91.685 -148.560 91.935 ;
        RECT -148.390 91.495 -148.220 92.095 ;
        RECT -148.915 90.865 -148.220 91.495 ;
        RECT -146.560 91.495 -146.390 92.095 ;
        RECT -143.935 92.005 -143.600 92.255 ;
        RECT -146.220 91.685 -145.885 91.935 ;
        RECT -143.430 91.845 -143.260 92.445 ;
        RECT -141.600 92.445 -140.905 93.075 ;
        RECT -141.600 91.845 -141.430 92.445 ;
        RECT -141.260 92.005 -140.925 92.255 ;
        RECT -138.565 92.095 -138.235 93.075 ;
        RECT -136.705 92.095 -136.375 93.075 ;
        RECT -134.035 92.445 -133.340 93.075 ;
        RECT -146.560 90.865 -145.865 91.495 ;
        RECT -143.525 90.865 -143.195 91.845 ;
        RECT -141.665 90.865 -141.335 91.845 ;
        RECT -138.975 91.685 -138.640 91.935 ;
        RECT -138.470 91.495 -138.300 92.095 ;
        RECT -138.995 90.865 -138.300 91.495 ;
        RECT -136.640 91.495 -136.470 92.095 ;
        RECT -134.015 92.005 -133.680 92.255 ;
        RECT -136.300 91.685 -135.965 91.935 ;
        RECT -133.510 91.845 -133.340 92.445 ;
        RECT -131.680 92.445 -130.985 93.075 ;
        RECT -131.680 91.845 -131.510 92.445 ;
        RECT -131.340 92.005 -131.005 92.255 ;
        RECT -128.645 92.095 -128.315 93.075 ;
        RECT -126.785 92.095 -126.455 93.075 ;
        RECT -124.115 92.445 -123.420 93.075 ;
        RECT -136.640 90.865 -135.945 91.495 ;
        RECT -133.605 90.865 -133.275 91.845 ;
        RECT -131.745 90.865 -131.415 91.845 ;
        RECT -129.055 91.685 -128.720 91.935 ;
        RECT -128.550 91.495 -128.380 92.095 ;
        RECT -129.075 90.865 -128.380 91.495 ;
        RECT -126.720 91.495 -126.550 92.095 ;
        RECT -124.095 92.005 -123.760 92.255 ;
        RECT -126.380 91.685 -126.045 91.935 ;
        RECT -123.590 91.845 -123.420 92.445 ;
        RECT -121.760 92.445 -121.065 93.075 ;
        RECT -121.760 91.845 -121.590 92.445 ;
        RECT -121.420 92.005 -121.085 92.255 ;
        RECT -118.725 92.095 -118.395 93.075 ;
        RECT -116.865 92.095 -116.535 93.075 ;
        RECT -114.195 92.445 -113.500 93.075 ;
        RECT -126.720 90.865 -126.025 91.495 ;
        RECT -123.685 90.865 -123.355 91.845 ;
        RECT -121.825 90.865 -121.495 91.845 ;
        RECT -119.135 91.685 -118.800 91.935 ;
        RECT -118.630 91.495 -118.460 92.095 ;
        RECT -119.155 90.865 -118.460 91.495 ;
        RECT -116.800 91.495 -116.630 92.095 ;
        RECT -114.175 92.005 -113.840 92.255 ;
        RECT -116.460 91.685 -116.125 91.935 ;
        RECT -113.670 91.845 -113.500 92.445 ;
        RECT -111.840 92.445 -111.145 93.075 ;
        RECT -111.840 91.845 -111.670 92.445 ;
        RECT -111.500 92.005 -111.165 92.255 ;
        RECT -108.805 92.095 -108.475 93.075 ;
        RECT -106.945 92.095 -106.615 93.075 ;
        RECT -104.275 92.445 -103.580 93.075 ;
        RECT -116.800 90.865 -116.105 91.495 ;
        RECT -113.765 90.865 -113.435 91.845 ;
        RECT -111.905 90.865 -111.575 91.845 ;
        RECT -109.215 91.685 -108.880 91.935 ;
        RECT -108.710 91.495 -108.540 92.095 ;
        RECT -109.235 90.865 -108.540 91.495 ;
        RECT -106.880 91.495 -106.710 92.095 ;
        RECT -104.255 92.005 -103.920 92.255 ;
        RECT -106.540 91.685 -106.205 91.935 ;
        RECT -103.750 91.845 -103.580 92.445 ;
        RECT -101.920 92.445 -101.225 93.075 ;
        RECT -101.920 91.845 -101.750 92.445 ;
        RECT -101.580 92.005 -101.245 92.255 ;
        RECT -98.885 92.095 -98.555 93.075 ;
        RECT -97.025 92.095 -96.695 93.075 ;
        RECT -94.355 92.445 -93.660 93.075 ;
        RECT -106.880 90.865 -106.185 91.495 ;
        RECT -103.845 90.865 -103.515 91.845 ;
        RECT -101.985 90.865 -101.655 91.845 ;
        RECT -99.295 91.685 -98.960 91.935 ;
        RECT -98.790 91.495 -98.620 92.095 ;
        RECT -99.315 90.865 -98.620 91.495 ;
        RECT -96.960 91.495 -96.790 92.095 ;
        RECT -94.335 92.005 -94.000 92.255 ;
        RECT -96.620 91.685 -96.285 91.935 ;
        RECT -93.830 91.845 -93.660 92.445 ;
        RECT -92.000 92.445 -91.305 93.075 ;
        RECT -92.000 91.845 -91.830 92.445 ;
        RECT -91.660 92.005 -91.325 92.255 ;
        RECT -88.965 92.095 -88.635 93.075 ;
        RECT -87.105 92.095 -86.775 93.075 ;
        RECT -84.435 92.445 -83.740 93.075 ;
        RECT -96.960 90.865 -96.265 91.495 ;
        RECT -93.925 90.865 -93.595 91.845 ;
        RECT -92.065 90.865 -91.735 91.845 ;
        RECT -89.375 91.685 -89.040 91.935 ;
        RECT -88.870 91.495 -88.700 92.095 ;
        RECT -89.395 90.865 -88.700 91.495 ;
        RECT -87.040 91.495 -86.870 92.095 ;
        RECT -84.415 92.005 -84.080 92.255 ;
        RECT -86.700 91.685 -86.365 91.935 ;
        RECT -83.910 91.845 -83.740 92.445 ;
        RECT -82.080 92.445 -81.385 93.075 ;
        RECT -82.080 91.845 -81.910 92.445 ;
        RECT -81.740 92.005 -81.405 92.255 ;
        RECT -79.045 92.095 -78.715 93.075 ;
        RECT -77.185 92.095 -76.855 93.075 ;
        RECT -74.515 92.445 -73.820 93.075 ;
        RECT -87.040 90.865 -86.345 91.495 ;
        RECT -84.005 90.865 -83.675 91.845 ;
        RECT -82.145 90.865 -81.815 91.845 ;
        RECT -79.455 91.685 -79.120 91.935 ;
        RECT -78.950 91.495 -78.780 92.095 ;
        RECT -79.475 90.865 -78.780 91.495 ;
        RECT -77.120 91.495 -76.950 92.095 ;
        RECT -74.495 92.005 -74.160 92.255 ;
        RECT -76.780 91.685 -76.445 91.935 ;
        RECT -73.990 91.845 -73.820 92.445 ;
        RECT -72.160 92.445 -71.465 93.075 ;
        RECT -72.160 91.845 -71.990 92.445 ;
        RECT -71.820 92.005 -71.485 92.255 ;
        RECT -69.125 92.095 -68.795 93.075 ;
        RECT -67.265 92.095 -66.935 93.075 ;
        RECT -64.595 92.445 -63.900 93.075 ;
        RECT -77.120 90.865 -76.425 91.495 ;
        RECT -74.085 90.865 -73.755 91.845 ;
        RECT -72.225 90.865 -71.895 91.845 ;
        RECT -69.535 91.685 -69.200 91.935 ;
        RECT -69.030 91.495 -68.860 92.095 ;
        RECT -69.555 90.865 -68.860 91.495 ;
        RECT -67.200 91.495 -67.030 92.095 ;
        RECT -64.575 92.005 -64.240 92.255 ;
        RECT -66.860 91.685 -66.525 91.935 ;
        RECT -64.070 91.845 -63.900 92.445 ;
        RECT -62.240 92.445 -61.545 93.075 ;
        RECT -62.240 91.845 -62.070 92.445 ;
        RECT -61.900 92.005 -61.565 92.255 ;
        RECT -59.205 92.095 -58.875 93.075 ;
        RECT -57.345 92.095 -57.015 93.075 ;
        RECT -54.675 92.445 -53.980 93.075 ;
        RECT -67.200 90.865 -66.505 91.495 ;
        RECT -64.165 90.865 -63.835 91.845 ;
        RECT -62.305 90.865 -61.975 91.845 ;
        RECT -59.615 91.685 -59.280 91.935 ;
        RECT -59.110 91.495 -58.940 92.095 ;
        RECT -59.635 90.865 -58.940 91.495 ;
        RECT -57.280 91.495 -57.110 92.095 ;
        RECT -54.655 92.005 -54.320 92.255 ;
        RECT -56.940 91.685 -56.605 91.935 ;
        RECT -54.150 91.845 -53.980 92.445 ;
        RECT -52.320 92.445 -51.625 93.075 ;
        RECT -52.320 91.845 -52.150 92.445 ;
        RECT -51.980 92.005 -51.645 92.255 ;
        RECT -49.285 92.095 -48.955 93.075 ;
        RECT -47.425 92.095 -47.095 93.075 ;
        RECT -44.755 92.445 -44.060 93.075 ;
        RECT -57.280 90.865 -56.585 91.495 ;
        RECT -54.245 90.865 -53.915 91.845 ;
        RECT -52.385 90.865 -52.055 91.845 ;
        RECT -49.695 91.685 -49.360 91.935 ;
        RECT -49.190 91.495 -49.020 92.095 ;
        RECT -49.715 90.865 -49.020 91.495 ;
        RECT -47.360 91.495 -47.190 92.095 ;
        RECT -44.735 92.005 -44.400 92.255 ;
        RECT -47.020 91.685 -46.685 91.935 ;
        RECT -44.230 91.845 -44.060 92.445 ;
        RECT -42.400 92.445 -41.705 93.075 ;
        RECT -42.400 91.845 -42.230 92.445 ;
        RECT -42.060 92.005 -41.725 92.255 ;
        RECT -39.365 92.095 -39.035 93.075 ;
        RECT -37.505 92.095 -37.175 93.075 ;
        RECT -34.835 92.445 -34.140 93.075 ;
        RECT -47.360 90.865 -46.665 91.495 ;
        RECT -44.325 90.865 -43.995 91.845 ;
        RECT -42.465 90.865 -42.135 91.845 ;
        RECT -39.775 91.685 -39.440 91.935 ;
        RECT -39.270 91.495 -39.100 92.095 ;
        RECT -39.795 90.865 -39.100 91.495 ;
        RECT -37.440 91.495 -37.270 92.095 ;
        RECT -34.815 92.005 -34.480 92.255 ;
        RECT -37.100 91.685 -36.765 91.935 ;
        RECT -34.310 91.845 -34.140 92.445 ;
        RECT -32.480 92.445 -31.785 93.075 ;
        RECT -32.480 91.845 -32.310 92.445 ;
        RECT -32.140 92.005 -31.805 92.255 ;
        RECT -29.445 92.095 -29.115 93.075 ;
        RECT -27.585 92.095 -27.255 93.075 ;
        RECT -24.915 92.445 -24.220 93.075 ;
        RECT -37.440 90.865 -36.745 91.495 ;
        RECT -34.405 90.865 -34.075 91.845 ;
        RECT -32.545 90.865 -32.215 91.845 ;
        RECT -29.855 91.685 -29.520 91.935 ;
        RECT -29.350 91.495 -29.180 92.095 ;
        RECT -29.875 90.865 -29.180 91.495 ;
        RECT -27.520 91.495 -27.350 92.095 ;
        RECT -24.895 92.005 -24.560 92.255 ;
        RECT -27.180 91.685 -26.845 91.935 ;
        RECT -24.390 91.845 -24.220 92.445 ;
        RECT -22.560 92.445 -21.865 93.075 ;
        RECT -22.560 91.845 -22.390 92.445 ;
        RECT -22.220 92.005 -21.885 92.255 ;
        RECT -19.525 92.095 -19.195 93.075 ;
        RECT -17.665 92.095 -17.335 93.075 ;
        RECT -14.995 92.445 -14.300 93.075 ;
        RECT -27.520 90.865 -26.825 91.495 ;
        RECT -24.485 90.865 -24.155 91.845 ;
        RECT -22.625 90.865 -22.295 91.845 ;
        RECT -19.935 91.685 -19.600 91.935 ;
        RECT -19.430 91.495 -19.260 92.095 ;
        RECT -19.955 90.865 -19.260 91.495 ;
        RECT -17.600 91.495 -17.430 92.095 ;
        RECT -14.975 92.005 -14.640 92.255 ;
        RECT -17.260 91.685 -16.925 91.935 ;
        RECT -14.470 91.845 -14.300 92.445 ;
        RECT -12.640 92.445 -11.945 93.075 ;
        RECT -12.640 91.845 -12.470 92.445 ;
        RECT -12.300 92.005 -11.965 92.255 ;
        RECT -9.605 92.095 -9.275 93.075 ;
        RECT -7.745 92.095 -7.415 93.075 ;
        RECT -5.075 92.445 -4.380 93.075 ;
        RECT -17.600 90.865 -16.905 91.495 ;
        RECT -14.565 90.865 -14.235 91.845 ;
        RECT -12.705 90.865 -12.375 91.845 ;
        RECT -10.015 91.685 -9.680 91.935 ;
        RECT -9.510 91.495 -9.340 92.095 ;
        RECT -10.035 90.865 -9.340 91.495 ;
        RECT -7.680 91.495 -7.510 92.095 ;
        RECT -5.055 92.005 -4.720 92.255 ;
        RECT -7.340 91.685 -7.005 91.935 ;
        RECT -4.550 91.845 -4.380 92.445 ;
        RECT -2.720 92.445 -2.025 93.075 ;
        RECT -2.720 91.845 -2.550 92.445 ;
        RECT -2.380 92.005 -2.045 92.255 ;
        RECT 0.315 92.095 0.645 93.075 ;
        RECT 2.175 92.095 2.505 93.075 ;
        RECT 4.845 92.445 5.540 93.075 ;
        RECT -7.680 90.865 -6.985 91.495 ;
        RECT -4.645 90.865 -4.315 91.845 ;
        RECT -2.785 90.865 -2.455 91.845 ;
        RECT -0.095 91.685 0.240 91.935 ;
        RECT 0.410 91.495 0.580 92.095 ;
        RECT -0.115 90.865 0.580 91.495 ;
        RECT 2.240 91.495 2.410 92.095 ;
        RECT 4.865 92.005 5.200 92.255 ;
        RECT 2.580 91.685 2.915 91.935 ;
        RECT 5.370 91.845 5.540 92.445 ;
        RECT 7.200 92.445 7.895 93.075 ;
        RECT 7.200 91.845 7.370 92.445 ;
        RECT 7.540 92.005 7.875 92.255 ;
        RECT 10.235 92.095 10.565 93.075 ;
        RECT 12.095 92.095 12.425 93.075 ;
        RECT 14.765 92.445 15.460 93.075 ;
        RECT 2.240 90.865 2.935 91.495 ;
        RECT 5.275 90.865 5.605 91.845 ;
        RECT 7.135 90.865 7.465 91.845 ;
        RECT 9.825 91.685 10.160 91.935 ;
        RECT 10.330 91.495 10.500 92.095 ;
        RECT 9.805 90.865 10.500 91.495 ;
        RECT 12.160 91.495 12.330 92.095 ;
        RECT 14.785 92.005 15.120 92.255 ;
        RECT 12.500 91.685 12.835 91.935 ;
        RECT 15.290 91.845 15.460 92.445 ;
        RECT 17.120 92.445 17.815 93.075 ;
        RECT 17.120 91.845 17.290 92.445 ;
        RECT 17.460 92.005 17.795 92.255 ;
        RECT 20.155 92.095 20.485 93.075 ;
        RECT 22.015 92.095 22.345 93.075 ;
        RECT 24.685 92.445 25.380 93.075 ;
        RECT 25.585 92.445 25.895 93.245 ;
        RECT 26.065 92.520 26.355 93.245 ;
        RECT 12.160 90.865 12.855 91.495 ;
        RECT 15.195 90.865 15.525 91.845 ;
        RECT 17.055 90.865 17.385 91.845 ;
        RECT 19.745 91.685 20.080 91.935 ;
        RECT 20.250 91.495 20.420 92.095 ;
        RECT 19.725 90.865 20.420 91.495 ;
        RECT 22.080 91.495 22.250 92.095 ;
        RECT 24.705 92.005 25.040 92.255 ;
        RECT 22.420 91.685 22.755 91.935 ;
        RECT 25.210 91.845 25.380 92.445 ;
        RECT 22.080 90.865 22.775 91.495 ;
        RECT 25.115 90.865 25.445 91.845 ;
        RECT -291.460 90.525 -289.620 90.695 ;
        RECT -290.075 89.140 -289.785 89.850 ;
        RECT -289.545 89.655 -289.375 90.180 ;
        RECT -289.205 89.835 -288.655 90.005 ;
        RECT -289.545 89.325 -288.995 89.655 ;
        RECT -288.825 89.510 -288.655 89.835 ;
        RECT -288.475 89.735 -288.105 90.075 ;
        RECT -287.925 89.835 -286.995 90.015 ;
        RECT -285.545 89.835 -284.615 90.015 ;
        RECT -287.925 89.510 -287.755 89.835 ;
        RECT -288.825 89.340 -287.755 89.510 ;
        RECT -284.785 89.510 -284.615 89.835 ;
        RECT -284.435 89.735 -284.065 90.075 ;
        RECT -283.885 89.835 -283.335 90.005 ;
        RECT -279.285 89.835 -278.735 90.005 ;
        RECT -283.885 89.510 -283.715 89.835 ;
        RECT -284.785 89.340 -283.715 89.510 ;
        RECT -278.905 89.510 -278.735 89.835 ;
        RECT -278.555 89.735 -278.185 90.075 ;
        RECT -278.005 89.835 -277.075 90.015 ;
        RECT -275.625 89.835 -274.695 90.015 ;
        RECT -278.005 89.510 -277.835 89.835 ;
        RECT -278.905 89.340 -277.835 89.510 ;
        RECT -274.865 89.510 -274.695 89.835 ;
        RECT -274.515 89.735 -274.145 90.075 ;
        RECT -273.965 89.835 -273.415 90.005 ;
        RECT -269.365 89.835 -268.815 90.005 ;
        RECT -273.965 89.510 -273.795 89.835 ;
        RECT -274.865 89.340 -273.795 89.510 ;
        RECT -268.985 89.510 -268.815 89.835 ;
        RECT -268.635 89.735 -268.265 90.075 ;
        RECT -268.085 89.835 -267.155 90.015 ;
        RECT -265.705 89.835 -264.775 90.015 ;
        RECT -268.085 89.510 -267.915 89.835 ;
        RECT -268.985 89.340 -267.915 89.510 ;
        RECT -264.945 89.510 -264.775 89.835 ;
        RECT -264.595 89.735 -264.225 90.075 ;
        RECT -264.045 89.835 -263.495 90.005 ;
        RECT -259.445 89.835 -258.895 90.005 ;
        RECT -264.045 89.510 -263.875 89.835 ;
        RECT -264.945 89.340 -263.875 89.510 ;
        RECT -259.065 89.510 -258.895 89.835 ;
        RECT -258.715 89.735 -258.345 90.075 ;
        RECT -258.165 89.835 -257.235 90.015 ;
        RECT -255.785 89.835 -254.855 90.015 ;
        RECT -258.165 89.510 -257.995 89.835 ;
        RECT -259.065 89.340 -257.995 89.510 ;
        RECT -255.025 89.510 -254.855 89.835 ;
        RECT -254.675 89.735 -254.305 90.075 ;
        RECT -254.125 89.835 -253.575 90.005 ;
        RECT -249.525 89.835 -248.975 90.005 ;
        RECT -254.125 89.510 -253.955 89.835 ;
        RECT -255.025 89.340 -253.955 89.510 ;
        RECT -249.145 89.510 -248.975 89.835 ;
        RECT -248.795 89.735 -248.425 90.075 ;
        RECT -248.245 89.835 -247.315 90.015 ;
        RECT -245.865 89.835 -244.935 90.015 ;
        RECT -248.245 89.510 -248.075 89.835 ;
        RECT -249.145 89.340 -248.075 89.510 ;
        RECT -245.105 89.510 -244.935 89.835 ;
        RECT -244.755 89.735 -244.385 90.075 ;
        RECT -244.205 89.835 -243.655 90.005 ;
        RECT -239.605 89.835 -239.055 90.005 ;
        RECT -244.205 89.510 -244.035 89.835 ;
        RECT -245.105 89.340 -244.035 89.510 ;
        RECT -239.225 89.510 -239.055 89.835 ;
        RECT -238.875 89.735 -238.505 90.075 ;
        RECT -238.325 89.835 -237.395 90.015 ;
        RECT -235.945 89.835 -235.015 90.015 ;
        RECT -238.325 89.510 -238.155 89.835 ;
        RECT -239.225 89.340 -238.155 89.510 ;
        RECT -235.185 89.510 -235.015 89.835 ;
        RECT -234.835 89.735 -234.465 90.075 ;
        RECT -234.285 89.835 -233.735 90.005 ;
        RECT -229.685 89.835 -229.135 90.005 ;
        RECT -234.285 89.510 -234.115 89.835 ;
        RECT -235.185 89.340 -234.115 89.510 ;
        RECT -229.305 89.510 -229.135 89.835 ;
        RECT -228.955 89.735 -228.585 90.075 ;
        RECT -228.405 89.835 -227.475 90.015 ;
        RECT -226.025 89.835 -225.095 90.015 ;
        RECT -228.405 89.510 -228.235 89.835 ;
        RECT -229.305 89.340 -228.235 89.510 ;
        RECT -225.265 89.510 -225.095 89.835 ;
        RECT -224.915 89.735 -224.545 90.075 ;
        RECT -224.365 89.835 -223.815 90.005 ;
        RECT -219.765 89.835 -219.215 90.005 ;
        RECT -224.365 89.510 -224.195 89.835 ;
        RECT -225.265 89.340 -224.195 89.510 ;
        RECT -219.385 89.510 -219.215 89.835 ;
        RECT -219.035 89.735 -218.665 90.075 ;
        RECT -218.485 89.835 -217.555 90.015 ;
        RECT -216.105 89.835 -215.175 90.015 ;
        RECT -218.485 89.510 -218.315 89.835 ;
        RECT -219.385 89.340 -218.315 89.510 ;
        RECT -215.345 89.510 -215.175 89.835 ;
        RECT -214.995 89.735 -214.625 90.075 ;
        RECT -214.445 89.835 -213.895 90.005 ;
        RECT -209.845 89.835 -209.295 90.005 ;
        RECT -214.445 89.510 -214.275 89.835 ;
        RECT -215.345 89.340 -214.275 89.510 ;
        RECT -209.465 89.510 -209.295 89.835 ;
        RECT -209.115 89.735 -208.745 90.075 ;
        RECT -208.565 89.835 -207.635 90.015 ;
        RECT -206.185 89.835 -205.255 90.015 ;
        RECT -208.565 89.510 -208.395 89.835 ;
        RECT -209.465 89.340 -208.395 89.510 ;
        RECT -205.425 89.510 -205.255 89.835 ;
        RECT -205.075 89.735 -204.705 90.075 ;
        RECT -204.525 89.835 -203.975 90.005 ;
        RECT -199.925 89.835 -199.375 90.005 ;
        RECT -204.525 89.510 -204.355 89.835 ;
        RECT -205.425 89.340 -204.355 89.510 ;
        RECT -199.545 89.510 -199.375 89.835 ;
        RECT -199.195 89.735 -198.825 90.075 ;
        RECT -198.645 89.835 -197.715 90.015 ;
        RECT -196.265 89.835 -195.335 90.015 ;
        RECT -198.645 89.510 -198.475 89.835 ;
        RECT -199.545 89.340 -198.475 89.510 ;
        RECT -195.505 89.510 -195.335 89.835 ;
        RECT -195.155 89.735 -194.785 90.075 ;
        RECT -194.605 89.835 -194.055 90.005 ;
        RECT -190.005 89.835 -189.455 90.005 ;
        RECT -194.605 89.510 -194.435 89.835 ;
        RECT -195.505 89.340 -194.435 89.510 ;
        RECT -189.625 89.510 -189.455 89.835 ;
        RECT -189.275 89.735 -188.905 90.075 ;
        RECT -188.725 89.835 -187.795 90.015 ;
        RECT -186.345 89.835 -185.415 90.015 ;
        RECT -188.725 89.510 -188.555 89.835 ;
        RECT -189.625 89.340 -188.555 89.510 ;
        RECT -185.585 89.510 -185.415 89.835 ;
        RECT -185.235 89.735 -184.865 90.075 ;
        RECT -184.685 89.835 -184.135 90.005 ;
        RECT -180.085 89.835 -179.535 90.005 ;
        RECT -184.685 89.510 -184.515 89.835 ;
        RECT -185.585 89.340 -184.515 89.510 ;
        RECT -179.705 89.510 -179.535 89.835 ;
        RECT -179.355 89.735 -178.985 90.075 ;
        RECT -178.805 89.835 -177.875 90.015 ;
        RECT -176.425 89.835 -175.495 90.015 ;
        RECT -178.805 89.510 -178.635 89.835 ;
        RECT -179.705 89.340 -178.635 89.510 ;
        RECT -175.665 89.510 -175.495 89.835 ;
        RECT -175.315 89.735 -174.945 90.075 ;
        RECT -174.765 89.835 -174.215 90.005 ;
        RECT -170.165 89.835 -169.615 90.005 ;
        RECT -174.765 89.510 -174.595 89.835 ;
        RECT -175.665 89.340 -174.595 89.510 ;
        RECT -169.785 89.510 -169.615 89.835 ;
        RECT -169.435 89.735 -169.065 90.075 ;
        RECT -168.885 89.835 -167.955 90.015 ;
        RECT -166.505 89.835 -165.575 90.015 ;
        RECT -168.885 89.510 -168.715 89.835 ;
        RECT -169.785 89.340 -168.715 89.510 ;
        RECT -165.745 89.510 -165.575 89.835 ;
        RECT -165.395 89.735 -165.025 90.075 ;
        RECT -164.845 89.835 -164.295 90.005 ;
        RECT -160.245 89.835 -159.695 90.005 ;
        RECT -164.845 89.510 -164.675 89.835 ;
        RECT -165.745 89.340 -164.675 89.510 ;
        RECT -159.865 89.510 -159.695 89.835 ;
        RECT -159.515 89.735 -159.145 90.075 ;
        RECT -158.965 89.835 -158.035 90.015 ;
        RECT -156.585 89.835 -155.655 90.015 ;
        RECT -158.965 89.510 -158.795 89.835 ;
        RECT -159.865 89.340 -158.795 89.510 ;
        RECT -155.825 89.510 -155.655 89.835 ;
        RECT -155.475 89.735 -155.105 90.075 ;
        RECT -154.925 89.835 -154.375 90.005 ;
        RECT -150.325 89.835 -149.775 90.005 ;
        RECT -154.925 89.510 -154.755 89.835 ;
        RECT -155.825 89.340 -154.755 89.510 ;
        RECT -149.945 89.510 -149.775 89.835 ;
        RECT -149.595 89.735 -149.225 90.075 ;
        RECT -149.045 89.835 -148.115 90.015 ;
        RECT -146.665 89.835 -145.735 90.015 ;
        RECT -149.045 89.510 -148.875 89.835 ;
        RECT -149.945 89.340 -148.875 89.510 ;
        RECT -145.905 89.510 -145.735 89.835 ;
        RECT -145.555 89.735 -145.185 90.075 ;
        RECT -145.005 89.835 -144.455 90.005 ;
        RECT -140.405 89.835 -139.855 90.005 ;
        RECT -145.005 89.510 -144.835 89.835 ;
        RECT -145.905 89.340 -144.835 89.510 ;
        RECT -140.025 89.510 -139.855 89.835 ;
        RECT -139.675 89.735 -139.305 90.075 ;
        RECT -139.125 89.835 -138.195 90.015 ;
        RECT -136.745 89.835 -135.815 90.015 ;
        RECT -139.125 89.510 -138.955 89.835 ;
        RECT -140.025 89.340 -138.955 89.510 ;
        RECT -135.985 89.510 -135.815 89.835 ;
        RECT -135.635 89.735 -135.265 90.075 ;
        RECT -135.085 89.835 -134.535 90.005 ;
        RECT -130.485 89.835 -129.935 90.005 ;
        RECT -135.085 89.510 -134.915 89.835 ;
        RECT -135.985 89.340 -134.915 89.510 ;
        RECT -130.105 89.510 -129.935 89.835 ;
        RECT -129.755 89.735 -129.385 90.075 ;
        RECT -129.205 89.835 -128.275 90.015 ;
        RECT -126.825 89.835 -125.895 90.015 ;
        RECT -129.205 89.510 -129.035 89.835 ;
        RECT -130.105 89.340 -129.035 89.510 ;
        RECT -126.065 89.510 -125.895 89.835 ;
        RECT -125.715 89.735 -125.345 90.075 ;
        RECT -125.165 89.835 -124.615 90.005 ;
        RECT -120.565 89.835 -120.015 90.005 ;
        RECT -125.165 89.510 -124.995 89.835 ;
        RECT -126.065 89.340 -124.995 89.510 ;
        RECT -120.185 89.510 -120.015 89.835 ;
        RECT -119.835 89.735 -119.465 90.075 ;
        RECT -119.285 89.835 -118.355 90.015 ;
        RECT -116.905 89.835 -115.975 90.015 ;
        RECT -119.285 89.510 -119.115 89.835 ;
        RECT -120.185 89.340 -119.115 89.510 ;
        RECT -116.145 89.510 -115.975 89.835 ;
        RECT -115.795 89.735 -115.425 90.075 ;
        RECT -115.245 89.835 -114.695 90.005 ;
        RECT -110.645 89.835 -110.095 90.005 ;
        RECT -115.245 89.510 -115.075 89.835 ;
        RECT -116.145 89.340 -115.075 89.510 ;
        RECT -110.265 89.510 -110.095 89.835 ;
        RECT -109.915 89.735 -109.545 90.075 ;
        RECT -109.365 89.835 -108.435 90.015 ;
        RECT -106.985 89.835 -106.055 90.015 ;
        RECT -109.365 89.510 -109.195 89.835 ;
        RECT -110.265 89.340 -109.195 89.510 ;
        RECT -106.225 89.510 -106.055 89.835 ;
        RECT -105.875 89.735 -105.505 90.075 ;
        RECT -105.325 89.835 -104.775 90.005 ;
        RECT -100.725 89.835 -100.175 90.005 ;
        RECT -105.325 89.510 -105.155 89.835 ;
        RECT -106.225 89.340 -105.155 89.510 ;
        RECT -100.345 89.510 -100.175 89.835 ;
        RECT -99.995 89.735 -99.625 90.075 ;
        RECT -99.445 89.835 -98.515 90.015 ;
        RECT -97.065 89.835 -96.135 90.015 ;
        RECT -99.445 89.510 -99.275 89.835 ;
        RECT -100.345 89.340 -99.275 89.510 ;
        RECT -96.305 89.510 -96.135 89.835 ;
        RECT -95.955 89.735 -95.585 90.075 ;
        RECT -95.405 89.835 -94.855 90.005 ;
        RECT -90.805 89.835 -90.255 90.005 ;
        RECT -95.405 89.510 -95.235 89.835 ;
        RECT -96.305 89.340 -95.235 89.510 ;
        RECT -90.425 89.510 -90.255 89.835 ;
        RECT -90.075 89.735 -89.705 90.075 ;
        RECT -89.525 89.835 -88.595 90.015 ;
        RECT -87.145 89.835 -86.215 90.015 ;
        RECT -89.525 89.510 -89.355 89.835 ;
        RECT -90.425 89.340 -89.355 89.510 ;
        RECT -86.385 89.510 -86.215 89.835 ;
        RECT -86.035 89.735 -85.665 90.075 ;
        RECT -85.485 89.835 -84.935 90.005 ;
        RECT -80.885 89.835 -80.335 90.005 ;
        RECT -85.485 89.510 -85.315 89.835 ;
        RECT -86.385 89.340 -85.315 89.510 ;
        RECT -80.505 89.510 -80.335 89.835 ;
        RECT -80.155 89.735 -79.785 90.075 ;
        RECT -79.605 89.835 -78.675 90.015 ;
        RECT -77.225 89.835 -76.295 90.015 ;
        RECT -79.605 89.510 -79.435 89.835 ;
        RECT -80.505 89.340 -79.435 89.510 ;
        RECT -76.465 89.510 -76.295 89.835 ;
        RECT -76.115 89.735 -75.745 90.075 ;
        RECT -75.565 89.835 -75.015 90.005 ;
        RECT -70.965 89.835 -70.415 90.005 ;
        RECT -75.565 89.510 -75.395 89.835 ;
        RECT -76.465 89.340 -75.395 89.510 ;
        RECT -70.585 89.510 -70.415 89.835 ;
        RECT -70.235 89.735 -69.865 90.075 ;
        RECT -69.685 89.835 -68.755 90.015 ;
        RECT -67.305 89.835 -66.375 90.015 ;
        RECT -69.685 89.510 -69.515 89.835 ;
        RECT -70.585 89.340 -69.515 89.510 ;
        RECT -66.545 89.510 -66.375 89.835 ;
        RECT -66.195 89.735 -65.825 90.075 ;
        RECT -65.645 89.835 -65.095 90.005 ;
        RECT -61.045 89.835 -60.495 90.005 ;
        RECT -65.645 89.510 -65.475 89.835 ;
        RECT -66.545 89.340 -65.475 89.510 ;
        RECT -60.665 89.510 -60.495 89.835 ;
        RECT -60.315 89.735 -59.945 90.075 ;
        RECT -59.765 89.835 -58.835 90.015 ;
        RECT -57.385 89.835 -56.455 90.015 ;
        RECT -59.765 89.510 -59.595 89.835 ;
        RECT -60.665 89.340 -59.595 89.510 ;
        RECT -56.625 89.510 -56.455 89.835 ;
        RECT -56.275 89.735 -55.905 90.075 ;
        RECT -55.725 89.835 -55.175 90.005 ;
        RECT -51.125 89.835 -50.575 90.005 ;
        RECT -55.725 89.510 -55.555 89.835 ;
        RECT -56.625 89.340 -55.555 89.510 ;
        RECT -50.745 89.510 -50.575 89.835 ;
        RECT -50.395 89.735 -50.025 90.075 ;
        RECT -49.845 89.835 -48.915 90.015 ;
        RECT -47.465 89.835 -46.535 90.015 ;
        RECT -49.845 89.510 -49.675 89.835 ;
        RECT -50.745 89.340 -49.675 89.510 ;
        RECT -46.705 89.510 -46.535 89.835 ;
        RECT -46.355 89.735 -45.985 90.075 ;
        RECT -45.805 89.835 -45.255 90.005 ;
        RECT -41.205 89.835 -40.655 90.005 ;
        RECT -45.805 89.510 -45.635 89.835 ;
        RECT -46.705 89.340 -45.635 89.510 ;
        RECT -40.825 89.510 -40.655 89.835 ;
        RECT -40.475 89.735 -40.105 90.075 ;
        RECT -39.925 89.835 -38.995 90.015 ;
        RECT -37.545 89.835 -36.615 90.015 ;
        RECT -39.925 89.510 -39.755 89.835 ;
        RECT -40.825 89.340 -39.755 89.510 ;
        RECT -36.785 89.510 -36.615 89.835 ;
        RECT -36.435 89.735 -36.065 90.075 ;
        RECT -35.885 89.835 -35.335 90.005 ;
        RECT -31.285 89.835 -30.735 90.005 ;
        RECT -35.885 89.510 -35.715 89.835 ;
        RECT -36.785 89.340 -35.715 89.510 ;
        RECT -30.905 89.510 -30.735 89.835 ;
        RECT -30.555 89.735 -30.185 90.075 ;
        RECT -30.005 89.835 -29.075 90.015 ;
        RECT -27.625 89.835 -26.695 90.015 ;
        RECT -30.005 89.510 -29.835 89.835 ;
        RECT -30.905 89.340 -29.835 89.510 ;
        RECT -26.865 89.510 -26.695 89.835 ;
        RECT -26.515 89.735 -26.145 90.075 ;
        RECT -25.965 89.835 -25.415 90.005 ;
        RECT -21.365 89.835 -20.815 90.005 ;
        RECT -25.965 89.510 -25.795 89.835 ;
        RECT -26.865 89.340 -25.795 89.510 ;
        RECT -20.985 89.510 -20.815 89.835 ;
        RECT -20.635 89.735 -20.265 90.075 ;
        RECT -20.085 89.835 -19.155 90.015 ;
        RECT -17.705 89.835 -16.775 90.015 ;
        RECT -20.085 89.510 -19.915 89.835 ;
        RECT -20.985 89.340 -19.915 89.510 ;
        RECT -16.945 89.510 -16.775 89.835 ;
        RECT -16.595 89.735 -16.225 90.075 ;
        RECT -16.045 89.835 -15.495 90.005 ;
        RECT -11.445 89.835 -10.895 90.005 ;
        RECT -16.045 89.510 -15.875 89.835 ;
        RECT -16.945 89.340 -15.875 89.510 ;
        RECT -11.065 89.510 -10.895 89.835 ;
        RECT -10.715 89.735 -10.345 90.075 ;
        RECT -10.165 89.835 -9.235 90.015 ;
        RECT -7.785 89.835 -6.855 90.015 ;
        RECT -10.165 89.510 -9.995 89.835 ;
        RECT -11.065 89.340 -9.995 89.510 ;
        RECT -7.025 89.510 -6.855 89.835 ;
        RECT -6.675 89.735 -6.305 90.075 ;
        RECT -6.125 89.835 -5.575 90.005 ;
        RECT -1.525 89.835 -0.975 90.005 ;
        RECT -6.125 89.510 -5.955 89.835 ;
        RECT -7.025 89.340 -5.955 89.510 ;
        RECT -1.145 89.510 -0.975 89.835 ;
        RECT -0.795 89.735 -0.425 90.075 ;
        RECT -0.245 89.835 0.685 90.015 ;
        RECT 2.135 89.835 3.065 90.015 ;
        RECT -0.245 89.510 -0.075 89.835 ;
        RECT -1.145 89.340 -0.075 89.510 ;
        RECT 2.895 89.510 3.065 89.835 ;
        RECT 3.245 89.735 3.615 90.075 ;
        RECT 3.795 89.835 4.345 90.005 ;
        RECT 8.395 89.835 8.945 90.005 ;
        RECT 3.795 89.510 3.965 89.835 ;
        RECT 2.895 89.340 3.965 89.510 ;
        RECT 8.775 89.510 8.945 89.835 ;
        RECT 9.125 89.735 9.495 90.075 ;
        RECT 9.675 89.835 10.605 90.015 ;
        RECT 12.055 89.835 12.985 90.015 ;
        RECT 9.675 89.510 9.845 89.835 ;
        RECT 8.775 89.340 9.845 89.510 ;
        RECT 12.815 89.510 12.985 89.835 ;
        RECT 13.165 89.735 13.535 90.075 ;
        RECT 13.715 89.835 14.265 90.005 ;
        RECT 18.315 89.835 18.865 90.005 ;
        RECT 13.715 89.510 13.885 89.835 ;
        RECT 12.815 89.340 13.885 89.510 ;
        RECT 18.695 89.510 18.865 89.835 ;
        RECT 19.045 89.735 19.415 90.075 ;
        RECT 19.595 89.835 20.525 90.015 ;
        RECT 21.975 89.835 22.905 90.015 ;
        RECT 19.595 89.510 19.765 89.835 ;
        RECT 18.695 89.340 19.765 89.510 ;
        RECT 22.735 89.510 22.905 89.835 ;
        RECT 23.085 89.735 23.455 90.075 ;
        RECT 23.635 89.835 24.185 90.005 ;
        RECT 23.635 89.510 23.805 89.835 ;
        RECT 24.355 89.655 24.525 90.180 ;
        RECT 22.735 89.340 23.805 89.510 ;
        RECT -289.545 89.140 -289.375 89.325 ;
        RECT -288.400 89.235 -288.070 89.340 ;
        RECT -284.470 89.235 -284.140 89.340 ;
        RECT -278.480 89.235 -278.150 89.340 ;
        RECT -274.550 89.235 -274.220 89.340 ;
        RECT -268.560 89.235 -268.230 89.340 ;
        RECT -264.630 89.235 -264.300 89.340 ;
        RECT -258.640 89.235 -258.310 89.340 ;
        RECT -254.710 89.235 -254.380 89.340 ;
        RECT -248.720 89.235 -248.390 89.340 ;
        RECT -244.790 89.235 -244.460 89.340 ;
        RECT -238.800 89.235 -238.470 89.340 ;
        RECT -234.870 89.235 -234.540 89.340 ;
        RECT -228.880 89.235 -228.550 89.340 ;
        RECT -224.950 89.235 -224.620 89.340 ;
        RECT -218.960 89.235 -218.630 89.340 ;
        RECT -215.030 89.235 -214.700 89.340 ;
        RECT -209.040 89.235 -208.710 89.340 ;
        RECT -205.110 89.235 -204.780 89.340 ;
        RECT -199.120 89.235 -198.790 89.340 ;
        RECT -195.190 89.235 -194.860 89.340 ;
        RECT -189.200 89.235 -188.870 89.340 ;
        RECT -185.270 89.235 -184.940 89.340 ;
        RECT -179.280 89.235 -178.950 89.340 ;
        RECT -175.350 89.235 -175.020 89.340 ;
        RECT -169.360 89.235 -169.030 89.340 ;
        RECT -165.430 89.235 -165.100 89.340 ;
        RECT -159.440 89.235 -159.110 89.340 ;
        RECT -155.510 89.235 -155.180 89.340 ;
        RECT -149.520 89.235 -149.190 89.340 ;
        RECT -145.590 89.235 -145.260 89.340 ;
        RECT -139.600 89.235 -139.270 89.340 ;
        RECT -135.670 89.235 -135.340 89.340 ;
        RECT -129.680 89.235 -129.350 89.340 ;
        RECT -125.750 89.235 -125.420 89.340 ;
        RECT -119.760 89.235 -119.430 89.340 ;
        RECT -115.830 89.235 -115.500 89.340 ;
        RECT -109.840 89.235 -109.510 89.340 ;
        RECT -105.910 89.235 -105.580 89.340 ;
        RECT -99.920 89.235 -99.590 89.340 ;
        RECT -95.990 89.235 -95.660 89.340 ;
        RECT -90.000 89.235 -89.670 89.340 ;
        RECT -86.070 89.235 -85.740 89.340 ;
        RECT -80.080 89.235 -79.750 89.340 ;
        RECT -76.150 89.235 -75.820 89.340 ;
        RECT -70.160 89.235 -69.830 89.340 ;
        RECT -66.230 89.235 -65.900 89.340 ;
        RECT -60.240 89.235 -59.910 89.340 ;
        RECT -56.310 89.235 -55.980 89.340 ;
        RECT -50.320 89.235 -49.990 89.340 ;
        RECT -46.390 89.235 -46.060 89.340 ;
        RECT -40.400 89.235 -40.070 89.340 ;
        RECT -36.470 89.235 -36.140 89.340 ;
        RECT -30.480 89.235 -30.150 89.340 ;
        RECT -26.550 89.235 -26.220 89.340 ;
        RECT -20.560 89.235 -20.230 89.340 ;
        RECT -16.630 89.235 -16.300 89.340 ;
        RECT -10.640 89.235 -10.310 89.340 ;
        RECT -6.710 89.235 -6.380 89.340 ;
        RECT -0.720 89.235 -0.390 89.340 ;
        RECT 3.210 89.235 3.540 89.340 ;
        RECT 9.200 89.235 9.530 89.340 ;
        RECT 13.130 89.235 13.460 89.340 ;
        RECT 19.120 89.235 19.450 89.340 ;
        RECT 23.050 89.235 23.380 89.340 ;
        RECT 23.975 89.325 24.525 89.655 ;
        RECT -290.075 89.125 -289.375 89.140 ;
        RECT -290.160 88.955 -289.375 89.125 ;
        RECT -289.840 88.950 -289.375 88.955 ;
        RECT -289.545 88.800 -289.375 88.950 ;
        RECT -285.545 89.065 -284.640 89.155 ;
        RECT -283.840 89.065 -283.335 89.145 ;
        RECT -285.545 88.885 -283.335 89.065 ;
        RECT -275.625 89.065 -274.720 89.155 ;
        RECT -273.920 89.065 -273.415 89.145 ;
        RECT -275.625 88.885 -273.415 89.065 ;
        RECT -265.705 89.065 -264.800 89.155 ;
        RECT -264.000 89.065 -263.495 89.145 ;
        RECT -265.705 88.885 -263.495 89.065 ;
        RECT -255.785 89.065 -254.880 89.155 ;
        RECT -254.080 89.065 -253.575 89.145 ;
        RECT -255.785 88.885 -253.575 89.065 ;
        RECT -245.865 89.065 -244.960 89.155 ;
        RECT -244.160 89.065 -243.655 89.145 ;
        RECT -245.865 88.885 -243.655 89.065 ;
        RECT -235.945 89.065 -235.040 89.155 ;
        RECT -234.240 89.065 -233.735 89.145 ;
        RECT -235.945 88.885 -233.735 89.065 ;
        RECT -226.025 89.065 -225.120 89.155 ;
        RECT -224.320 89.065 -223.815 89.145 ;
        RECT -226.025 88.885 -223.815 89.065 ;
        RECT -216.105 89.065 -215.200 89.155 ;
        RECT -214.400 89.065 -213.895 89.145 ;
        RECT -216.105 88.885 -213.895 89.065 ;
        RECT -206.185 89.065 -205.280 89.155 ;
        RECT -204.480 89.065 -203.975 89.145 ;
        RECT -206.185 88.885 -203.975 89.065 ;
        RECT -196.265 89.065 -195.360 89.155 ;
        RECT -194.560 89.065 -194.055 89.145 ;
        RECT -196.265 88.885 -194.055 89.065 ;
        RECT -186.345 89.065 -185.440 89.155 ;
        RECT -184.640 89.065 -184.135 89.145 ;
        RECT -186.345 88.885 -184.135 89.065 ;
        RECT -176.425 89.065 -175.520 89.155 ;
        RECT -174.720 89.065 -174.215 89.145 ;
        RECT -176.425 88.885 -174.215 89.065 ;
        RECT -166.505 89.065 -165.600 89.155 ;
        RECT -164.800 89.065 -164.295 89.145 ;
        RECT -166.505 88.885 -164.295 89.065 ;
        RECT -156.585 89.065 -155.680 89.155 ;
        RECT -154.880 89.065 -154.375 89.145 ;
        RECT -156.585 88.885 -154.375 89.065 ;
        RECT -146.665 89.065 -145.760 89.155 ;
        RECT -144.960 89.065 -144.455 89.145 ;
        RECT -146.665 88.885 -144.455 89.065 ;
        RECT -136.745 89.065 -135.840 89.155 ;
        RECT -135.040 89.065 -134.535 89.145 ;
        RECT -136.745 88.885 -134.535 89.065 ;
        RECT -126.825 89.065 -125.920 89.155 ;
        RECT -125.120 89.065 -124.615 89.145 ;
        RECT -126.825 88.885 -124.615 89.065 ;
        RECT -116.905 89.065 -116.000 89.155 ;
        RECT -115.200 89.065 -114.695 89.145 ;
        RECT -116.905 88.885 -114.695 89.065 ;
        RECT -106.985 89.065 -106.080 89.155 ;
        RECT -105.280 89.065 -104.775 89.145 ;
        RECT -106.985 88.885 -104.775 89.065 ;
        RECT -97.065 89.065 -96.160 89.155 ;
        RECT -95.360 89.065 -94.855 89.145 ;
        RECT -97.065 88.885 -94.855 89.065 ;
        RECT -87.145 89.065 -86.240 89.155 ;
        RECT -85.440 89.065 -84.935 89.145 ;
        RECT -87.145 88.885 -84.935 89.065 ;
        RECT -77.225 89.065 -76.320 89.155 ;
        RECT -75.520 89.065 -75.015 89.145 ;
        RECT -77.225 88.885 -75.015 89.065 ;
        RECT -67.305 89.065 -66.400 89.155 ;
        RECT -65.600 89.065 -65.095 89.145 ;
        RECT -67.305 88.885 -65.095 89.065 ;
        RECT -57.385 89.065 -56.480 89.155 ;
        RECT -55.680 89.065 -55.175 89.145 ;
        RECT -57.385 88.885 -55.175 89.065 ;
        RECT -47.465 89.065 -46.560 89.155 ;
        RECT -45.760 89.065 -45.255 89.145 ;
        RECT -47.465 88.885 -45.255 89.065 ;
        RECT -37.545 89.065 -36.640 89.155 ;
        RECT -35.840 89.065 -35.335 89.145 ;
        RECT -37.545 88.885 -35.335 89.065 ;
        RECT -27.625 89.065 -26.720 89.155 ;
        RECT -25.920 89.065 -25.415 89.145 ;
        RECT -27.625 88.885 -25.415 89.065 ;
        RECT -17.705 89.065 -16.800 89.155 ;
        RECT -16.000 89.065 -15.495 89.145 ;
        RECT -17.705 88.885 -15.495 89.065 ;
        RECT -7.785 89.065 -6.880 89.155 ;
        RECT -6.080 89.065 -5.575 89.145 ;
        RECT -7.785 88.885 -5.575 89.065 ;
        RECT 2.135 89.065 3.040 89.155 ;
        RECT 3.840 89.065 4.345 89.145 ;
        RECT 2.135 88.885 4.345 89.065 ;
        RECT 12.055 89.065 12.960 89.155 ;
        RECT 13.760 89.065 14.265 89.145 ;
        RECT 12.055 88.885 14.265 89.065 ;
        RECT 21.975 89.065 22.880 89.155 ;
        RECT 23.680 89.065 24.185 89.145 ;
        RECT 21.975 88.885 24.185 89.065 ;
        RECT 24.355 89.130 24.525 89.325 ;
        RECT 24.765 89.130 25.055 89.850 ;
        RECT 24.355 89.125 25.055 89.130 ;
        RECT 24.355 88.955 25.140 89.125 ;
        RECT 24.355 88.950 24.820 88.955 ;
        RECT 24.355 88.800 24.525 88.950 ;
        RECT -292.865 10.940 -292.695 11.090 ;
        RECT -293.480 10.770 -292.695 10.940 ;
        RECT -293.395 9.605 -293.105 10.770 ;
        RECT -292.865 10.565 -292.695 10.770 ;
        RECT -292.525 10.825 -290.315 11.005 ;
        RECT -292.525 10.735 -291.620 10.825 ;
        RECT -290.820 10.745 -290.315 10.825 ;
        RECT -282.605 10.825 -280.395 11.005 ;
        RECT -282.605 10.735 -281.700 10.825 ;
        RECT -280.900 10.745 -280.395 10.825 ;
        RECT -272.685 10.825 -270.475 11.005 ;
        RECT -272.685 10.735 -271.780 10.825 ;
        RECT -270.980 10.745 -270.475 10.825 ;
        RECT -262.765 10.825 -260.555 11.005 ;
        RECT -262.765 10.735 -261.860 10.825 ;
        RECT -261.060 10.745 -260.555 10.825 ;
        RECT -252.845 10.825 -250.635 11.005 ;
        RECT -252.845 10.735 -251.940 10.825 ;
        RECT -251.140 10.745 -250.635 10.825 ;
        RECT -242.925 10.825 -240.715 11.005 ;
        RECT -242.925 10.735 -242.020 10.825 ;
        RECT -241.220 10.745 -240.715 10.825 ;
        RECT -233.005 10.825 -230.795 11.005 ;
        RECT -233.005 10.735 -232.100 10.825 ;
        RECT -231.300 10.745 -230.795 10.825 ;
        RECT -223.085 10.825 -220.875 11.005 ;
        RECT -223.085 10.735 -222.180 10.825 ;
        RECT -221.380 10.745 -220.875 10.825 ;
        RECT -213.165 10.825 -210.955 11.005 ;
        RECT -213.165 10.735 -212.260 10.825 ;
        RECT -211.460 10.745 -210.955 10.825 ;
        RECT -203.245 10.825 -201.035 11.005 ;
        RECT -203.245 10.735 -202.340 10.825 ;
        RECT -201.540 10.745 -201.035 10.825 ;
        RECT -193.325 10.825 -191.115 11.005 ;
        RECT -193.325 10.735 -192.420 10.825 ;
        RECT -191.620 10.745 -191.115 10.825 ;
        RECT -183.405 10.825 -181.195 11.005 ;
        RECT -183.405 10.735 -182.500 10.825 ;
        RECT -181.700 10.745 -181.195 10.825 ;
        RECT -173.485 10.825 -171.275 11.005 ;
        RECT -173.485 10.735 -172.580 10.825 ;
        RECT -171.780 10.745 -171.275 10.825 ;
        RECT -163.565 10.825 -161.355 11.005 ;
        RECT -163.565 10.735 -162.660 10.825 ;
        RECT -161.860 10.745 -161.355 10.825 ;
        RECT -153.645 10.825 -151.435 11.005 ;
        RECT -153.645 10.735 -152.740 10.825 ;
        RECT -151.940 10.745 -151.435 10.825 ;
        RECT -143.725 10.825 -141.515 11.005 ;
        RECT -143.725 10.735 -142.820 10.825 ;
        RECT -142.020 10.745 -141.515 10.825 ;
        RECT -133.805 10.825 -131.595 11.005 ;
        RECT -133.805 10.735 -132.900 10.825 ;
        RECT -132.100 10.745 -131.595 10.825 ;
        RECT -123.885 10.825 -121.675 11.005 ;
        RECT -123.885 10.735 -122.980 10.825 ;
        RECT -122.180 10.745 -121.675 10.825 ;
        RECT -113.965 10.825 -111.755 11.005 ;
        RECT -113.965 10.735 -113.060 10.825 ;
        RECT -112.260 10.745 -111.755 10.825 ;
        RECT -104.045 10.825 -101.835 11.005 ;
        RECT -104.045 10.735 -103.140 10.825 ;
        RECT -102.340 10.745 -101.835 10.825 ;
        RECT -94.125 10.825 -91.915 11.005 ;
        RECT -94.125 10.735 -93.220 10.825 ;
        RECT -92.420 10.745 -91.915 10.825 ;
        RECT -84.205 10.825 -81.995 11.005 ;
        RECT -84.205 10.735 -83.300 10.825 ;
        RECT -82.500 10.745 -81.995 10.825 ;
        RECT -74.285 10.825 -72.075 11.005 ;
        RECT -74.285 10.735 -73.380 10.825 ;
        RECT -72.580 10.745 -72.075 10.825 ;
        RECT -64.365 10.825 -62.155 11.005 ;
        RECT -64.365 10.735 -63.460 10.825 ;
        RECT -62.660 10.745 -62.155 10.825 ;
        RECT -54.445 10.825 -52.235 11.005 ;
        RECT -54.445 10.735 -53.540 10.825 ;
        RECT -52.740 10.745 -52.235 10.825 ;
        RECT -44.525 10.825 -42.315 11.005 ;
        RECT -44.525 10.735 -43.620 10.825 ;
        RECT -42.820 10.745 -42.315 10.825 ;
        RECT -34.605 10.825 -32.395 11.005 ;
        RECT -34.605 10.735 -33.700 10.825 ;
        RECT -32.900 10.745 -32.395 10.825 ;
        RECT -24.685 10.825 -22.475 11.005 ;
        RECT -24.685 10.735 -23.780 10.825 ;
        RECT -22.980 10.745 -22.475 10.825 ;
        RECT -14.765 10.825 -12.555 11.005 ;
        RECT -14.765 10.735 -13.860 10.825 ;
        RECT -13.060 10.745 -12.555 10.825 ;
        RECT -4.845 10.825 -2.635 11.005 ;
        RECT -4.845 10.735 -3.940 10.825 ;
        RECT -3.140 10.745 -2.635 10.825 ;
        RECT 5.075 10.825 7.285 11.005 ;
        RECT 5.075 10.735 5.980 10.825 ;
        RECT 6.780 10.745 7.285 10.825 ;
        RECT 14.995 10.825 17.205 11.005 ;
        RECT 14.995 10.735 15.900 10.825 ;
        RECT 16.700 10.745 17.205 10.825 ;
        RECT -292.865 10.235 -291.935 10.565 ;
        RECT -291.450 10.550 -291.120 10.655 ;
        RECT -285.460 10.550 -285.130 10.655 ;
        RECT -281.530 10.550 -281.200 10.655 ;
        RECT -275.540 10.550 -275.210 10.655 ;
        RECT -271.610 10.550 -271.280 10.655 ;
        RECT -265.620 10.550 -265.290 10.655 ;
        RECT -261.690 10.550 -261.360 10.655 ;
        RECT -255.700 10.550 -255.370 10.655 ;
        RECT -251.770 10.550 -251.440 10.655 ;
        RECT -245.780 10.550 -245.450 10.655 ;
        RECT -241.850 10.550 -241.520 10.655 ;
        RECT -235.860 10.550 -235.530 10.655 ;
        RECT -231.930 10.550 -231.600 10.655 ;
        RECT -225.940 10.550 -225.610 10.655 ;
        RECT -222.010 10.550 -221.680 10.655 ;
        RECT -216.020 10.550 -215.690 10.655 ;
        RECT -212.090 10.550 -211.760 10.655 ;
        RECT -206.100 10.550 -205.770 10.655 ;
        RECT -202.170 10.550 -201.840 10.655 ;
        RECT -196.180 10.550 -195.850 10.655 ;
        RECT -192.250 10.550 -191.920 10.655 ;
        RECT -186.260 10.550 -185.930 10.655 ;
        RECT -182.330 10.550 -182.000 10.655 ;
        RECT -176.340 10.550 -176.010 10.655 ;
        RECT -172.410 10.550 -172.080 10.655 ;
        RECT -166.420 10.550 -166.090 10.655 ;
        RECT -162.490 10.550 -162.160 10.655 ;
        RECT -156.500 10.550 -156.170 10.655 ;
        RECT -152.570 10.550 -152.240 10.655 ;
        RECT -146.580 10.550 -146.250 10.655 ;
        RECT -142.650 10.550 -142.320 10.655 ;
        RECT -136.660 10.550 -136.330 10.655 ;
        RECT -132.730 10.550 -132.400 10.655 ;
        RECT -126.740 10.550 -126.410 10.655 ;
        RECT -122.810 10.550 -122.480 10.655 ;
        RECT -116.820 10.550 -116.490 10.655 ;
        RECT -112.890 10.550 -112.560 10.655 ;
        RECT -106.900 10.550 -106.570 10.655 ;
        RECT -102.970 10.550 -102.640 10.655 ;
        RECT -96.980 10.550 -96.650 10.655 ;
        RECT -93.050 10.550 -92.720 10.655 ;
        RECT -87.060 10.550 -86.730 10.655 ;
        RECT -83.130 10.550 -82.800 10.655 ;
        RECT -77.140 10.550 -76.810 10.655 ;
        RECT -73.210 10.550 -72.880 10.655 ;
        RECT -67.220 10.550 -66.890 10.655 ;
        RECT -63.290 10.550 -62.960 10.655 ;
        RECT -57.300 10.550 -56.970 10.655 ;
        RECT -53.370 10.550 -53.040 10.655 ;
        RECT -47.380 10.550 -47.050 10.655 ;
        RECT -43.450 10.550 -43.120 10.655 ;
        RECT -37.460 10.550 -37.130 10.655 ;
        RECT -33.530 10.550 -33.200 10.655 ;
        RECT -27.540 10.550 -27.210 10.655 ;
        RECT -23.610 10.550 -23.280 10.655 ;
        RECT -17.620 10.550 -17.290 10.655 ;
        RECT -13.690 10.550 -13.360 10.655 ;
        RECT -7.700 10.550 -7.370 10.655 ;
        RECT -3.770 10.550 -3.440 10.655 ;
        RECT 2.220 10.550 2.550 10.655 ;
        RECT 6.150 10.550 6.480 10.655 ;
        RECT 12.140 10.550 12.470 10.655 ;
        RECT 16.070 10.550 16.400 10.655 ;
        RECT 22.060 10.550 22.390 10.655 ;
        RECT -291.765 10.380 -290.695 10.550 ;
        RECT -292.865 9.710 -292.695 10.235 ;
        RECT -291.765 10.055 -291.595 10.380 ;
        RECT -292.525 9.875 -291.595 10.055 ;
        RECT -291.415 9.815 -291.045 10.155 ;
        RECT -290.865 10.055 -290.695 10.380 ;
        RECT -285.885 10.380 -284.815 10.550 ;
        RECT -285.885 10.055 -285.715 10.380 ;
        RECT -290.865 9.885 -290.315 10.055 ;
        RECT -286.265 9.885 -285.715 10.055 ;
        RECT -285.535 9.815 -285.165 10.155 ;
        RECT -284.985 10.055 -284.815 10.380 ;
        RECT -281.845 10.380 -280.775 10.550 ;
        RECT -281.845 10.055 -281.675 10.380 ;
        RECT -284.985 9.875 -284.055 10.055 ;
        RECT -282.605 9.875 -281.675 10.055 ;
        RECT -281.495 9.815 -281.125 10.155 ;
        RECT -280.945 10.055 -280.775 10.380 ;
        RECT -275.965 10.380 -274.895 10.550 ;
        RECT -275.965 10.055 -275.795 10.380 ;
        RECT -280.945 9.885 -280.395 10.055 ;
        RECT -276.345 9.885 -275.795 10.055 ;
        RECT -275.615 9.815 -275.245 10.155 ;
        RECT -275.065 10.055 -274.895 10.380 ;
        RECT -271.925 10.380 -270.855 10.550 ;
        RECT -271.925 10.055 -271.755 10.380 ;
        RECT -275.065 9.875 -274.135 10.055 ;
        RECT -272.685 9.875 -271.755 10.055 ;
        RECT -271.575 9.815 -271.205 10.155 ;
        RECT -271.025 10.055 -270.855 10.380 ;
        RECT -266.045 10.380 -264.975 10.550 ;
        RECT -266.045 10.055 -265.875 10.380 ;
        RECT -271.025 9.885 -270.475 10.055 ;
        RECT -266.425 9.885 -265.875 10.055 ;
        RECT -265.695 9.815 -265.325 10.155 ;
        RECT -265.145 10.055 -264.975 10.380 ;
        RECT -262.005 10.380 -260.935 10.550 ;
        RECT -262.005 10.055 -261.835 10.380 ;
        RECT -265.145 9.875 -264.215 10.055 ;
        RECT -262.765 9.875 -261.835 10.055 ;
        RECT -261.655 9.815 -261.285 10.155 ;
        RECT -261.105 10.055 -260.935 10.380 ;
        RECT -256.125 10.380 -255.055 10.550 ;
        RECT -256.125 10.055 -255.955 10.380 ;
        RECT -261.105 9.885 -260.555 10.055 ;
        RECT -256.505 9.885 -255.955 10.055 ;
        RECT -255.775 9.815 -255.405 10.155 ;
        RECT -255.225 10.055 -255.055 10.380 ;
        RECT -252.085 10.380 -251.015 10.550 ;
        RECT -252.085 10.055 -251.915 10.380 ;
        RECT -255.225 9.875 -254.295 10.055 ;
        RECT -252.845 9.875 -251.915 10.055 ;
        RECT -251.735 9.815 -251.365 10.155 ;
        RECT -251.185 10.055 -251.015 10.380 ;
        RECT -246.205 10.380 -245.135 10.550 ;
        RECT -246.205 10.055 -246.035 10.380 ;
        RECT -251.185 9.885 -250.635 10.055 ;
        RECT -246.585 9.885 -246.035 10.055 ;
        RECT -245.855 9.815 -245.485 10.155 ;
        RECT -245.305 10.055 -245.135 10.380 ;
        RECT -242.165 10.380 -241.095 10.550 ;
        RECT -242.165 10.055 -241.995 10.380 ;
        RECT -245.305 9.875 -244.375 10.055 ;
        RECT -242.925 9.875 -241.995 10.055 ;
        RECT -241.815 9.815 -241.445 10.155 ;
        RECT -241.265 10.055 -241.095 10.380 ;
        RECT -236.285 10.380 -235.215 10.550 ;
        RECT -236.285 10.055 -236.115 10.380 ;
        RECT -241.265 9.885 -240.715 10.055 ;
        RECT -236.665 9.885 -236.115 10.055 ;
        RECT -235.935 9.815 -235.565 10.155 ;
        RECT -235.385 10.055 -235.215 10.380 ;
        RECT -232.245 10.380 -231.175 10.550 ;
        RECT -232.245 10.055 -232.075 10.380 ;
        RECT -235.385 9.875 -234.455 10.055 ;
        RECT -233.005 9.875 -232.075 10.055 ;
        RECT -231.895 9.815 -231.525 10.155 ;
        RECT -231.345 10.055 -231.175 10.380 ;
        RECT -226.365 10.380 -225.295 10.550 ;
        RECT -226.365 10.055 -226.195 10.380 ;
        RECT -231.345 9.885 -230.795 10.055 ;
        RECT -226.745 9.885 -226.195 10.055 ;
        RECT -226.015 9.815 -225.645 10.155 ;
        RECT -225.465 10.055 -225.295 10.380 ;
        RECT -222.325 10.380 -221.255 10.550 ;
        RECT -222.325 10.055 -222.155 10.380 ;
        RECT -225.465 9.875 -224.535 10.055 ;
        RECT -223.085 9.875 -222.155 10.055 ;
        RECT -221.975 9.815 -221.605 10.155 ;
        RECT -221.425 10.055 -221.255 10.380 ;
        RECT -216.445 10.380 -215.375 10.550 ;
        RECT -216.445 10.055 -216.275 10.380 ;
        RECT -221.425 9.885 -220.875 10.055 ;
        RECT -216.825 9.885 -216.275 10.055 ;
        RECT -216.095 9.815 -215.725 10.155 ;
        RECT -215.545 10.055 -215.375 10.380 ;
        RECT -212.405 10.380 -211.335 10.550 ;
        RECT -212.405 10.055 -212.235 10.380 ;
        RECT -215.545 9.875 -214.615 10.055 ;
        RECT -213.165 9.875 -212.235 10.055 ;
        RECT -212.055 9.815 -211.685 10.155 ;
        RECT -211.505 10.055 -211.335 10.380 ;
        RECT -206.525 10.380 -205.455 10.550 ;
        RECT -206.525 10.055 -206.355 10.380 ;
        RECT -211.505 9.885 -210.955 10.055 ;
        RECT -206.905 9.885 -206.355 10.055 ;
        RECT -206.175 9.815 -205.805 10.155 ;
        RECT -205.625 10.055 -205.455 10.380 ;
        RECT -202.485 10.380 -201.415 10.550 ;
        RECT -202.485 10.055 -202.315 10.380 ;
        RECT -205.625 9.875 -204.695 10.055 ;
        RECT -203.245 9.875 -202.315 10.055 ;
        RECT -202.135 9.815 -201.765 10.155 ;
        RECT -201.585 10.055 -201.415 10.380 ;
        RECT -196.605 10.380 -195.535 10.550 ;
        RECT -196.605 10.055 -196.435 10.380 ;
        RECT -201.585 9.885 -201.035 10.055 ;
        RECT -196.985 9.885 -196.435 10.055 ;
        RECT -196.255 9.815 -195.885 10.155 ;
        RECT -195.705 10.055 -195.535 10.380 ;
        RECT -192.565 10.380 -191.495 10.550 ;
        RECT -192.565 10.055 -192.395 10.380 ;
        RECT -195.705 9.875 -194.775 10.055 ;
        RECT -193.325 9.875 -192.395 10.055 ;
        RECT -192.215 9.815 -191.845 10.155 ;
        RECT -191.665 10.055 -191.495 10.380 ;
        RECT -186.685 10.380 -185.615 10.550 ;
        RECT -186.685 10.055 -186.515 10.380 ;
        RECT -191.665 9.885 -191.115 10.055 ;
        RECT -187.065 9.885 -186.515 10.055 ;
        RECT -186.335 9.815 -185.965 10.155 ;
        RECT -185.785 10.055 -185.615 10.380 ;
        RECT -182.645 10.380 -181.575 10.550 ;
        RECT -182.645 10.055 -182.475 10.380 ;
        RECT -185.785 9.875 -184.855 10.055 ;
        RECT -183.405 9.875 -182.475 10.055 ;
        RECT -182.295 9.815 -181.925 10.155 ;
        RECT -181.745 10.055 -181.575 10.380 ;
        RECT -176.765 10.380 -175.695 10.550 ;
        RECT -176.765 10.055 -176.595 10.380 ;
        RECT -181.745 9.885 -181.195 10.055 ;
        RECT -177.145 9.885 -176.595 10.055 ;
        RECT -176.415 9.815 -176.045 10.155 ;
        RECT -175.865 10.055 -175.695 10.380 ;
        RECT -172.725 10.380 -171.655 10.550 ;
        RECT -172.725 10.055 -172.555 10.380 ;
        RECT -175.865 9.875 -174.935 10.055 ;
        RECT -173.485 9.875 -172.555 10.055 ;
        RECT -172.375 9.815 -172.005 10.155 ;
        RECT -171.825 10.055 -171.655 10.380 ;
        RECT -166.845 10.380 -165.775 10.550 ;
        RECT -166.845 10.055 -166.675 10.380 ;
        RECT -171.825 9.885 -171.275 10.055 ;
        RECT -167.225 9.885 -166.675 10.055 ;
        RECT -166.495 9.815 -166.125 10.155 ;
        RECT -165.945 10.055 -165.775 10.380 ;
        RECT -162.805 10.380 -161.735 10.550 ;
        RECT -162.805 10.055 -162.635 10.380 ;
        RECT -165.945 9.875 -165.015 10.055 ;
        RECT -163.565 9.875 -162.635 10.055 ;
        RECT -162.455 9.815 -162.085 10.155 ;
        RECT -161.905 10.055 -161.735 10.380 ;
        RECT -156.925 10.380 -155.855 10.550 ;
        RECT -156.925 10.055 -156.755 10.380 ;
        RECT -161.905 9.885 -161.355 10.055 ;
        RECT -157.305 9.885 -156.755 10.055 ;
        RECT -156.575 9.815 -156.205 10.155 ;
        RECT -156.025 10.055 -155.855 10.380 ;
        RECT -152.885 10.380 -151.815 10.550 ;
        RECT -152.885 10.055 -152.715 10.380 ;
        RECT -156.025 9.875 -155.095 10.055 ;
        RECT -153.645 9.875 -152.715 10.055 ;
        RECT -152.535 9.815 -152.165 10.155 ;
        RECT -151.985 10.055 -151.815 10.380 ;
        RECT -147.005 10.380 -145.935 10.550 ;
        RECT -147.005 10.055 -146.835 10.380 ;
        RECT -151.985 9.885 -151.435 10.055 ;
        RECT -147.385 9.885 -146.835 10.055 ;
        RECT -146.655 9.815 -146.285 10.155 ;
        RECT -146.105 10.055 -145.935 10.380 ;
        RECT -142.965 10.380 -141.895 10.550 ;
        RECT -142.965 10.055 -142.795 10.380 ;
        RECT -146.105 9.875 -145.175 10.055 ;
        RECT -143.725 9.875 -142.795 10.055 ;
        RECT -142.615 9.815 -142.245 10.155 ;
        RECT -142.065 10.055 -141.895 10.380 ;
        RECT -137.085 10.380 -136.015 10.550 ;
        RECT -137.085 10.055 -136.915 10.380 ;
        RECT -142.065 9.885 -141.515 10.055 ;
        RECT -137.465 9.885 -136.915 10.055 ;
        RECT -136.735 9.815 -136.365 10.155 ;
        RECT -136.185 10.055 -136.015 10.380 ;
        RECT -133.045 10.380 -131.975 10.550 ;
        RECT -133.045 10.055 -132.875 10.380 ;
        RECT -136.185 9.875 -135.255 10.055 ;
        RECT -133.805 9.875 -132.875 10.055 ;
        RECT -132.695 9.815 -132.325 10.155 ;
        RECT -132.145 10.055 -131.975 10.380 ;
        RECT -127.165 10.380 -126.095 10.550 ;
        RECT -127.165 10.055 -126.995 10.380 ;
        RECT -132.145 9.885 -131.595 10.055 ;
        RECT -127.545 9.885 -126.995 10.055 ;
        RECT -126.815 9.815 -126.445 10.155 ;
        RECT -126.265 10.055 -126.095 10.380 ;
        RECT -123.125 10.380 -122.055 10.550 ;
        RECT -123.125 10.055 -122.955 10.380 ;
        RECT -126.265 9.875 -125.335 10.055 ;
        RECT -123.885 9.875 -122.955 10.055 ;
        RECT -122.775 9.815 -122.405 10.155 ;
        RECT -122.225 10.055 -122.055 10.380 ;
        RECT -117.245 10.380 -116.175 10.550 ;
        RECT -117.245 10.055 -117.075 10.380 ;
        RECT -122.225 9.885 -121.675 10.055 ;
        RECT -117.625 9.885 -117.075 10.055 ;
        RECT -116.895 9.815 -116.525 10.155 ;
        RECT -116.345 10.055 -116.175 10.380 ;
        RECT -113.205 10.380 -112.135 10.550 ;
        RECT -113.205 10.055 -113.035 10.380 ;
        RECT -116.345 9.875 -115.415 10.055 ;
        RECT -113.965 9.875 -113.035 10.055 ;
        RECT -112.855 9.815 -112.485 10.155 ;
        RECT -112.305 10.055 -112.135 10.380 ;
        RECT -107.325 10.380 -106.255 10.550 ;
        RECT -107.325 10.055 -107.155 10.380 ;
        RECT -112.305 9.885 -111.755 10.055 ;
        RECT -107.705 9.885 -107.155 10.055 ;
        RECT -106.975 9.815 -106.605 10.155 ;
        RECT -106.425 10.055 -106.255 10.380 ;
        RECT -103.285 10.380 -102.215 10.550 ;
        RECT -103.285 10.055 -103.115 10.380 ;
        RECT -106.425 9.875 -105.495 10.055 ;
        RECT -104.045 9.875 -103.115 10.055 ;
        RECT -102.935 9.815 -102.565 10.155 ;
        RECT -102.385 10.055 -102.215 10.380 ;
        RECT -97.405 10.380 -96.335 10.550 ;
        RECT -97.405 10.055 -97.235 10.380 ;
        RECT -102.385 9.885 -101.835 10.055 ;
        RECT -97.785 9.885 -97.235 10.055 ;
        RECT -97.055 9.815 -96.685 10.155 ;
        RECT -96.505 10.055 -96.335 10.380 ;
        RECT -93.365 10.380 -92.295 10.550 ;
        RECT -93.365 10.055 -93.195 10.380 ;
        RECT -96.505 9.875 -95.575 10.055 ;
        RECT -94.125 9.875 -93.195 10.055 ;
        RECT -93.015 9.815 -92.645 10.155 ;
        RECT -92.465 10.055 -92.295 10.380 ;
        RECT -87.485 10.380 -86.415 10.550 ;
        RECT -87.485 10.055 -87.315 10.380 ;
        RECT -92.465 9.885 -91.915 10.055 ;
        RECT -87.865 9.885 -87.315 10.055 ;
        RECT -87.135 9.815 -86.765 10.155 ;
        RECT -86.585 10.055 -86.415 10.380 ;
        RECT -83.445 10.380 -82.375 10.550 ;
        RECT -83.445 10.055 -83.275 10.380 ;
        RECT -86.585 9.875 -85.655 10.055 ;
        RECT -84.205 9.875 -83.275 10.055 ;
        RECT -83.095 9.815 -82.725 10.155 ;
        RECT -82.545 10.055 -82.375 10.380 ;
        RECT -77.565 10.380 -76.495 10.550 ;
        RECT -77.565 10.055 -77.395 10.380 ;
        RECT -82.545 9.885 -81.995 10.055 ;
        RECT -77.945 9.885 -77.395 10.055 ;
        RECT -77.215 9.815 -76.845 10.155 ;
        RECT -76.665 10.055 -76.495 10.380 ;
        RECT -73.525 10.380 -72.455 10.550 ;
        RECT -73.525 10.055 -73.355 10.380 ;
        RECT -76.665 9.875 -75.735 10.055 ;
        RECT -74.285 9.875 -73.355 10.055 ;
        RECT -73.175 9.815 -72.805 10.155 ;
        RECT -72.625 10.055 -72.455 10.380 ;
        RECT -67.645 10.380 -66.575 10.550 ;
        RECT -67.645 10.055 -67.475 10.380 ;
        RECT -72.625 9.885 -72.075 10.055 ;
        RECT -68.025 9.885 -67.475 10.055 ;
        RECT -67.295 9.815 -66.925 10.155 ;
        RECT -66.745 10.055 -66.575 10.380 ;
        RECT -63.605 10.380 -62.535 10.550 ;
        RECT -63.605 10.055 -63.435 10.380 ;
        RECT -66.745 9.875 -65.815 10.055 ;
        RECT -64.365 9.875 -63.435 10.055 ;
        RECT -63.255 9.815 -62.885 10.155 ;
        RECT -62.705 10.055 -62.535 10.380 ;
        RECT -57.725 10.380 -56.655 10.550 ;
        RECT -57.725 10.055 -57.555 10.380 ;
        RECT -62.705 9.885 -62.155 10.055 ;
        RECT -58.105 9.885 -57.555 10.055 ;
        RECT -57.375 9.815 -57.005 10.155 ;
        RECT -56.825 10.055 -56.655 10.380 ;
        RECT -53.685 10.380 -52.615 10.550 ;
        RECT -53.685 10.055 -53.515 10.380 ;
        RECT -56.825 9.875 -55.895 10.055 ;
        RECT -54.445 9.875 -53.515 10.055 ;
        RECT -53.335 9.815 -52.965 10.155 ;
        RECT -52.785 10.055 -52.615 10.380 ;
        RECT -47.805 10.380 -46.735 10.550 ;
        RECT -47.805 10.055 -47.635 10.380 ;
        RECT -52.785 9.885 -52.235 10.055 ;
        RECT -48.185 9.885 -47.635 10.055 ;
        RECT -47.455 9.815 -47.085 10.155 ;
        RECT -46.905 10.055 -46.735 10.380 ;
        RECT -43.765 10.380 -42.695 10.550 ;
        RECT -43.765 10.055 -43.595 10.380 ;
        RECT -46.905 9.875 -45.975 10.055 ;
        RECT -44.525 9.875 -43.595 10.055 ;
        RECT -43.415 9.815 -43.045 10.155 ;
        RECT -42.865 10.055 -42.695 10.380 ;
        RECT -37.885 10.380 -36.815 10.550 ;
        RECT -37.885 10.055 -37.715 10.380 ;
        RECT -42.865 9.885 -42.315 10.055 ;
        RECT -38.265 9.885 -37.715 10.055 ;
        RECT -37.535 9.815 -37.165 10.155 ;
        RECT -36.985 10.055 -36.815 10.380 ;
        RECT -33.845 10.380 -32.775 10.550 ;
        RECT -33.845 10.055 -33.675 10.380 ;
        RECT -36.985 9.875 -36.055 10.055 ;
        RECT -34.605 9.875 -33.675 10.055 ;
        RECT -33.495 9.815 -33.125 10.155 ;
        RECT -32.945 10.055 -32.775 10.380 ;
        RECT -27.965 10.380 -26.895 10.550 ;
        RECT -27.965 10.055 -27.795 10.380 ;
        RECT -32.945 9.885 -32.395 10.055 ;
        RECT -28.345 9.885 -27.795 10.055 ;
        RECT -27.615 9.815 -27.245 10.155 ;
        RECT -27.065 10.055 -26.895 10.380 ;
        RECT -23.925 10.380 -22.855 10.550 ;
        RECT -23.925 10.055 -23.755 10.380 ;
        RECT -27.065 9.875 -26.135 10.055 ;
        RECT -24.685 9.875 -23.755 10.055 ;
        RECT -23.575 9.815 -23.205 10.155 ;
        RECT -23.025 10.055 -22.855 10.380 ;
        RECT -18.045 10.380 -16.975 10.550 ;
        RECT -18.045 10.055 -17.875 10.380 ;
        RECT -23.025 9.885 -22.475 10.055 ;
        RECT -18.425 9.885 -17.875 10.055 ;
        RECT -17.695 9.815 -17.325 10.155 ;
        RECT -17.145 10.055 -16.975 10.380 ;
        RECT -14.005 10.380 -12.935 10.550 ;
        RECT -14.005 10.055 -13.835 10.380 ;
        RECT -17.145 9.875 -16.215 10.055 ;
        RECT -14.765 9.875 -13.835 10.055 ;
        RECT -13.655 9.815 -13.285 10.155 ;
        RECT -13.105 10.055 -12.935 10.380 ;
        RECT -8.125 10.380 -7.055 10.550 ;
        RECT -8.125 10.055 -7.955 10.380 ;
        RECT -13.105 9.885 -12.555 10.055 ;
        RECT -8.505 9.885 -7.955 10.055 ;
        RECT -7.775 9.815 -7.405 10.155 ;
        RECT -7.225 10.055 -7.055 10.380 ;
        RECT -4.085 10.380 -3.015 10.550 ;
        RECT -4.085 10.055 -3.915 10.380 ;
        RECT -7.225 9.875 -6.295 10.055 ;
        RECT -4.845 9.875 -3.915 10.055 ;
        RECT -3.735 9.815 -3.365 10.155 ;
        RECT -3.185 10.055 -3.015 10.380 ;
        RECT 1.795 10.380 2.865 10.550 ;
        RECT 1.795 10.055 1.965 10.380 ;
        RECT -3.185 9.885 -2.635 10.055 ;
        RECT 1.415 9.885 1.965 10.055 ;
        RECT 2.145 9.815 2.515 10.155 ;
        RECT 2.695 10.055 2.865 10.380 ;
        RECT 5.835 10.380 6.905 10.550 ;
        RECT 5.835 10.055 6.005 10.380 ;
        RECT 2.695 9.875 3.625 10.055 ;
        RECT 5.075 9.875 6.005 10.055 ;
        RECT 6.185 9.815 6.555 10.155 ;
        RECT 6.735 10.055 6.905 10.380 ;
        RECT 11.715 10.380 12.785 10.550 ;
        RECT 11.715 10.055 11.885 10.380 ;
        RECT 6.735 9.885 7.285 10.055 ;
        RECT 11.335 9.885 11.885 10.055 ;
        RECT 12.065 9.815 12.435 10.155 ;
        RECT 12.615 10.055 12.785 10.380 ;
        RECT 15.755 10.380 16.825 10.550 ;
        RECT 15.755 10.055 15.925 10.380 ;
        RECT 12.615 9.875 13.545 10.055 ;
        RECT 14.995 9.875 15.925 10.055 ;
        RECT 16.105 9.815 16.475 10.155 ;
        RECT 16.655 10.055 16.825 10.380 ;
        RECT 21.635 10.380 22.705 10.550 ;
        RECT 21.635 10.055 21.805 10.380 ;
        RECT 16.655 9.885 17.205 10.055 ;
        RECT 21.255 9.885 21.805 10.055 ;
        RECT 21.985 9.815 22.355 10.155 ;
        RECT 22.535 10.055 22.705 10.380 ;
        RECT 22.535 9.875 23.465 10.055 ;
        RECT -293.480 9.195 -291.640 9.365 ;
        RECT 22.580 9.195 24.420 9.365 ;
        RECT -293.395 8.470 -293.105 9.195 ;
        RECT -292.935 8.395 -292.625 9.195 ;
        RECT -292.420 8.395 -291.725 9.025 ;
        RECT -293.395 6.645 -293.105 7.810 ;
        RECT -292.420 7.795 -292.250 8.395 ;
        RECT -292.080 7.955 -291.745 8.205 ;
        RECT -289.385 8.045 -289.055 9.025 ;
        RECT -287.525 8.045 -287.195 9.025 ;
        RECT -284.855 8.395 -284.160 9.025 ;
        RECT -292.935 6.645 -292.655 7.785 ;
        RECT -292.485 6.815 -292.155 7.795 ;
        RECT -291.985 6.645 -291.725 7.785 ;
        RECT -289.795 7.635 -289.460 7.885 ;
        RECT -289.290 7.445 -289.120 8.045 ;
        RECT -289.815 6.815 -289.120 7.445 ;
        RECT -287.460 7.445 -287.290 8.045 ;
        RECT -284.835 7.955 -284.500 8.205 ;
        RECT -287.120 7.635 -286.785 7.885 ;
        RECT -284.330 7.795 -284.160 8.395 ;
        RECT -282.500 8.395 -281.805 9.025 ;
        RECT -282.500 7.795 -282.330 8.395 ;
        RECT -282.160 7.955 -281.825 8.205 ;
        RECT -279.465 8.045 -279.135 9.025 ;
        RECT -277.605 8.045 -277.275 9.025 ;
        RECT -274.935 8.395 -274.240 9.025 ;
        RECT -287.460 6.815 -286.765 7.445 ;
        RECT -284.425 6.815 -284.095 7.795 ;
        RECT -282.565 6.815 -282.235 7.795 ;
        RECT -279.875 7.635 -279.540 7.885 ;
        RECT -279.370 7.445 -279.200 8.045 ;
        RECT -279.895 6.815 -279.200 7.445 ;
        RECT -277.540 7.445 -277.370 8.045 ;
        RECT -274.915 7.955 -274.580 8.205 ;
        RECT -277.200 7.635 -276.865 7.885 ;
        RECT -274.410 7.795 -274.240 8.395 ;
        RECT -272.580 8.395 -271.885 9.025 ;
        RECT -272.580 7.795 -272.410 8.395 ;
        RECT -272.240 7.955 -271.905 8.205 ;
        RECT -269.545 8.045 -269.215 9.025 ;
        RECT -267.685 8.045 -267.355 9.025 ;
        RECT -265.015 8.395 -264.320 9.025 ;
        RECT -277.540 6.815 -276.845 7.445 ;
        RECT -274.505 6.815 -274.175 7.795 ;
        RECT -272.645 6.815 -272.315 7.795 ;
        RECT -269.955 7.635 -269.620 7.885 ;
        RECT -269.450 7.445 -269.280 8.045 ;
        RECT -269.975 6.815 -269.280 7.445 ;
        RECT -267.620 7.445 -267.450 8.045 ;
        RECT -264.995 7.955 -264.660 8.205 ;
        RECT -267.280 7.635 -266.945 7.885 ;
        RECT -264.490 7.795 -264.320 8.395 ;
        RECT -262.660 8.395 -261.965 9.025 ;
        RECT -262.660 7.795 -262.490 8.395 ;
        RECT -262.320 7.955 -261.985 8.205 ;
        RECT -259.625 8.045 -259.295 9.025 ;
        RECT -257.765 8.045 -257.435 9.025 ;
        RECT -255.095 8.395 -254.400 9.025 ;
        RECT -267.620 6.815 -266.925 7.445 ;
        RECT -264.585 6.815 -264.255 7.795 ;
        RECT -262.725 6.815 -262.395 7.795 ;
        RECT -260.035 7.635 -259.700 7.885 ;
        RECT -259.530 7.445 -259.360 8.045 ;
        RECT -260.055 6.815 -259.360 7.445 ;
        RECT -257.700 7.445 -257.530 8.045 ;
        RECT -255.075 7.955 -254.740 8.205 ;
        RECT -257.360 7.635 -257.025 7.885 ;
        RECT -254.570 7.795 -254.400 8.395 ;
        RECT -252.740 8.395 -252.045 9.025 ;
        RECT -252.740 7.795 -252.570 8.395 ;
        RECT -252.400 7.955 -252.065 8.205 ;
        RECT -249.705 8.045 -249.375 9.025 ;
        RECT -247.845 8.045 -247.515 9.025 ;
        RECT -245.175 8.395 -244.480 9.025 ;
        RECT -257.700 6.815 -257.005 7.445 ;
        RECT -254.665 6.815 -254.335 7.795 ;
        RECT -252.805 6.815 -252.475 7.795 ;
        RECT -250.115 7.635 -249.780 7.885 ;
        RECT -249.610 7.445 -249.440 8.045 ;
        RECT -250.135 6.815 -249.440 7.445 ;
        RECT -247.780 7.445 -247.610 8.045 ;
        RECT -245.155 7.955 -244.820 8.205 ;
        RECT -247.440 7.635 -247.105 7.885 ;
        RECT -244.650 7.795 -244.480 8.395 ;
        RECT -242.820 8.395 -242.125 9.025 ;
        RECT -242.820 7.795 -242.650 8.395 ;
        RECT -242.480 7.955 -242.145 8.205 ;
        RECT -239.785 8.045 -239.455 9.025 ;
        RECT -237.925 8.045 -237.595 9.025 ;
        RECT -235.255 8.395 -234.560 9.025 ;
        RECT -247.780 6.815 -247.085 7.445 ;
        RECT -244.745 6.815 -244.415 7.795 ;
        RECT -242.885 6.815 -242.555 7.795 ;
        RECT -240.195 7.635 -239.860 7.885 ;
        RECT -239.690 7.445 -239.520 8.045 ;
        RECT -240.215 6.815 -239.520 7.445 ;
        RECT -237.860 7.445 -237.690 8.045 ;
        RECT -235.235 7.955 -234.900 8.205 ;
        RECT -237.520 7.635 -237.185 7.885 ;
        RECT -234.730 7.795 -234.560 8.395 ;
        RECT -232.900 8.395 -232.205 9.025 ;
        RECT -232.900 7.795 -232.730 8.395 ;
        RECT -232.560 7.955 -232.225 8.205 ;
        RECT -229.865 8.045 -229.535 9.025 ;
        RECT -228.005 8.045 -227.675 9.025 ;
        RECT -225.335 8.395 -224.640 9.025 ;
        RECT -237.860 6.815 -237.165 7.445 ;
        RECT -234.825 6.815 -234.495 7.795 ;
        RECT -232.965 6.815 -232.635 7.795 ;
        RECT -230.275 7.635 -229.940 7.885 ;
        RECT -229.770 7.445 -229.600 8.045 ;
        RECT -230.295 6.815 -229.600 7.445 ;
        RECT -227.940 7.445 -227.770 8.045 ;
        RECT -225.315 7.955 -224.980 8.205 ;
        RECT -227.600 7.635 -227.265 7.885 ;
        RECT -224.810 7.795 -224.640 8.395 ;
        RECT -222.980 8.395 -222.285 9.025 ;
        RECT -222.980 7.795 -222.810 8.395 ;
        RECT -222.640 7.955 -222.305 8.205 ;
        RECT -219.945 8.045 -219.615 9.025 ;
        RECT -218.085 8.045 -217.755 9.025 ;
        RECT -215.415 8.395 -214.720 9.025 ;
        RECT -227.940 6.815 -227.245 7.445 ;
        RECT -224.905 6.815 -224.575 7.795 ;
        RECT -223.045 6.815 -222.715 7.795 ;
        RECT -220.355 7.635 -220.020 7.885 ;
        RECT -219.850 7.445 -219.680 8.045 ;
        RECT -220.375 6.815 -219.680 7.445 ;
        RECT -218.020 7.445 -217.850 8.045 ;
        RECT -215.395 7.955 -215.060 8.205 ;
        RECT -217.680 7.635 -217.345 7.885 ;
        RECT -214.890 7.795 -214.720 8.395 ;
        RECT -213.060 8.395 -212.365 9.025 ;
        RECT -213.060 7.795 -212.890 8.395 ;
        RECT -212.720 7.955 -212.385 8.205 ;
        RECT -210.025 8.045 -209.695 9.025 ;
        RECT -208.165 8.045 -207.835 9.025 ;
        RECT -205.495 8.395 -204.800 9.025 ;
        RECT -218.020 6.815 -217.325 7.445 ;
        RECT -214.985 6.815 -214.655 7.795 ;
        RECT -213.125 6.815 -212.795 7.795 ;
        RECT -210.435 7.635 -210.100 7.885 ;
        RECT -209.930 7.445 -209.760 8.045 ;
        RECT -210.455 6.815 -209.760 7.445 ;
        RECT -208.100 7.445 -207.930 8.045 ;
        RECT -205.475 7.955 -205.140 8.205 ;
        RECT -207.760 7.635 -207.425 7.885 ;
        RECT -204.970 7.795 -204.800 8.395 ;
        RECT -203.140 8.395 -202.445 9.025 ;
        RECT -203.140 7.795 -202.970 8.395 ;
        RECT -202.800 7.955 -202.465 8.205 ;
        RECT -200.105 8.045 -199.775 9.025 ;
        RECT -198.245 8.045 -197.915 9.025 ;
        RECT -195.575 8.395 -194.880 9.025 ;
        RECT -208.100 6.815 -207.405 7.445 ;
        RECT -205.065 6.815 -204.735 7.795 ;
        RECT -203.205 6.815 -202.875 7.795 ;
        RECT -200.515 7.635 -200.180 7.885 ;
        RECT -200.010 7.445 -199.840 8.045 ;
        RECT -200.535 6.815 -199.840 7.445 ;
        RECT -198.180 7.445 -198.010 8.045 ;
        RECT -195.555 7.955 -195.220 8.205 ;
        RECT -197.840 7.635 -197.505 7.885 ;
        RECT -195.050 7.795 -194.880 8.395 ;
        RECT -193.220 8.395 -192.525 9.025 ;
        RECT -193.220 7.795 -193.050 8.395 ;
        RECT -192.880 7.955 -192.545 8.205 ;
        RECT -190.185 8.045 -189.855 9.025 ;
        RECT -188.325 8.045 -187.995 9.025 ;
        RECT -185.655 8.395 -184.960 9.025 ;
        RECT -198.180 6.815 -197.485 7.445 ;
        RECT -195.145 6.815 -194.815 7.795 ;
        RECT -193.285 6.815 -192.955 7.795 ;
        RECT -190.595 7.635 -190.260 7.885 ;
        RECT -190.090 7.445 -189.920 8.045 ;
        RECT -190.615 6.815 -189.920 7.445 ;
        RECT -188.260 7.445 -188.090 8.045 ;
        RECT -185.635 7.955 -185.300 8.205 ;
        RECT -187.920 7.635 -187.585 7.885 ;
        RECT -185.130 7.795 -184.960 8.395 ;
        RECT -183.300 8.395 -182.605 9.025 ;
        RECT -183.300 7.795 -183.130 8.395 ;
        RECT -182.960 7.955 -182.625 8.205 ;
        RECT -180.265 8.045 -179.935 9.025 ;
        RECT -178.405 8.045 -178.075 9.025 ;
        RECT -175.735 8.395 -175.040 9.025 ;
        RECT -188.260 6.815 -187.565 7.445 ;
        RECT -185.225 6.815 -184.895 7.795 ;
        RECT -183.365 6.815 -183.035 7.795 ;
        RECT -180.675 7.635 -180.340 7.885 ;
        RECT -180.170 7.445 -180.000 8.045 ;
        RECT -180.695 6.815 -180.000 7.445 ;
        RECT -178.340 7.445 -178.170 8.045 ;
        RECT -175.715 7.955 -175.380 8.205 ;
        RECT -178.000 7.635 -177.665 7.885 ;
        RECT -175.210 7.795 -175.040 8.395 ;
        RECT -173.380 8.395 -172.685 9.025 ;
        RECT -173.380 7.795 -173.210 8.395 ;
        RECT -173.040 7.955 -172.705 8.205 ;
        RECT -170.345 8.045 -170.015 9.025 ;
        RECT -168.485 8.045 -168.155 9.025 ;
        RECT -165.815 8.395 -165.120 9.025 ;
        RECT -178.340 6.815 -177.645 7.445 ;
        RECT -175.305 6.815 -174.975 7.795 ;
        RECT -173.445 6.815 -173.115 7.795 ;
        RECT -170.755 7.635 -170.420 7.885 ;
        RECT -170.250 7.445 -170.080 8.045 ;
        RECT -170.775 6.815 -170.080 7.445 ;
        RECT -168.420 7.445 -168.250 8.045 ;
        RECT -165.795 7.955 -165.460 8.205 ;
        RECT -168.080 7.635 -167.745 7.885 ;
        RECT -165.290 7.795 -165.120 8.395 ;
        RECT -163.460 8.395 -162.765 9.025 ;
        RECT -163.460 7.795 -163.290 8.395 ;
        RECT -163.120 7.955 -162.785 8.205 ;
        RECT -160.425 8.045 -160.095 9.025 ;
        RECT -158.565 8.045 -158.235 9.025 ;
        RECT -155.895 8.395 -155.200 9.025 ;
        RECT -168.420 6.815 -167.725 7.445 ;
        RECT -165.385 6.815 -165.055 7.795 ;
        RECT -163.525 6.815 -163.195 7.795 ;
        RECT -160.835 7.635 -160.500 7.885 ;
        RECT -160.330 7.445 -160.160 8.045 ;
        RECT -160.855 6.815 -160.160 7.445 ;
        RECT -158.500 7.445 -158.330 8.045 ;
        RECT -155.875 7.955 -155.540 8.205 ;
        RECT -158.160 7.635 -157.825 7.885 ;
        RECT -155.370 7.795 -155.200 8.395 ;
        RECT -153.540 8.395 -152.845 9.025 ;
        RECT -153.540 7.795 -153.370 8.395 ;
        RECT -153.200 7.955 -152.865 8.205 ;
        RECT -150.505 8.045 -150.175 9.025 ;
        RECT -148.645 8.045 -148.315 9.025 ;
        RECT -145.975 8.395 -145.280 9.025 ;
        RECT -158.500 6.815 -157.805 7.445 ;
        RECT -155.465 6.815 -155.135 7.795 ;
        RECT -153.605 6.815 -153.275 7.795 ;
        RECT -150.915 7.635 -150.580 7.885 ;
        RECT -150.410 7.445 -150.240 8.045 ;
        RECT -150.935 6.815 -150.240 7.445 ;
        RECT -148.580 7.445 -148.410 8.045 ;
        RECT -145.955 7.955 -145.620 8.205 ;
        RECT -148.240 7.635 -147.905 7.885 ;
        RECT -145.450 7.795 -145.280 8.395 ;
        RECT -143.620 8.395 -142.925 9.025 ;
        RECT -143.620 7.795 -143.450 8.395 ;
        RECT -143.280 7.955 -142.945 8.205 ;
        RECT -140.585 8.045 -140.255 9.025 ;
        RECT -138.725 8.045 -138.395 9.025 ;
        RECT -136.055 8.395 -135.360 9.025 ;
        RECT -148.580 6.815 -147.885 7.445 ;
        RECT -145.545 6.815 -145.215 7.795 ;
        RECT -143.685 6.815 -143.355 7.795 ;
        RECT -140.995 7.635 -140.660 7.885 ;
        RECT -140.490 7.445 -140.320 8.045 ;
        RECT -141.015 6.815 -140.320 7.445 ;
        RECT -138.660 7.445 -138.490 8.045 ;
        RECT -136.035 7.955 -135.700 8.205 ;
        RECT -138.320 7.635 -137.985 7.885 ;
        RECT -135.530 7.795 -135.360 8.395 ;
        RECT -133.700 8.395 -133.005 9.025 ;
        RECT -133.700 7.795 -133.530 8.395 ;
        RECT -133.360 7.955 -133.025 8.205 ;
        RECT -130.665 8.045 -130.335 9.025 ;
        RECT -128.805 8.045 -128.475 9.025 ;
        RECT -126.135 8.395 -125.440 9.025 ;
        RECT -138.660 6.815 -137.965 7.445 ;
        RECT -135.625 6.815 -135.295 7.795 ;
        RECT -133.765 6.815 -133.435 7.795 ;
        RECT -131.075 7.635 -130.740 7.885 ;
        RECT -130.570 7.445 -130.400 8.045 ;
        RECT -131.095 6.815 -130.400 7.445 ;
        RECT -128.740 7.445 -128.570 8.045 ;
        RECT -126.115 7.955 -125.780 8.205 ;
        RECT -128.400 7.635 -128.065 7.885 ;
        RECT -125.610 7.795 -125.440 8.395 ;
        RECT -123.780 8.395 -123.085 9.025 ;
        RECT -123.780 7.795 -123.610 8.395 ;
        RECT -123.440 7.955 -123.105 8.205 ;
        RECT -120.745 8.045 -120.415 9.025 ;
        RECT -118.885 8.045 -118.555 9.025 ;
        RECT -116.215 8.395 -115.520 9.025 ;
        RECT -128.740 6.815 -128.045 7.445 ;
        RECT -125.705 6.815 -125.375 7.795 ;
        RECT -123.845 6.815 -123.515 7.795 ;
        RECT -121.155 7.635 -120.820 7.885 ;
        RECT -120.650 7.445 -120.480 8.045 ;
        RECT -121.175 6.815 -120.480 7.445 ;
        RECT -118.820 7.445 -118.650 8.045 ;
        RECT -116.195 7.955 -115.860 8.205 ;
        RECT -118.480 7.635 -118.145 7.885 ;
        RECT -115.690 7.795 -115.520 8.395 ;
        RECT -113.860 8.395 -113.165 9.025 ;
        RECT -113.860 7.795 -113.690 8.395 ;
        RECT -113.520 7.955 -113.185 8.205 ;
        RECT -110.825 8.045 -110.495 9.025 ;
        RECT -108.965 8.045 -108.635 9.025 ;
        RECT -106.295 8.395 -105.600 9.025 ;
        RECT -118.820 6.815 -118.125 7.445 ;
        RECT -115.785 6.815 -115.455 7.795 ;
        RECT -113.925 6.815 -113.595 7.795 ;
        RECT -111.235 7.635 -110.900 7.885 ;
        RECT -110.730 7.445 -110.560 8.045 ;
        RECT -111.255 6.815 -110.560 7.445 ;
        RECT -108.900 7.445 -108.730 8.045 ;
        RECT -106.275 7.955 -105.940 8.205 ;
        RECT -108.560 7.635 -108.225 7.885 ;
        RECT -105.770 7.795 -105.600 8.395 ;
        RECT -103.940 8.395 -103.245 9.025 ;
        RECT -103.940 7.795 -103.770 8.395 ;
        RECT -103.600 7.955 -103.265 8.205 ;
        RECT -100.905 8.045 -100.575 9.025 ;
        RECT -99.045 8.045 -98.715 9.025 ;
        RECT -96.375 8.395 -95.680 9.025 ;
        RECT -108.900 6.815 -108.205 7.445 ;
        RECT -105.865 6.815 -105.535 7.795 ;
        RECT -104.005 6.815 -103.675 7.795 ;
        RECT -101.315 7.635 -100.980 7.885 ;
        RECT -100.810 7.445 -100.640 8.045 ;
        RECT -101.335 6.815 -100.640 7.445 ;
        RECT -98.980 7.445 -98.810 8.045 ;
        RECT -96.355 7.955 -96.020 8.205 ;
        RECT -98.640 7.635 -98.305 7.885 ;
        RECT -95.850 7.795 -95.680 8.395 ;
        RECT -94.020 8.395 -93.325 9.025 ;
        RECT -94.020 7.795 -93.850 8.395 ;
        RECT -93.680 7.955 -93.345 8.205 ;
        RECT -90.985 8.045 -90.655 9.025 ;
        RECT -89.125 8.045 -88.795 9.025 ;
        RECT -86.455 8.395 -85.760 9.025 ;
        RECT -98.980 6.815 -98.285 7.445 ;
        RECT -95.945 6.815 -95.615 7.795 ;
        RECT -94.085 6.815 -93.755 7.795 ;
        RECT -91.395 7.635 -91.060 7.885 ;
        RECT -90.890 7.445 -90.720 8.045 ;
        RECT -91.415 6.815 -90.720 7.445 ;
        RECT -89.060 7.445 -88.890 8.045 ;
        RECT -86.435 7.955 -86.100 8.205 ;
        RECT -88.720 7.635 -88.385 7.885 ;
        RECT -85.930 7.795 -85.760 8.395 ;
        RECT -84.100 8.395 -83.405 9.025 ;
        RECT -84.100 7.795 -83.930 8.395 ;
        RECT -83.760 7.955 -83.425 8.205 ;
        RECT -81.065 8.045 -80.735 9.025 ;
        RECT -79.205 8.045 -78.875 9.025 ;
        RECT -76.535 8.395 -75.840 9.025 ;
        RECT -89.060 6.815 -88.365 7.445 ;
        RECT -86.025 6.815 -85.695 7.795 ;
        RECT -84.165 6.815 -83.835 7.795 ;
        RECT -81.475 7.635 -81.140 7.885 ;
        RECT -80.970 7.445 -80.800 8.045 ;
        RECT -81.495 6.815 -80.800 7.445 ;
        RECT -79.140 7.445 -78.970 8.045 ;
        RECT -76.515 7.955 -76.180 8.205 ;
        RECT -78.800 7.635 -78.465 7.885 ;
        RECT -76.010 7.795 -75.840 8.395 ;
        RECT -74.180 8.395 -73.485 9.025 ;
        RECT -74.180 7.795 -74.010 8.395 ;
        RECT -73.840 7.955 -73.505 8.205 ;
        RECT -71.145 8.045 -70.815 9.025 ;
        RECT -69.285 8.045 -68.955 9.025 ;
        RECT -66.615 8.395 -65.920 9.025 ;
        RECT -79.140 6.815 -78.445 7.445 ;
        RECT -76.105 6.815 -75.775 7.795 ;
        RECT -74.245 6.815 -73.915 7.795 ;
        RECT -71.555 7.635 -71.220 7.885 ;
        RECT -71.050 7.445 -70.880 8.045 ;
        RECT -71.575 6.815 -70.880 7.445 ;
        RECT -69.220 7.445 -69.050 8.045 ;
        RECT -66.595 7.955 -66.260 8.205 ;
        RECT -68.880 7.635 -68.545 7.885 ;
        RECT -66.090 7.795 -65.920 8.395 ;
        RECT -64.260 8.395 -63.565 9.025 ;
        RECT -64.260 7.795 -64.090 8.395 ;
        RECT -63.920 7.955 -63.585 8.205 ;
        RECT -61.225 8.045 -60.895 9.025 ;
        RECT -59.365 8.045 -59.035 9.025 ;
        RECT -56.695 8.395 -56.000 9.025 ;
        RECT -69.220 6.815 -68.525 7.445 ;
        RECT -66.185 6.815 -65.855 7.795 ;
        RECT -64.325 6.815 -63.995 7.795 ;
        RECT -61.635 7.635 -61.300 7.885 ;
        RECT -61.130 7.445 -60.960 8.045 ;
        RECT -61.655 6.815 -60.960 7.445 ;
        RECT -59.300 7.445 -59.130 8.045 ;
        RECT -56.675 7.955 -56.340 8.205 ;
        RECT -58.960 7.635 -58.625 7.885 ;
        RECT -56.170 7.795 -56.000 8.395 ;
        RECT -54.340 8.395 -53.645 9.025 ;
        RECT -54.340 7.795 -54.170 8.395 ;
        RECT -54.000 7.955 -53.665 8.205 ;
        RECT -51.305 8.045 -50.975 9.025 ;
        RECT -49.445 8.045 -49.115 9.025 ;
        RECT -46.775 8.395 -46.080 9.025 ;
        RECT -59.300 6.815 -58.605 7.445 ;
        RECT -56.265 6.815 -55.935 7.795 ;
        RECT -54.405 6.815 -54.075 7.795 ;
        RECT -51.715 7.635 -51.380 7.885 ;
        RECT -51.210 7.445 -51.040 8.045 ;
        RECT -51.735 6.815 -51.040 7.445 ;
        RECT -49.380 7.445 -49.210 8.045 ;
        RECT -46.755 7.955 -46.420 8.205 ;
        RECT -49.040 7.635 -48.705 7.885 ;
        RECT -46.250 7.795 -46.080 8.395 ;
        RECT -44.420 8.395 -43.725 9.025 ;
        RECT -44.420 7.795 -44.250 8.395 ;
        RECT -44.080 7.955 -43.745 8.205 ;
        RECT -41.385 8.045 -41.055 9.025 ;
        RECT -39.525 8.045 -39.195 9.025 ;
        RECT -36.855 8.395 -36.160 9.025 ;
        RECT -49.380 6.815 -48.685 7.445 ;
        RECT -46.345 6.815 -46.015 7.795 ;
        RECT -44.485 6.815 -44.155 7.795 ;
        RECT -41.795 7.635 -41.460 7.885 ;
        RECT -41.290 7.445 -41.120 8.045 ;
        RECT -41.815 6.815 -41.120 7.445 ;
        RECT -39.460 7.445 -39.290 8.045 ;
        RECT -36.835 7.955 -36.500 8.205 ;
        RECT -39.120 7.635 -38.785 7.885 ;
        RECT -36.330 7.795 -36.160 8.395 ;
        RECT -34.500 8.395 -33.805 9.025 ;
        RECT -34.500 7.795 -34.330 8.395 ;
        RECT -34.160 7.955 -33.825 8.205 ;
        RECT -31.465 8.045 -31.135 9.025 ;
        RECT -29.605 8.045 -29.275 9.025 ;
        RECT -26.935 8.395 -26.240 9.025 ;
        RECT -39.460 6.815 -38.765 7.445 ;
        RECT -36.425 6.815 -36.095 7.795 ;
        RECT -34.565 6.815 -34.235 7.795 ;
        RECT -31.875 7.635 -31.540 7.885 ;
        RECT -31.370 7.445 -31.200 8.045 ;
        RECT -31.895 6.815 -31.200 7.445 ;
        RECT -29.540 7.445 -29.370 8.045 ;
        RECT -26.915 7.955 -26.580 8.205 ;
        RECT -29.200 7.635 -28.865 7.885 ;
        RECT -26.410 7.795 -26.240 8.395 ;
        RECT -24.580 8.395 -23.885 9.025 ;
        RECT -24.580 7.795 -24.410 8.395 ;
        RECT -24.240 7.955 -23.905 8.205 ;
        RECT -21.545 8.045 -21.215 9.025 ;
        RECT -19.685 8.045 -19.355 9.025 ;
        RECT -17.015 8.395 -16.320 9.025 ;
        RECT -29.540 6.815 -28.845 7.445 ;
        RECT -26.505 6.815 -26.175 7.795 ;
        RECT -24.645 6.815 -24.315 7.795 ;
        RECT -21.955 7.635 -21.620 7.885 ;
        RECT -21.450 7.445 -21.280 8.045 ;
        RECT -21.975 6.815 -21.280 7.445 ;
        RECT -19.620 7.445 -19.450 8.045 ;
        RECT -16.995 7.955 -16.660 8.205 ;
        RECT -19.280 7.635 -18.945 7.885 ;
        RECT -16.490 7.795 -16.320 8.395 ;
        RECT -14.660 8.395 -13.965 9.025 ;
        RECT -14.660 7.795 -14.490 8.395 ;
        RECT -14.320 7.955 -13.985 8.205 ;
        RECT -11.625 8.045 -11.295 9.025 ;
        RECT -9.765 8.045 -9.435 9.025 ;
        RECT -7.095 8.395 -6.400 9.025 ;
        RECT -19.620 6.815 -18.925 7.445 ;
        RECT -16.585 6.815 -16.255 7.795 ;
        RECT -14.725 6.815 -14.395 7.795 ;
        RECT -12.035 7.635 -11.700 7.885 ;
        RECT -11.530 7.445 -11.360 8.045 ;
        RECT -12.055 6.815 -11.360 7.445 ;
        RECT -9.700 7.445 -9.530 8.045 ;
        RECT -7.075 7.955 -6.740 8.205 ;
        RECT -9.360 7.635 -9.025 7.885 ;
        RECT -6.570 7.795 -6.400 8.395 ;
        RECT -4.740 8.395 -4.045 9.025 ;
        RECT -4.740 7.795 -4.570 8.395 ;
        RECT -4.400 7.955 -4.065 8.205 ;
        RECT -1.705 8.045 -1.375 9.025 ;
        RECT 0.155 8.045 0.485 9.025 ;
        RECT 2.825 8.395 3.520 9.025 ;
        RECT -9.700 6.815 -9.005 7.445 ;
        RECT -6.665 6.815 -6.335 7.795 ;
        RECT -4.805 6.815 -4.475 7.795 ;
        RECT -2.115 7.635 -1.780 7.885 ;
        RECT -1.610 7.445 -1.440 8.045 ;
        RECT -2.135 6.815 -1.440 7.445 ;
        RECT 0.220 7.445 0.390 8.045 ;
        RECT 2.845 7.955 3.180 8.205 ;
        RECT 0.560 7.635 0.895 7.885 ;
        RECT 3.350 7.795 3.520 8.395 ;
        RECT 5.180 8.395 5.875 9.025 ;
        RECT 5.180 7.795 5.350 8.395 ;
        RECT 5.520 7.955 5.855 8.205 ;
        RECT 8.215 8.045 8.545 9.025 ;
        RECT 10.075 8.045 10.405 9.025 ;
        RECT 12.745 8.395 13.440 9.025 ;
        RECT 0.220 6.815 0.915 7.445 ;
        RECT 3.255 6.815 3.585 7.795 ;
        RECT 5.115 6.815 5.445 7.795 ;
        RECT 7.805 7.635 8.140 7.885 ;
        RECT 8.310 7.445 8.480 8.045 ;
        RECT 7.785 6.815 8.480 7.445 ;
        RECT 10.140 7.445 10.310 8.045 ;
        RECT 12.765 7.955 13.100 8.205 ;
        RECT 10.480 7.635 10.815 7.885 ;
        RECT 13.270 7.795 13.440 8.395 ;
        RECT 15.100 8.395 15.795 9.025 ;
        RECT 15.100 7.795 15.270 8.395 ;
        RECT 15.440 7.955 15.775 8.205 ;
        RECT 18.135 8.045 18.465 9.025 ;
        RECT 19.995 8.045 20.325 9.025 ;
        RECT 22.665 8.395 23.360 9.025 ;
        RECT 23.565 8.395 23.875 9.195 ;
        RECT 24.045 8.470 24.335 9.195 ;
        RECT 10.140 6.815 10.835 7.445 ;
        RECT 13.175 6.815 13.505 7.795 ;
        RECT 15.035 6.815 15.365 7.795 ;
        RECT 17.725 7.635 18.060 7.885 ;
        RECT 18.230 7.445 18.400 8.045 ;
        RECT 17.705 6.815 18.400 7.445 ;
        RECT 20.060 7.445 20.230 8.045 ;
        RECT 22.685 7.955 23.020 8.205 ;
        RECT 20.400 7.635 20.735 7.885 ;
        RECT 23.190 7.795 23.360 8.395 ;
        RECT 20.060 6.815 20.755 7.445 ;
        RECT 23.095 6.815 23.425 7.795 ;
        RECT -293.480 6.475 -291.640 6.645 ;
        RECT -292.095 5.090 -291.805 5.800 ;
        RECT -291.565 5.605 -291.395 6.130 ;
        RECT -291.225 5.785 -290.675 5.955 ;
        RECT -291.565 5.275 -291.015 5.605 ;
        RECT -290.845 5.460 -290.675 5.785 ;
        RECT -290.495 5.685 -290.125 6.025 ;
        RECT -289.945 5.785 -289.015 5.965 ;
        RECT -287.565 5.785 -286.635 5.965 ;
        RECT -289.945 5.460 -289.775 5.785 ;
        RECT -290.845 5.290 -289.775 5.460 ;
        RECT -286.805 5.460 -286.635 5.785 ;
        RECT -286.455 5.685 -286.085 6.025 ;
        RECT -285.905 5.785 -285.355 5.955 ;
        RECT -281.305 5.785 -280.755 5.955 ;
        RECT -285.905 5.460 -285.735 5.785 ;
        RECT -286.805 5.290 -285.735 5.460 ;
        RECT -280.925 5.460 -280.755 5.785 ;
        RECT -280.575 5.685 -280.205 6.025 ;
        RECT -280.025 5.785 -279.095 5.965 ;
        RECT -277.645 5.785 -276.715 5.965 ;
        RECT -280.025 5.460 -279.855 5.785 ;
        RECT -280.925 5.290 -279.855 5.460 ;
        RECT -276.885 5.460 -276.715 5.785 ;
        RECT -276.535 5.685 -276.165 6.025 ;
        RECT -275.985 5.785 -275.435 5.955 ;
        RECT -271.385 5.785 -270.835 5.955 ;
        RECT -275.985 5.460 -275.815 5.785 ;
        RECT -276.885 5.290 -275.815 5.460 ;
        RECT -271.005 5.460 -270.835 5.785 ;
        RECT -270.655 5.685 -270.285 6.025 ;
        RECT -270.105 5.785 -269.175 5.965 ;
        RECT -267.725 5.785 -266.795 5.965 ;
        RECT -270.105 5.460 -269.935 5.785 ;
        RECT -271.005 5.290 -269.935 5.460 ;
        RECT -266.965 5.460 -266.795 5.785 ;
        RECT -266.615 5.685 -266.245 6.025 ;
        RECT -266.065 5.785 -265.515 5.955 ;
        RECT -261.465 5.785 -260.915 5.955 ;
        RECT -266.065 5.460 -265.895 5.785 ;
        RECT -266.965 5.290 -265.895 5.460 ;
        RECT -261.085 5.460 -260.915 5.785 ;
        RECT -260.735 5.685 -260.365 6.025 ;
        RECT -260.185 5.785 -259.255 5.965 ;
        RECT -257.805 5.785 -256.875 5.965 ;
        RECT -260.185 5.460 -260.015 5.785 ;
        RECT -261.085 5.290 -260.015 5.460 ;
        RECT -257.045 5.460 -256.875 5.785 ;
        RECT -256.695 5.685 -256.325 6.025 ;
        RECT -256.145 5.785 -255.595 5.955 ;
        RECT -251.545 5.785 -250.995 5.955 ;
        RECT -256.145 5.460 -255.975 5.785 ;
        RECT -257.045 5.290 -255.975 5.460 ;
        RECT -251.165 5.460 -250.995 5.785 ;
        RECT -250.815 5.685 -250.445 6.025 ;
        RECT -250.265 5.785 -249.335 5.965 ;
        RECT -247.885 5.785 -246.955 5.965 ;
        RECT -250.265 5.460 -250.095 5.785 ;
        RECT -251.165 5.290 -250.095 5.460 ;
        RECT -247.125 5.460 -246.955 5.785 ;
        RECT -246.775 5.685 -246.405 6.025 ;
        RECT -246.225 5.785 -245.675 5.955 ;
        RECT -241.625 5.785 -241.075 5.955 ;
        RECT -246.225 5.460 -246.055 5.785 ;
        RECT -247.125 5.290 -246.055 5.460 ;
        RECT -241.245 5.460 -241.075 5.785 ;
        RECT -240.895 5.685 -240.525 6.025 ;
        RECT -240.345 5.785 -239.415 5.965 ;
        RECT -237.965 5.785 -237.035 5.965 ;
        RECT -240.345 5.460 -240.175 5.785 ;
        RECT -241.245 5.290 -240.175 5.460 ;
        RECT -237.205 5.460 -237.035 5.785 ;
        RECT -236.855 5.685 -236.485 6.025 ;
        RECT -236.305 5.785 -235.755 5.955 ;
        RECT -231.705 5.785 -231.155 5.955 ;
        RECT -236.305 5.460 -236.135 5.785 ;
        RECT -237.205 5.290 -236.135 5.460 ;
        RECT -231.325 5.460 -231.155 5.785 ;
        RECT -230.975 5.685 -230.605 6.025 ;
        RECT -230.425 5.785 -229.495 5.965 ;
        RECT -228.045 5.785 -227.115 5.965 ;
        RECT -230.425 5.460 -230.255 5.785 ;
        RECT -231.325 5.290 -230.255 5.460 ;
        RECT -227.285 5.460 -227.115 5.785 ;
        RECT -226.935 5.685 -226.565 6.025 ;
        RECT -226.385 5.785 -225.835 5.955 ;
        RECT -221.785 5.785 -221.235 5.955 ;
        RECT -226.385 5.460 -226.215 5.785 ;
        RECT -227.285 5.290 -226.215 5.460 ;
        RECT -221.405 5.460 -221.235 5.785 ;
        RECT -221.055 5.685 -220.685 6.025 ;
        RECT -220.505 5.785 -219.575 5.965 ;
        RECT -218.125 5.785 -217.195 5.965 ;
        RECT -220.505 5.460 -220.335 5.785 ;
        RECT -221.405 5.290 -220.335 5.460 ;
        RECT -217.365 5.460 -217.195 5.785 ;
        RECT -217.015 5.685 -216.645 6.025 ;
        RECT -216.465 5.785 -215.915 5.955 ;
        RECT -211.865 5.785 -211.315 5.955 ;
        RECT -216.465 5.460 -216.295 5.785 ;
        RECT -217.365 5.290 -216.295 5.460 ;
        RECT -211.485 5.460 -211.315 5.785 ;
        RECT -211.135 5.685 -210.765 6.025 ;
        RECT -210.585 5.785 -209.655 5.965 ;
        RECT -208.205 5.785 -207.275 5.965 ;
        RECT -210.585 5.460 -210.415 5.785 ;
        RECT -211.485 5.290 -210.415 5.460 ;
        RECT -207.445 5.460 -207.275 5.785 ;
        RECT -207.095 5.685 -206.725 6.025 ;
        RECT -206.545 5.785 -205.995 5.955 ;
        RECT -201.945 5.785 -201.395 5.955 ;
        RECT -206.545 5.460 -206.375 5.785 ;
        RECT -207.445 5.290 -206.375 5.460 ;
        RECT -201.565 5.460 -201.395 5.785 ;
        RECT -201.215 5.685 -200.845 6.025 ;
        RECT -200.665 5.785 -199.735 5.965 ;
        RECT -198.285 5.785 -197.355 5.965 ;
        RECT -200.665 5.460 -200.495 5.785 ;
        RECT -201.565 5.290 -200.495 5.460 ;
        RECT -197.525 5.460 -197.355 5.785 ;
        RECT -197.175 5.685 -196.805 6.025 ;
        RECT -196.625 5.785 -196.075 5.955 ;
        RECT -192.025 5.785 -191.475 5.955 ;
        RECT -196.625 5.460 -196.455 5.785 ;
        RECT -197.525 5.290 -196.455 5.460 ;
        RECT -191.645 5.460 -191.475 5.785 ;
        RECT -191.295 5.685 -190.925 6.025 ;
        RECT -190.745 5.785 -189.815 5.965 ;
        RECT -188.365 5.785 -187.435 5.965 ;
        RECT -190.745 5.460 -190.575 5.785 ;
        RECT -191.645 5.290 -190.575 5.460 ;
        RECT -187.605 5.460 -187.435 5.785 ;
        RECT -187.255 5.685 -186.885 6.025 ;
        RECT -186.705 5.785 -186.155 5.955 ;
        RECT -182.105 5.785 -181.555 5.955 ;
        RECT -186.705 5.460 -186.535 5.785 ;
        RECT -187.605 5.290 -186.535 5.460 ;
        RECT -181.725 5.460 -181.555 5.785 ;
        RECT -181.375 5.685 -181.005 6.025 ;
        RECT -180.825 5.785 -179.895 5.965 ;
        RECT -178.445 5.785 -177.515 5.965 ;
        RECT -180.825 5.460 -180.655 5.785 ;
        RECT -181.725 5.290 -180.655 5.460 ;
        RECT -177.685 5.460 -177.515 5.785 ;
        RECT -177.335 5.685 -176.965 6.025 ;
        RECT -176.785 5.785 -176.235 5.955 ;
        RECT -172.185 5.785 -171.635 5.955 ;
        RECT -176.785 5.460 -176.615 5.785 ;
        RECT -177.685 5.290 -176.615 5.460 ;
        RECT -171.805 5.460 -171.635 5.785 ;
        RECT -171.455 5.685 -171.085 6.025 ;
        RECT -170.905 5.785 -169.975 5.965 ;
        RECT -168.525 5.785 -167.595 5.965 ;
        RECT -170.905 5.460 -170.735 5.785 ;
        RECT -171.805 5.290 -170.735 5.460 ;
        RECT -167.765 5.460 -167.595 5.785 ;
        RECT -167.415 5.685 -167.045 6.025 ;
        RECT -166.865 5.785 -166.315 5.955 ;
        RECT -162.265 5.785 -161.715 5.955 ;
        RECT -166.865 5.460 -166.695 5.785 ;
        RECT -167.765 5.290 -166.695 5.460 ;
        RECT -161.885 5.460 -161.715 5.785 ;
        RECT -161.535 5.685 -161.165 6.025 ;
        RECT -160.985 5.785 -160.055 5.965 ;
        RECT -158.605 5.785 -157.675 5.965 ;
        RECT -160.985 5.460 -160.815 5.785 ;
        RECT -161.885 5.290 -160.815 5.460 ;
        RECT -157.845 5.460 -157.675 5.785 ;
        RECT -157.495 5.685 -157.125 6.025 ;
        RECT -156.945 5.785 -156.395 5.955 ;
        RECT -152.345 5.785 -151.795 5.955 ;
        RECT -156.945 5.460 -156.775 5.785 ;
        RECT -157.845 5.290 -156.775 5.460 ;
        RECT -151.965 5.460 -151.795 5.785 ;
        RECT -151.615 5.685 -151.245 6.025 ;
        RECT -151.065 5.785 -150.135 5.965 ;
        RECT -148.685 5.785 -147.755 5.965 ;
        RECT -151.065 5.460 -150.895 5.785 ;
        RECT -151.965 5.290 -150.895 5.460 ;
        RECT -147.925 5.460 -147.755 5.785 ;
        RECT -147.575 5.685 -147.205 6.025 ;
        RECT -147.025 5.785 -146.475 5.955 ;
        RECT -142.425 5.785 -141.875 5.955 ;
        RECT -147.025 5.460 -146.855 5.785 ;
        RECT -147.925 5.290 -146.855 5.460 ;
        RECT -142.045 5.460 -141.875 5.785 ;
        RECT -141.695 5.685 -141.325 6.025 ;
        RECT -141.145 5.785 -140.215 5.965 ;
        RECT -138.765 5.785 -137.835 5.965 ;
        RECT -141.145 5.460 -140.975 5.785 ;
        RECT -142.045 5.290 -140.975 5.460 ;
        RECT -138.005 5.460 -137.835 5.785 ;
        RECT -137.655 5.685 -137.285 6.025 ;
        RECT -137.105 5.785 -136.555 5.955 ;
        RECT -132.505 5.785 -131.955 5.955 ;
        RECT -137.105 5.460 -136.935 5.785 ;
        RECT -138.005 5.290 -136.935 5.460 ;
        RECT -132.125 5.460 -131.955 5.785 ;
        RECT -131.775 5.685 -131.405 6.025 ;
        RECT -131.225 5.785 -130.295 5.965 ;
        RECT -128.845 5.785 -127.915 5.965 ;
        RECT -131.225 5.460 -131.055 5.785 ;
        RECT -132.125 5.290 -131.055 5.460 ;
        RECT -128.085 5.460 -127.915 5.785 ;
        RECT -127.735 5.685 -127.365 6.025 ;
        RECT -127.185 5.785 -126.635 5.955 ;
        RECT -122.585 5.785 -122.035 5.955 ;
        RECT -127.185 5.460 -127.015 5.785 ;
        RECT -128.085 5.290 -127.015 5.460 ;
        RECT -122.205 5.460 -122.035 5.785 ;
        RECT -121.855 5.685 -121.485 6.025 ;
        RECT -121.305 5.785 -120.375 5.965 ;
        RECT -118.925 5.785 -117.995 5.965 ;
        RECT -121.305 5.460 -121.135 5.785 ;
        RECT -122.205 5.290 -121.135 5.460 ;
        RECT -118.165 5.460 -117.995 5.785 ;
        RECT -117.815 5.685 -117.445 6.025 ;
        RECT -117.265 5.785 -116.715 5.955 ;
        RECT -112.665 5.785 -112.115 5.955 ;
        RECT -117.265 5.460 -117.095 5.785 ;
        RECT -118.165 5.290 -117.095 5.460 ;
        RECT -112.285 5.460 -112.115 5.785 ;
        RECT -111.935 5.685 -111.565 6.025 ;
        RECT -111.385 5.785 -110.455 5.965 ;
        RECT -109.005 5.785 -108.075 5.965 ;
        RECT -111.385 5.460 -111.215 5.785 ;
        RECT -112.285 5.290 -111.215 5.460 ;
        RECT -108.245 5.460 -108.075 5.785 ;
        RECT -107.895 5.685 -107.525 6.025 ;
        RECT -107.345 5.785 -106.795 5.955 ;
        RECT -102.745 5.785 -102.195 5.955 ;
        RECT -107.345 5.460 -107.175 5.785 ;
        RECT -108.245 5.290 -107.175 5.460 ;
        RECT -102.365 5.460 -102.195 5.785 ;
        RECT -102.015 5.685 -101.645 6.025 ;
        RECT -101.465 5.785 -100.535 5.965 ;
        RECT -99.085 5.785 -98.155 5.965 ;
        RECT -101.465 5.460 -101.295 5.785 ;
        RECT -102.365 5.290 -101.295 5.460 ;
        RECT -98.325 5.460 -98.155 5.785 ;
        RECT -97.975 5.685 -97.605 6.025 ;
        RECT -97.425 5.785 -96.875 5.955 ;
        RECT -92.825 5.785 -92.275 5.955 ;
        RECT -97.425 5.460 -97.255 5.785 ;
        RECT -98.325 5.290 -97.255 5.460 ;
        RECT -92.445 5.460 -92.275 5.785 ;
        RECT -92.095 5.685 -91.725 6.025 ;
        RECT -91.545 5.785 -90.615 5.965 ;
        RECT -89.165 5.785 -88.235 5.965 ;
        RECT -91.545 5.460 -91.375 5.785 ;
        RECT -92.445 5.290 -91.375 5.460 ;
        RECT -88.405 5.460 -88.235 5.785 ;
        RECT -88.055 5.685 -87.685 6.025 ;
        RECT -87.505 5.785 -86.955 5.955 ;
        RECT -82.905 5.785 -82.355 5.955 ;
        RECT -87.505 5.460 -87.335 5.785 ;
        RECT -88.405 5.290 -87.335 5.460 ;
        RECT -82.525 5.460 -82.355 5.785 ;
        RECT -82.175 5.685 -81.805 6.025 ;
        RECT -81.625 5.785 -80.695 5.965 ;
        RECT -79.245 5.785 -78.315 5.965 ;
        RECT -81.625 5.460 -81.455 5.785 ;
        RECT -82.525 5.290 -81.455 5.460 ;
        RECT -78.485 5.460 -78.315 5.785 ;
        RECT -78.135 5.685 -77.765 6.025 ;
        RECT -77.585 5.785 -77.035 5.955 ;
        RECT -72.985 5.785 -72.435 5.955 ;
        RECT -77.585 5.460 -77.415 5.785 ;
        RECT -78.485 5.290 -77.415 5.460 ;
        RECT -72.605 5.460 -72.435 5.785 ;
        RECT -72.255 5.685 -71.885 6.025 ;
        RECT -71.705 5.785 -70.775 5.965 ;
        RECT -69.325 5.785 -68.395 5.965 ;
        RECT -71.705 5.460 -71.535 5.785 ;
        RECT -72.605 5.290 -71.535 5.460 ;
        RECT -68.565 5.460 -68.395 5.785 ;
        RECT -68.215 5.685 -67.845 6.025 ;
        RECT -67.665 5.785 -67.115 5.955 ;
        RECT -63.065 5.785 -62.515 5.955 ;
        RECT -67.665 5.460 -67.495 5.785 ;
        RECT -68.565 5.290 -67.495 5.460 ;
        RECT -62.685 5.460 -62.515 5.785 ;
        RECT -62.335 5.685 -61.965 6.025 ;
        RECT -61.785 5.785 -60.855 5.965 ;
        RECT -59.405 5.785 -58.475 5.965 ;
        RECT -61.785 5.460 -61.615 5.785 ;
        RECT -62.685 5.290 -61.615 5.460 ;
        RECT -58.645 5.460 -58.475 5.785 ;
        RECT -58.295 5.685 -57.925 6.025 ;
        RECT -57.745 5.785 -57.195 5.955 ;
        RECT -53.145 5.785 -52.595 5.955 ;
        RECT -57.745 5.460 -57.575 5.785 ;
        RECT -58.645 5.290 -57.575 5.460 ;
        RECT -52.765 5.460 -52.595 5.785 ;
        RECT -52.415 5.685 -52.045 6.025 ;
        RECT -51.865 5.785 -50.935 5.965 ;
        RECT -49.485 5.785 -48.555 5.965 ;
        RECT -51.865 5.460 -51.695 5.785 ;
        RECT -52.765 5.290 -51.695 5.460 ;
        RECT -48.725 5.460 -48.555 5.785 ;
        RECT -48.375 5.685 -48.005 6.025 ;
        RECT -47.825 5.785 -47.275 5.955 ;
        RECT -43.225 5.785 -42.675 5.955 ;
        RECT -47.825 5.460 -47.655 5.785 ;
        RECT -48.725 5.290 -47.655 5.460 ;
        RECT -42.845 5.460 -42.675 5.785 ;
        RECT -42.495 5.685 -42.125 6.025 ;
        RECT -41.945 5.785 -41.015 5.965 ;
        RECT -39.565 5.785 -38.635 5.965 ;
        RECT -41.945 5.460 -41.775 5.785 ;
        RECT -42.845 5.290 -41.775 5.460 ;
        RECT -38.805 5.460 -38.635 5.785 ;
        RECT -38.455 5.685 -38.085 6.025 ;
        RECT -37.905 5.785 -37.355 5.955 ;
        RECT -33.305 5.785 -32.755 5.955 ;
        RECT -37.905 5.460 -37.735 5.785 ;
        RECT -38.805 5.290 -37.735 5.460 ;
        RECT -32.925 5.460 -32.755 5.785 ;
        RECT -32.575 5.685 -32.205 6.025 ;
        RECT -32.025 5.785 -31.095 5.965 ;
        RECT -29.645 5.785 -28.715 5.965 ;
        RECT -32.025 5.460 -31.855 5.785 ;
        RECT -32.925 5.290 -31.855 5.460 ;
        RECT -28.885 5.460 -28.715 5.785 ;
        RECT -28.535 5.685 -28.165 6.025 ;
        RECT -27.985 5.785 -27.435 5.955 ;
        RECT -23.385 5.785 -22.835 5.955 ;
        RECT -27.985 5.460 -27.815 5.785 ;
        RECT -28.885 5.290 -27.815 5.460 ;
        RECT -23.005 5.460 -22.835 5.785 ;
        RECT -22.655 5.685 -22.285 6.025 ;
        RECT -22.105 5.785 -21.175 5.965 ;
        RECT -19.725 5.785 -18.795 5.965 ;
        RECT -22.105 5.460 -21.935 5.785 ;
        RECT -23.005 5.290 -21.935 5.460 ;
        RECT -18.965 5.460 -18.795 5.785 ;
        RECT -18.615 5.685 -18.245 6.025 ;
        RECT -18.065 5.785 -17.515 5.955 ;
        RECT -13.465 5.785 -12.915 5.955 ;
        RECT -18.065 5.460 -17.895 5.785 ;
        RECT -18.965 5.290 -17.895 5.460 ;
        RECT -13.085 5.460 -12.915 5.785 ;
        RECT -12.735 5.685 -12.365 6.025 ;
        RECT -12.185 5.785 -11.255 5.965 ;
        RECT -9.805 5.785 -8.875 5.965 ;
        RECT -12.185 5.460 -12.015 5.785 ;
        RECT -13.085 5.290 -12.015 5.460 ;
        RECT -9.045 5.460 -8.875 5.785 ;
        RECT -8.695 5.685 -8.325 6.025 ;
        RECT -8.145 5.785 -7.595 5.955 ;
        RECT -3.545 5.785 -2.995 5.955 ;
        RECT -8.145 5.460 -7.975 5.785 ;
        RECT -9.045 5.290 -7.975 5.460 ;
        RECT -3.165 5.460 -2.995 5.785 ;
        RECT -2.815 5.685 -2.445 6.025 ;
        RECT -2.265 5.785 -1.335 5.965 ;
        RECT 0.115 5.785 1.045 5.965 ;
        RECT -2.265 5.460 -2.095 5.785 ;
        RECT -3.165 5.290 -2.095 5.460 ;
        RECT 0.875 5.460 1.045 5.785 ;
        RECT 1.225 5.685 1.595 6.025 ;
        RECT 1.775 5.785 2.325 5.955 ;
        RECT 6.375 5.785 6.925 5.955 ;
        RECT 1.775 5.460 1.945 5.785 ;
        RECT 0.875 5.290 1.945 5.460 ;
        RECT 6.755 5.460 6.925 5.785 ;
        RECT 7.105 5.685 7.475 6.025 ;
        RECT 7.655 5.785 8.585 5.965 ;
        RECT 10.035 5.785 10.965 5.965 ;
        RECT 7.655 5.460 7.825 5.785 ;
        RECT 6.755 5.290 7.825 5.460 ;
        RECT 10.795 5.460 10.965 5.785 ;
        RECT 11.145 5.685 11.515 6.025 ;
        RECT 11.695 5.785 12.245 5.955 ;
        RECT 16.295 5.785 16.845 5.955 ;
        RECT 11.695 5.460 11.865 5.785 ;
        RECT 10.795 5.290 11.865 5.460 ;
        RECT 16.675 5.460 16.845 5.785 ;
        RECT 17.025 5.685 17.395 6.025 ;
        RECT 17.575 5.785 18.505 5.965 ;
        RECT 19.955 5.785 20.885 5.965 ;
        RECT 17.575 5.460 17.745 5.785 ;
        RECT 16.675 5.290 17.745 5.460 ;
        RECT 20.715 5.460 20.885 5.785 ;
        RECT 21.065 5.685 21.435 6.025 ;
        RECT 21.615 5.785 22.165 5.955 ;
        RECT 21.615 5.460 21.785 5.785 ;
        RECT 22.335 5.605 22.505 6.130 ;
        RECT 20.715 5.290 21.785 5.460 ;
        RECT -291.565 5.090 -291.395 5.275 ;
        RECT -290.420 5.185 -290.090 5.290 ;
        RECT -286.490 5.185 -286.160 5.290 ;
        RECT -280.500 5.185 -280.170 5.290 ;
        RECT -276.570 5.185 -276.240 5.290 ;
        RECT -270.580 5.185 -270.250 5.290 ;
        RECT -266.650 5.185 -266.320 5.290 ;
        RECT -260.660 5.185 -260.330 5.290 ;
        RECT -256.730 5.185 -256.400 5.290 ;
        RECT -250.740 5.185 -250.410 5.290 ;
        RECT -246.810 5.185 -246.480 5.290 ;
        RECT -240.820 5.185 -240.490 5.290 ;
        RECT -236.890 5.185 -236.560 5.290 ;
        RECT -230.900 5.185 -230.570 5.290 ;
        RECT -226.970 5.185 -226.640 5.290 ;
        RECT -220.980 5.185 -220.650 5.290 ;
        RECT -217.050 5.185 -216.720 5.290 ;
        RECT -211.060 5.185 -210.730 5.290 ;
        RECT -207.130 5.185 -206.800 5.290 ;
        RECT -201.140 5.185 -200.810 5.290 ;
        RECT -197.210 5.185 -196.880 5.290 ;
        RECT -191.220 5.185 -190.890 5.290 ;
        RECT -187.290 5.185 -186.960 5.290 ;
        RECT -181.300 5.185 -180.970 5.290 ;
        RECT -177.370 5.185 -177.040 5.290 ;
        RECT -171.380 5.185 -171.050 5.290 ;
        RECT -167.450 5.185 -167.120 5.290 ;
        RECT -161.460 5.185 -161.130 5.290 ;
        RECT -157.530 5.185 -157.200 5.290 ;
        RECT -151.540 5.185 -151.210 5.290 ;
        RECT -147.610 5.185 -147.280 5.290 ;
        RECT -141.620 5.185 -141.290 5.290 ;
        RECT -137.690 5.185 -137.360 5.290 ;
        RECT -131.700 5.185 -131.370 5.290 ;
        RECT -127.770 5.185 -127.440 5.290 ;
        RECT -121.780 5.185 -121.450 5.290 ;
        RECT -117.850 5.185 -117.520 5.290 ;
        RECT -111.860 5.185 -111.530 5.290 ;
        RECT -107.930 5.185 -107.600 5.290 ;
        RECT -101.940 5.185 -101.610 5.290 ;
        RECT -98.010 5.185 -97.680 5.290 ;
        RECT -92.020 5.185 -91.690 5.290 ;
        RECT -88.090 5.185 -87.760 5.290 ;
        RECT -82.100 5.185 -81.770 5.290 ;
        RECT -78.170 5.185 -77.840 5.290 ;
        RECT -72.180 5.185 -71.850 5.290 ;
        RECT -68.250 5.185 -67.920 5.290 ;
        RECT -62.260 5.185 -61.930 5.290 ;
        RECT -58.330 5.185 -58.000 5.290 ;
        RECT -52.340 5.185 -52.010 5.290 ;
        RECT -48.410 5.185 -48.080 5.290 ;
        RECT -42.420 5.185 -42.090 5.290 ;
        RECT -38.490 5.185 -38.160 5.290 ;
        RECT -32.500 5.185 -32.170 5.290 ;
        RECT -28.570 5.185 -28.240 5.290 ;
        RECT -22.580 5.185 -22.250 5.290 ;
        RECT -18.650 5.185 -18.320 5.290 ;
        RECT -12.660 5.185 -12.330 5.290 ;
        RECT -8.730 5.185 -8.400 5.290 ;
        RECT -2.740 5.185 -2.410 5.290 ;
        RECT 1.190 5.185 1.520 5.290 ;
        RECT 7.180 5.185 7.510 5.290 ;
        RECT 11.110 5.185 11.440 5.290 ;
        RECT 17.100 5.185 17.430 5.290 ;
        RECT 21.030 5.185 21.360 5.290 ;
        RECT 21.955 5.275 22.505 5.605 ;
        RECT -292.095 5.075 -291.395 5.090 ;
        RECT -292.180 4.905 -291.395 5.075 ;
        RECT -291.860 4.900 -291.395 4.905 ;
        RECT -291.565 4.750 -291.395 4.900 ;
        RECT -287.565 5.015 -286.660 5.105 ;
        RECT -285.860 5.015 -285.355 5.095 ;
        RECT -287.565 4.835 -285.355 5.015 ;
        RECT -277.645 5.015 -276.740 5.105 ;
        RECT -275.940 5.015 -275.435 5.095 ;
        RECT -277.645 4.835 -275.435 5.015 ;
        RECT -267.725 5.015 -266.820 5.105 ;
        RECT -266.020 5.015 -265.515 5.095 ;
        RECT -267.725 4.835 -265.515 5.015 ;
        RECT -257.805 5.015 -256.900 5.105 ;
        RECT -256.100 5.015 -255.595 5.095 ;
        RECT -257.805 4.835 -255.595 5.015 ;
        RECT -247.885 5.015 -246.980 5.105 ;
        RECT -246.180 5.015 -245.675 5.095 ;
        RECT -247.885 4.835 -245.675 5.015 ;
        RECT -237.965 5.015 -237.060 5.105 ;
        RECT -236.260 5.015 -235.755 5.095 ;
        RECT -237.965 4.835 -235.755 5.015 ;
        RECT -228.045 5.015 -227.140 5.105 ;
        RECT -226.340 5.015 -225.835 5.095 ;
        RECT -228.045 4.835 -225.835 5.015 ;
        RECT -218.125 5.015 -217.220 5.105 ;
        RECT -216.420 5.015 -215.915 5.095 ;
        RECT -218.125 4.835 -215.915 5.015 ;
        RECT -208.205 5.015 -207.300 5.105 ;
        RECT -206.500 5.015 -205.995 5.095 ;
        RECT -208.205 4.835 -205.995 5.015 ;
        RECT -198.285 5.015 -197.380 5.105 ;
        RECT -196.580 5.015 -196.075 5.095 ;
        RECT -198.285 4.835 -196.075 5.015 ;
        RECT -188.365 5.015 -187.460 5.105 ;
        RECT -186.660 5.015 -186.155 5.095 ;
        RECT -188.365 4.835 -186.155 5.015 ;
        RECT -178.445 5.015 -177.540 5.105 ;
        RECT -176.740 5.015 -176.235 5.095 ;
        RECT -178.445 4.835 -176.235 5.015 ;
        RECT -168.525 5.015 -167.620 5.105 ;
        RECT -166.820 5.015 -166.315 5.095 ;
        RECT -168.525 4.835 -166.315 5.015 ;
        RECT -158.605 5.015 -157.700 5.105 ;
        RECT -156.900 5.015 -156.395 5.095 ;
        RECT -158.605 4.835 -156.395 5.015 ;
        RECT -148.685 5.015 -147.780 5.105 ;
        RECT -146.980 5.015 -146.475 5.095 ;
        RECT -148.685 4.835 -146.475 5.015 ;
        RECT -138.765 5.015 -137.860 5.105 ;
        RECT -137.060 5.015 -136.555 5.095 ;
        RECT -138.765 4.835 -136.555 5.015 ;
        RECT -128.845 5.015 -127.940 5.105 ;
        RECT -127.140 5.015 -126.635 5.095 ;
        RECT -128.845 4.835 -126.635 5.015 ;
        RECT -118.925 5.015 -118.020 5.105 ;
        RECT -117.220 5.015 -116.715 5.095 ;
        RECT -118.925 4.835 -116.715 5.015 ;
        RECT -109.005 5.015 -108.100 5.105 ;
        RECT -107.300 5.015 -106.795 5.095 ;
        RECT -109.005 4.835 -106.795 5.015 ;
        RECT -99.085 5.015 -98.180 5.105 ;
        RECT -97.380 5.015 -96.875 5.095 ;
        RECT -99.085 4.835 -96.875 5.015 ;
        RECT -89.165 5.015 -88.260 5.105 ;
        RECT -87.460 5.015 -86.955 5.095 ;
        RECT -89.165 4.835 -86.955 5.015 ;
        RECT -79.245 5.015 -78.340 5.105 ;
        RECT -77.540 5.015 -77.035 5.095 ;
        RECT -79.245 4.835 -77.035 5.015 ;
        RECT -69.325 5.015 -68.420 5.105 ;
        RECT -67.620 5.015 -67.115 5.095 ;
        RECT -69.325 4.835 -67.115 5.015 ;
        RECT -59.405 5.015 -58.500 5.105 ;
        RECT -57.700 5.015 -57.195 5.095 ;
        RECT -59.405 4.835 -57.195 5.015 ;
        RECT -49.485 5.015 -48.580 5.105 ;
        RECT -47.780 5.015 -47.275 5.095 ;
        RECT -49.485 4.835 -47.275 5.015 ;
        RECT -39.565 5.015 -38.660 5.105 ;
        RECT -37.860 5.015 -37.355 5.095 ;
        RECT -39.565 4.835 -37.355 5.015 ;
        RECT -29.645 5.015 -28.740 5.105 ;
        RECT -27.940 5.015 -27.435 5.095 ;
        RECT -29.645 4.835 -27.435 5.015 ;
        RECT -19.725 5.015 -18.820 5.105 ;
        RECT -18.020 5.015 -17.515 5.095 ;
        RECT -19.725 4.835 -17.515 5.015 ;
        RECT -9.805 5.015 -8.900 5.105 ;
        RECT -8.100 5.015 -7.595 5.095 ;
        RECT -9.805 4.835 -7.595 5.015 ;
        RECT 0.115 5.015 1.020 5.105 ;
        RECT 1.820 5.015 2.325 5.095 ;
        RECT 0.115 4.835 2.325 5.015 ;
        RECT 10.035 5.015 10.940 5.105 ;
        RECT 11.740 5.015 12.245 5.095 ;
        RECT 10.035 4.835 12.245 5.015 ;
        RECT 19.955 5.015 20.860 5.105 ;
        RECT 21.660 5.015 22.165 5.095 ;
        RECT 19.955 4.835 22.165 5.015 ;
        RECT 22.335 5.080 22.505 5.275 ;
        RECT 22.745 5.080 23.035 5.800 ;
        RECT 22.335 5.075 23.035 5.080 ;
        RECT 22.335 4.905 23.120 5.075 ;
        RECT 22.335 4.900 22.800 4.905 ;
        RECT 22.335 4.750 22.505 4.900 ;
        RECT -292.505 -78.010 -292.335 -77.860 ;
        RECT -293.120 -78.180 -292.335 -78.010 ;
        RECT -293.035 -79.345 -292.745 -78.180 ;
        RECT -292.505 -78.385 -292.335 -78.180 ;
        RECT -292.165 -78.125 -289.955 -77.945 ;
        RECT -292.165 -78.215 -291.260 -78.125 ;
        RECT -290.460 -78.205 -289.955 -78.125 ;
        RECT -282.245 -78.125 -280.035 -77.945 ;
        RECT -282.245 -78.215 -281.340 -78.125 ;
        RECT -280.540 -78.205 -280.035 -78.125 ;
        RECT -272.325 -78.125 -270.115 -77.945 ;
        RECT -272.325 -78.215 -271.420 -78.125 ;
        RECT -270.620 -78.205 -270.115 -78.125 ;
        RECT -262.405 -78.125 -260.195 -77.945 ;
        RECT -262.405 -78.215 -261.500 -78.125 ;
        RECT -260.700 -78.205 -260.195 -78.125 ;
        RECT -252.485 -78.125 -250.275 -77.945 ;
        RECT -252.485 -78.215 -251.580 -78.125 ;
        RECT -250.780 -78.205 -250.275 -78.125 ;
        RECT -242.565 -78.125 -240.355 -77.945 ;
        RECT -242.565 -78.215 -241.660 -78.125 ;
        RECT -240.860 -78.205 -240.355 -78.125 ;
        RECT -232.645 -78.125 -230.435 -77.945 ;
        RECT -232.645 -78.215 -231.740 -78.125 ;
        RECT -230.940 -78.205 -230.435 -78.125 ;
        RECT -222.725 -78.125 -220.515 -77.945 ;
        RECT -222.725 -78.215 -221.820 -78.125 ;
        RECT -221.020 -78.205 -220.515 -78.125 ;
        RECT -212.805 -78.125 -210.595 -77.945 ;
        RECT -212.805 -78.215 -211.900 -78.125 ;
        RECT -211.100 -78.205 -210.595 -78.125 ;
        RECT -202.885 -78.125 -200.675 -77.945 ;
        RECT -202.885 -78.215 -201.980 -78.125 ;
        RECT -201.180 -78.205 -200.675 -78.125 ;
        RECT -192.965 -78.125 -190.755 -77.945 ;
        RECT -192.965 -78.215 -192.060 -78.125 ;
        RECT -191.260 -78.205 -190.755 -78.125 ;
        RECT -183.045 -78.125 -180.835 -77.945 ;
        RECT -183.045 -78.215 -182.140 -78.125 ;
        RECT -181.340 -78.205 -180.835 -78.125 ;
        RECT -173.125 -78.125 -170.915 -77.945 ;
        RECT -173.125 -78.215 -172.220 -78.125 ;
        RECT -171.420 -78.205 -170.915 -78.125 ;
        RECT -163.205 -78.125 -160.995 -77.945 ;
        RECT -163.205 -78.215 -162.300 -78.125 ;
        RECT -161.500 -78.205 -160.995 -78.125 ;
        RECT -153.285 -78.125 -151.075 -77.945 ;
        RECT -153.285 -78.215 -152.380 -78.125 ;
        RECT -151.580 -78.205 -151.075 -78.125 ;
        RECT -143.365 -78.125 -141.155 -77.945 ;
        RECT -143.365 -78.215 -142.460 -78.125 ;
        RECT -141.660 -78.205 -141.155 -78.125 ;
        RECT -133.445 -78.125 -131.235 -77.945 ;
        RECT -133.445 -78.215 -132.540 -78.125 ;
        RECT -131.740 -78.205 -131.235 -78.125 ;
        RECT -123.525 -78.125 -121.315 -77.945 ;
        RECT -123.525 -78.215 -122.620 -78.125 ;
        RECT -121.820 -78.205 -121.315 -78.125 ;
        RECT -113.605 -78.125 -111.395 -77.945 ;
        RECT -113.605 -78.215 -112.700 -78.125 ;
        RECT -111.900 -78.205 -111.395 -78.125 ;
        RECT -103.685 -78.125 -101.475 -77.945 ;
        RECT -103.685 -78.215 -102.780 -78.125 ;
        RECT -101.980 -78.205 -101.475 -78.125 ;
        RECT -93.765 -78.125 -91.555 -77.945 ;
        RECT -93.765 -78.215 -92.860 -78.125 ;
        RECT -92.060 -78.205 -91.555 -78.125 ;
        RECT -83.845 -78.125 -81.635 -77.945 ;
        RECT -83.845 -78.215 -82.940 -78.125 ;
        RECT -82.140 -78.205 -81.635 -78.125 ;
        RECT -73.925 -78.125 -71.715 -77.945 ;
        RECT -73.925 -78.215 -73.020 -78.125 ;
        RECT -72.220 -78.205 -71.715 -78.125 ;
        RECT -64.005 -78.125 -61.795 -77.945 ;
        RECT -64.005 -78.215 -63.100 -78.125 ;
        RECT -62.300 -78.205 -61.795 -78.125 ;
        RECT -54.085 -78.125 -51.875 -77.945 ;
        RECT -54.085 -78.215 -53.180 -78.125 ;
        RECT -52.380 -78.205 -51.875 -78.125 ;
        RECT -44.165 -78.125 -41.955 -77.945 ;
        RECT -44.165 -78.215 -43.260 -78.125 ;
        RECT -42.460 -78.205 -41.955 -78.125 ;
        RECT -34.245 -78.125 -32.035 -77.945 ;
        RECT -34.245 -78.215 -33.340 -78.125 ;
        RECT -32.540 -78.205 -32.035 -78.125 ;
        RECT -24.325 -78.125 -22.115 -77.945 ;
        RECT -24.325 -78.215 -23.420 -78.125 ;
        RECT -22.620 -78.205 -22.115 -78.125 ;
        RECT -14.405 -78.125 -12.195 -77.945 ;
        RECT -14.405 -78.215 -13.500 -78.125 ;
        RECT -12.700 -78.205 -12.195 -78.125 ;
        RECT -4.485 -78.125 -2.275 -77.945 ;
        RECT -4.485 -78.215 -3.580 -78.125 ;
        RECT -2.780 -78.205 -2.275 -78.125 ;
        RECT 5.435 -78.125 7.645 -77.945 ;
        RECT 5.435 -78.215 6.340 -78.125 ;
        RECT 7.140 -78.205 7.645 -78.125 ;
        RECT 15.355 -78.125 17.565 -77.945 ;
        RECT 15.355 -78.215 16.260 -78.125 ;
        RECT 17.060 -78.205 17.565 -78.125 ;
        RECT -292.505 -78.715 -291.575 -78.385 ;
        RECT -291.090 -78.400 -290.760 -78.295 ;
        RECT -285.100 -78.400 -284.770 -78.295 ;
        RECT -281.170 -78.400 -280.840 -78.295 ;
        RECT -275.180 -78.400 -274.850 -78.295 ;
        RECT -271.250 -78.400 -270.920 -78.295 ;
        RECT -265.260 -78.400 -264.930 -78.295 ;
        RECT -261.330 -78.400 -261.000 -78.295 ;
        RECT -255.340 -78.400 -255.010 -78.295 ;
        RECT -251.410 -78.400 -251.080 -78.295 ;
        RECT -245.420 -78.400 -245.090 -78.295 ;
        RECT -241.490 -78.400 -241.160 -78.295 ;
        RECT -235.500 -78.400 -235.170 -78.295 ;
        RECT -231.570 -78.400 -231.240 -78.295 ;
        RECT -225.580 -78.400 -225.250 -78.295 ;
        RECT -221.650 -78.400 -221.320 -78.295 ;
        RECT -215.660 -78.400 -215.330 -78.295 ;
        RECT -211.730 -78.400 -211.400 -78.295 ;
        RECT -205.740 -78.400 -205.410 -78.295 ;
        RECT -201.810 -78.400 -201.480 -78.295 ;
        RECT -195.820 -78.400 -195.490 -78.295 ;
        RECT -191.890 -78.400 -191.560 -78.295 ;
        RECT -185.900 -78.400 -185.570 -78.295 ;
        RECT -181.970 -78.400 -181.640 -78.295 ;
        RECT -175.980 -78.400 -175.650 -78.295 ;
        RECT -172.050 -78.400 -171.720 -78.295 ;
        RECT -166.060 -78.400 -165.730 -78.295 ;
        RECT -162.130 -78.400 -161.800 -78.295 ;
        RECT -156.140 -78.400 -155.810 -78.295 ;
        RECT -152.210 -78.400 -151.880 -78.295 ;
        RECT -146.220 -78.400 -145.890 -78.295 ;
        RECT -142.290 -78.400 -141.960 -78.295 ;
        RECT -136.300 -78.400 -135.970 -78.295 ;
        RECT -132.370 -78.400 -132.040 -78.295 ;
        RECT -126.380 -78.400 -126.050 -78.295 ;
        RECT -122.450 -78.400 -122.120 -78.295 ;
        RECT -116.460 -78.400 -116.130 -78.295 ;
        RECT -112.530 -78.400 -112.200 -78.295 ;
        RECT -106.540 -78.400 -106.210 -78.295 ;
        RECT -102.610 -78.400 -102.280 -78.295 ;
        RECT -96.620 -78.400 -96.290 -78.295 ;
        RECT -92.690 -78.400 -92.360 -78.295 ;
        RECT -86.700 -78.400 -86.370 -78.295 ;
        RECT -82.770 -78.400 -82.440 -78.295 ;
        RECT -76.780 -78.400 -76.450 -78.295 ;
        RECT -72.850 -78.400 -72.520 -78.295 ;
        RECT -66.860 -78.400 -66.530 -78.295 ;
        RECT -62.930 -78.400 -62.600 -78.295 ;
        RECT -56.940 -78.400 -56.610 -78.295 ;
        RECT -53.010 -78.400 -52.680 -78.295 ;
        RECT -47.020 -78.400 -46.690 -78.295 ;
        RECT -43.090 -78.400 -42.760 -78.295 ;
        RECT -37.100 -78.400 -36.770 -78.295 ;
        RECT -33.170 -78.400 -32.840 -78.295 ;
        RECT -27.180 -78.400 -26.850 -78.295 ;
        RECT -23.250 -78.400 -22.920 -78.295 ;
        RECT -17.260 -78.400 -16.930 -78.295 ;
        RECT -13.330 -78.400 -13.000 -78.295 ;
        RECT -7.340 -78.400 -7.010 -78.295 ;
        RECT -3.410 -78.400 -3.080 -78.295 ;
        RECT 2.580 -78.400 2.910 -78.295 ;
        RECT 6.510 -78.400 6.840 -78.295 ;
        RECT 12.500 -78.400 12.830 -78.295 ;
        RECT 16.430 -78.400 16.760 -78.295 ;
        RECT 22.420 -78.400 22.750 -78.295 ;
        RECT -291.405 -78.570 -290.335 -78.400 ;
        RECT -292.505 -79.240 -292.335 -78.715 ;
        RECT -291.405 -78.895 -291.235 -78.570 ;
        RECT -292.165 -79.075 -291.235 -78.895 ;
        RECT -291.055 -79.135 -290.685 -78.795 ;
        RECT -290.505 -78.895 -290.335 -78.570 ;
        RECT -285.525 -78.570 -284.455 -78.400 ;
        RECT -285.525 -78.895 -285.355 -78.570 ;
        RECT -290.505 -79.065 -289.955 -78.895 ;
        RECT -285.905 -79.065 -285.355 -78.895 ;
        RECT -285.175 -79.135 -284.805 -78.795 ;
        RECT -284.625 -78.895 -284.455 -78.570 ;
        RECT -281.485 -78.570 -280.415 -78.400 ;
        RECT -281.485 -78.895 -281.315 -78.570 ;
        RECT -284.625 -79.075 -283.695 -78.895 ;
        RECT -282.245 -79.075 -281.315 -78.895 ;
        RECT -281.135 -79.135 -280.765 -78.795 ;
        RECT -280.585 -78.895 -280.415 -78.570 ;
        RECT -275.605 -78.570 -274.535 -78.400 ;
        RECT -275.605 -78.895 -275.435 -78.570 ;
        RECT -280.585 -79.065 -280.035 -78.895 ;
        RECT -275.985 -79.065 -275.435 -78.895 ;
        RECT -275.255 -79.135 -274.885 -78.795 ;
        RECT -274.705 -78.895 -274.535 -78.570 ;
        RECT -271.565 -78.570 -270.495 -78.400 ;
        RECT -271.565 -78.895 -271.395 -78.570 ;
        RECT -274.705 -79.075 -273.775 -78.895 ;
        RECT -272.325 -79.075 -271.395 -78.895 ;
        RECT -271.215 -79.135 -270.845 -78.795 ;
        RECT -270.665 -78.895 -270.495 -78.570 ;
        RECT -265.685 -78.570 -264.615 -78.400 ;
        RECT -265.685 -78.895 -265.515 -78.570 ;
        RECT -270.665 -79.065 -270.115 -78.895 ;
        RECT -266.065 -79.065 -265.515 -78.895 ;
        RECT -265.335 -79.135 -264.965 -78.795 ;
        RECT -264.785 -78.895 -264.615 -78.570 ;
        RECT -261.645 -78.570 -260.575 -78.400 ;
        RECT -261.645 -78.895 -261.475 -78.570 ;
        RECT -264.785 -79.075 -263.855 -78.895 ;
        RECT -262.405 -79.075 -261.475 -78.895 ;
        RECT -261.295 -79.135 -260.925 -78.795 ;
        RECT -260.745 -78.895 -260.575 -78.570 ;
        RECT -255.765 -78.570 -254.695 -78.400 ;
        RECT -255.765 -78.895 -255.595 -78.570 ;
        RECT -260.745 -79.065 -260.195 -78.895 ;
        RECT -256.145 -79.065 -255.595 -78.895 ;
        RECT -255.415 -79.135 -255.045 -78.795 ;
        RECT -254.865 -78.895 -254.695 -78.570 ;
        RECT -251.725 -78.570 -250.655 -78.400 ;
        RECT -251.725 -78.895 -251.555 -78.570 ;
        RECT -254.865 -79.075 -253.935 -78.895 ;
        RECT -252.485 -79.075 -251.555 -78.895 ;
        RECT -251.375 -79.135 -251.005 -78.795 ;
        RECT -250.825 -78.895 -250.655 -78.570 ;
        RECT -245.845 -78.570 -244.775 -78.400 ;
        RECT -245.845 -78.895 -245.675 -78.570 ;
        RECT -250.825 -79.065 -250.275 -78.895 ;
        RECT -246.225 -79.065 -245.675 -78.895 ;
        RECT -245.495 -79.135 -245.125 -78.795 ;
        RECT -244.945 -78.895 -244.775 -78.570 ;
        RECT -241.805 -78.570 -240.735 -78.400 ;
        RECT -241.805 -78.895 -241.635 -78.570 ;
        RECT -244.945 -79.075 -244.015 -78.895 ;
        RECT -242.565 -79.075 -241.635 -78.895 ;
        RECT -241.455 -79.135 -241.085 -78.795 ;
        RECT -240.905 -78.895 -240.735 -78.570 ;
        RECT -235.925 -78.570 -234.855 -78.400 ;
        RECT -235.925 -78.895 -235.755 -78.570 ;
        RECT -240.905 -79.065 -240.355 -78.895 ;
        RECT -236.305 -79.065 -235.755 -78.895 ;
        RECT -235.575 -79.135 -235.205 -78.795 ;
        RECT -235.025 -78.895 -234.855 -78.570 ;
        RECT -231.885 -78.570 -230.815 -78.400 ;
        RECT -231.885 -78.895 -231.715 -78.570 ;
        RECT -235.025 -79.075 -234.095 -78.895 ;
        RECT -232.645 -79.075 -231.715 -78.895 ;
        RECT -231.535 -79.135 -231.165 -78.795 ;
        RECT -230.985 -78.895 -230.815 -78.570 ;
        RECT -226.005 -78.570 -224.935 -78.400 ;
        RECT -226.005 -78.895 -225.835 -78.570 ;
        RECT -230.985 -79.065 -230.435 -78.895 ;
        RECT -226.385 -79.065 -225.835 -78.895 ;
        RECT -225.655 -79.135 -225.285 -78.795 ;
        RECT -225.105 -78.895 -224.935 -78.570 ;
        RECT -221.965 -78.570 -220.895 -78.400 ;
        RECT -221.965 -78.895 -221.795 -78.570 ;
        RECT -225.105 -79.075 -224.175 -78.895 ;
        RECT -222.725 -79.075 -221.795 -78.895 ;
        RECT -221.615 -79.135 -221.245 -78.795 ;
        RECT -221.065 -78.895 -220.895 -78.570 ;
        RECT -216.085 -78.570 -215.015 -78.400 ;
        RECT -216.085 -78.895 -215.915 -78.570 ;
        RECT -221.065 -79.065 -220.515 -78.895 ;
        RECT -216.465 -79.065 -215.915 -78.895 ;
        RECT -215.735 -79.135 -215.365 -78.795 ;
        RECT -215.185 -78.895 -215.015 -78.570 ;
        RECT -212.045 -78.570 -210.975 -78.400 ;
        RECT -212.045 -78.895 -211.875 -78.570 ;
        RECT -215.185 -79.075 -214.255 -78.895 ;
        RECT -212.805 -79.075 -211.875 -78.895 ;
        RECT -211.695 -79.135 -211.325 -78.795 ;
        RECT -211.145 -78.895 -210.975 -78.570 ;
        RECT -206.165 -78.570 -205.095 -78.400 ;
        RECT -206.165 -78.895 -205.995 -78.570 ;
        RECT -211.145 -79.065 -210.595 -78.895 ;
        RECT -206.545 -79.065 -205.995 -78.895 ;
        RECT -205.815 -79.135 -205.445 -78.795 ;
        RECT -205.265 -78.895 -205.095 -78.570 ;
        RECT -202.125 -78.570 -201.055 -78.400 ;
        RECT -202.125 -78.895 -201.955 -78.570 ;
        RECT -205.265 -79.075 -204.335 -78.895 ;
        RECT -202.885 -79.075 -201.955 -78.895 ;
        RECT -201.775 -79.135 -201.405 -78.795 ;
        RECT -201.225 -78.895 -201.055 -78.570 ;
        RECT -196.245 -78.570 -195.175 -78.400 ;
        RECT -196.245 -78.895 -196.075 -78.570 ;
        RECT -201.225 -79.065 -200.675 -78.895 ;
        RECT -196.625 -79.065 -196.075 -78.895 ;
        RECT -195.895 -79.135 -195.525 -78.795 ;
        RECT -195.345 -78.895 -195.175 -78.570 ;
        RECT -192.205 -78.570 -191.135 -78.400 ;
        RECT -192.205 -78.895 -192.035 -78.570 ;
        RECT -195.345 -79.075 -194.415 -78.895 ;
        RECT -192.965 -79.075 -192.035 -78.895 ;
        RECT -191.855 -79.135 -191.485 -78.795 ;
        RECT -191.305 -78.895 -191.135 -78.570 ;
        RECT -186.325 -78.570 -185.255 -78.400 ;
        RECT -186.325 -78.895 -186.155 -78.570 ;
        RECT -191.305 -79.065 -190.755 -78.895 ;
        RECT -186.705 -79.065 -186.155 -78.895 ;
        RECT -185.975 -79.135 -185.605 -78.795 ;
        RECT -185.425 -78.895 -185.255 -78.570 ;
        RECT -182.285 -78.570 -181.215 -78.400 ;
        RECT -182.285 -78.895 -182.115 -78.570 ;
        RECT -185.425 -79.075 -184.495 -78.895 ;
        RECT -183.045 -79.075 -182.115 -78.895 ;
        RECT -181.935 -79.135 -181.565 -78.795 ;
        RECT -181.385 -78.895 -181.215 -78.570 ;
        RECT -176.405 -78.570 -175.335 -78.400 ;
        RECT -176.405 -78.895 -176.235 -78.570 ;
        RECT -181.385 -79.065 -180.835 -78.895 ;
        RECT -176.785 -79.065 -176.235 -78.895 ;
        RECT -176.055 -79.135 -175.685 -78.795 ;
        RECT -175.505 -78.895 -175.335 -78.570 ;
        RECT -172.365 -78.570 -171.295 -78.400 ;
        RECT -172.365 -78.895 -172.195 -78.570 ;
        RECT -175.505 -79.075 -174.575 -78.895 ;
        RECT -173.125 -79.075 -172.195 -78.895 ;
        RECT -172.015 -79.135 -171.645 -78.795 ;
        RECT -171.465 -78.895 -171.295 -78.570 ;
        RECT -166.485 -78.570 -165.415 -78.400 ;
        RECT -166.485 -78.895 -166.315 -78.570 ;
        RECT -171.465 -79.065 -170.915 -78.895 ;
        RECT -166.865 -79.065 -166.315 -78.895 ;
        RECT -166.135 -79.135 -165.765 -78.795 ;
        RECT -165.585 -78.895 -165.415 -78.570 ;
        RECT -162.445 -78.570 -161.375 -78.400 ;
        RECT -162.445 -78.895 -162.275 -78.570 ;
        RECT -165.585 -79.075 -164.655 -78.895 ;
        RECT -163.205 -79.075 -162.275 -78.895 ;
        RECT -162.095 -79.135 -161.725 -78.795 ;
        RECT -161.545 -78.895 -161.375 -78.570 ;
        RECT -156.565 -78.570 -155.495 -78.400 ;
        RECT -156.565 -78.895 -156.395 -78.570 ;
        RECT -161.545 -79.065 -160.995 -78.895 ;
        RECT -156.945 -79.065 -156.395 -78.895 ;
        RECT -156.215 -79.135 -155.845 -78.795 ;
        RECT -155.665 -78.895 -155.495 -78.570 ;
        RECT -152.525 -78.570 -151.455 -78.400 ;
        RECT -152.525 -78.895 -152.355 -78.570 ;
        RECT -155.665 -79.075 -154.735 -78.895 ;
        RECT -153.285 -79.075 -152.355 -78.895 ;
        RECT -152.175 -79.135 -151.805 -78.795 ;
        RECT -151.625 -78.895 -151.455 -78.570 ;
        RECT -146.645 -78.570 -145.575 -78.400 ;
        RECT -146.645 -78.895 -146.475 -78.570 ;
        RECT -151.625 -79.065 -151.075 -78.895 ;
        RECT -147.025 -79.065 -146.475 -78.895 ;
        RECT -146.295 -79.135 -145.925 -78.795 ;
        RECT -145.745 -78.895 -145.575 -78.570 ;
        RECT -142.605 -78.570 -141.535 -78.400 ;
        RECT -142.605 -78.895 -142.435 -78.570 ;
        RECT -145.745 -79.075 -144.815 -78.895 ;
        RECT -143.365 -79.075 -142.435 -78.895 ;
        RECT -142.255 -79.135 -141.885 -78.795 ;
        RECT -141.705 -78.895 -141.535 -78.570 ;
        RECT -136.725 -78.570 -135.655 -78.400 ;
        RECT -136.725 -78.895 -136.555 -78.570 ;
        RECT -141.705 -79.065 -141.155 -78.895 ;
        RECT -137.105 -79.065 -136.555 -78.895 ;
        RECT -136.375 -79.135 -136.005 -78.795 ;
        RECT -135.825 -78.895 -135.655 -78.570 ;
        RECT -132.685 -78.570 -131.615 -78.400 ;
        RECT -132.685 -78.895 -132.515 -78.570 ;
        RECT -135.825 -79.075 -134.895 -78.895 ;
        RECT -133.445 -79.075 -132.515 -78.895 ;
        RECT -132.335 -79.135 -131.965 -78.795 ;
        RECT -131.785 -78.895 -131.615 -78.570 ;
        RECT -126.805 -78.570 -125.735 -78.400 ;
        RECT -126.805 -78.895 -126.635 -78.570 ;
        RECT -131.785 -79.065 -131.235 -78.895 ;
        RECT -127.185 -79.065 -126.635 -78.895 ;
        RECT -126.455 -79.135 -126.085 -78.795 ;
        RECT -125.905 -78.895 -125.735 -78.570 ;
        RECT -122.765 -78.570 -121.695 -78.400 ;
        RECT -122.765 -78.895 -122.595 -78.570 ;
        RECT -125.905 -79.075 -124.975 -78.895 ;
        RECT -123.525 -79.075 -122.595 -78.895 ;
        RECT -122.415 -79.135 -122.045 -78.795 ;
        RECT -121.865 -78.895 -121.695 -78.570 ;
        RECT -116.885 -78.570 -115.815 -78.400 ;
        RECT -116.885 -78.895 -116.715 -78.570 ;
        RECT -121.865 -79.065 -121.315 -78.895 ;
        RECT -117.265 -79.065 -116.715 -78.895 ;
        RECT -116.535 -79.135 -116.165 -78.795 ;
        RECT -115.985 -78.895 -115.815 -78.570 ;
        RECT -112.845 -78.570 -111.775 -78.400 ;
        RECT -112.845 -78.895 -112.675 -78.570 ;
        RECT -115.985 -79.075 -115.055 -78.895 ;
        RECT -113.605 -79.075 -112.675 -78.895 ;
        RECT -112.495 -79.135 -112.125 -78.795 ;
        RECT -111.945 -78.895 -111.775 -78.570 ;
        RECT -106.965 -78.570 -105.895 -78.400 ;
        RECT -106.965 -78.895 -106.795 -78.570 ;
        RECT -111.945 -79.065 -111.395 -78.895 ;
        RECT -107.345 -79.065 -106.795 -78.895 ;
        RECT -106.615 -79.135 -106.245 -78.795 ;
        RECT -106.065 -78.895 -105.895 -78.570 ;
        RECT -102.925 -78.570 -101.855 -78.400 ;
        RECT -102.925 -78.895 -102.755 -78.570 ;
        RECT -106.065 -79.075 -105.135 -78.895 ;
        RECT -103.685 -79.075 -102.755 -78.895 ;
        RECT -102.575 -79.135 -102.205 -78.795 ;
        RECT -102.025 -78.895 -101.855 -78.570 ;
        RECT -97.045 -78.570 -95.975 -78.400 ;
        RECT -97.045 -78.895 -96.875 -78.570 ;
        RECT -102.025 -79.065 -101.475 -78.895 ;
        RECT -97.425 -79.065 -96.875 -78.895 ;
        RECT -96.695 -79.135 -96.325 -78.795 ;
        RECT -96.145 -78.895 -95.975 -78.570 ;
        RECT -93.005 -78.570 -91.935 -78.400 ;
        RECT -93.005 -78.895 -92.835 -78.570 ;
        RECT -96.145 -79.075 -95.215 -78.895 ;
        RECT -93.765 -79.075 -92.835 -78.895 ;
        RECT -92.655 -79.135 -92.285 -78.795 ;
        RECT -92.105 -78.895 -91.935 -78.570 ;
        RECT -87.125 -78.570 -86.055 -78.400 ;
        RECT -87.125 -78.895 -86.955 -78.570 ;
        RECT -92.105 -79.065 -91.555 -78.895 ;
        RECT -87.505 -79.065 -86.955 -78.895 ;
        RECT -86.775 -79.135 -86.405 -78.795 ;
        RECT -86.225 -78.895 -86.055 -78.570 ;
        RECT -83.085 -78.570 -82.015 -78.400 ;
        RECT -83.085 -78.895 -82.915 -78.570 ;
        RECT -86.225 -79.075 -85.295 -78.895 ;
        RECT -83.845 -79.075 -82.915 -78.895 ;
        RECT -82.735 -79.135 -82.365 -78.795 ;
        RECT -82.185 -78.895 -82.015 -78.570 ;
        RECT -77.205 -78.570 -76.135 -78.400 ;
        RECT -77.205 -78.895 -77.035 -78.570 ;
        RECT -82.185 -79.065 -81.635 -78.895 ;
        RECT -77.585 -79.065 -77.035 -78.895 ;
        RECT -76.855 -79.135 -76.485 -78.795 ;
        RECT -76.305 -78.895 -76.135 -78.570 ;
        RECT -73.165 -78.570 -72.095 -78.400 ;
        RECT -73.165 -78.895 -72.995 -78.570 ;
        RECT -76.305 -79.075 -75.375 -78.895 ;
        RECT -73.925 -79.075 -72.995 -78.895 ;
        RECT -72.815 -79.135 -72.445 -78.795 ;
        RECT -72.265 -78.895 -72.095 -78.570 ;
        RECT -67.285 -78.570 -66.215 -78.400 ;
        RECT -67.285 -78.895 -67.115 -78.570 ;
        RECT -72.265 -79.065 -71.715 -78.895 ;
        RECT -67.665 -79.065 -67.115 -78.895 ;
        RECT -66.935 -79.135 -66.565 -78.795 ;
        RECT -66.385 -78.895 -66.215 -78.570 ;
        RECT -63.245 -78.570 -62.175 -78.400 ;
        RECT -63.245 -78.895 -63.075 -78.570 ;
        RECT -66.385 -79.075 -65.455 -78.895 ;
        RECT -64.005 -79.075 -63.075 -78.895 ;
        RECT -62.895 -79.135 -62.525 -78.795 ;
        RECT -62.345 -78.895 -62.175 -78.570 ;
        RECT -57.365 -78.570 -56.295 -78.400 ;
        RECT -57.365 -78.895 -57.195 -78.570 ;
        RECT -62.345 -79.065 -61.795 -78.895 ;
        RECT -57.745 -79.065 -57.195 -78.895 ;
        RECT -57.015 -79.135 -56.645 -78.795 ;
        RECT -56.465 -78.895 -56.295 -78.570 ;
        RECT -53.325 -78.570 -52.255 -78.400 ;
        RECT -53.325 -78.895 -53.155 -78.570 ;
        RECT -56.465 -79.075 -55.535 -78.895 ;
        RECT -54.085 -79.075 -53.155 -78.895 ;
        RECT -52.975 -79.135 -52.605 -78.795 ;
        RECT -52.425 -78.895 -52.255 -78.570 ;
        RECT -47.445 -78.570 -46.375 -78.400 ;
        RECT -47.445 -78.895 -47.275 -78.570 ;
        RECT -52.425 -79.065 -51.875 -78.895 ;
        RECT -47.825 -79.065 -47.275 -78.895 ;
        RECT -47.095 -79.135 -46.725 -78.795 ;
        RECT -46.545 -78.895 -46.375 -78.570 ;
        RECT -43.405 -78.570 -42.335 -78.400 ;
        RECT -43.405 -78.895 -43.235 -78.570 ;
        RECT -46.545 -79.075 -45.615 -78.895 ;
        RECT -44.165 -79.075 -43.235 -78.895 ;
        RECT -43.055 -79.135 -42.685 -78.795 ;
        RECT -42.505 -78.895 -42.335 -78.570 ;
        RECT -37.525 -78.570 -36.455 -78.400 ;
        RECT -37.525 -78.895 -37.355 -78.570 ;
        RECT -42.505 -79.065 -41.955 -78.895 ;
        RECT -37.905 -79.065 -37.355 -78.895 ;
        RECT -37.175 -79.135 -36.805 -78.795 ;
        RECT -36.625 -78.895 -36.455 -78.570 ;
        RECT -33.485 -78.570 -32.415 -78.400 ;
        RECT -33.485 -78.895 -33.315 -78.570 ;
        RECT -36.625 -79.075 -35.695 -78.895 ;
        RECT -34.245 -79.075 -33.315 -78.895 ;
        RECT -33.135 -79.135 -32.765 -78.795 ;
        RECT -32.585 -78.895 -32.415 -78.570 ;
        RECT -27.605 -78.570 -26.535 -78.400 ;
        RECT -27.605 -78.895 -27.435 -78.570 ;
        RECT -32.585 -79.065 -32.035 -78.895 ;
        RECT -27.985 -79.065 -27.435 -78.895 ;
        RECT -27.255 -79.135 -26.885 -78.795 ;
        RECT -26.705 -78.895 -26.535 -78.570 ;
        RECT -23.565 -78.570 -22.495 -78.400 ;
        RECT -23.565 -78.895 -23.395 -78.570 ;
        RECT -26.705 -79.075 -25.775 -78.895 ;
        RECT -24.325 -79.075 -23.395 -78.895 ;
        RECT -23.215 -79.135 -22.845 -78.795 ;
        RECT -22.665 -78.895 -22.495 -78.570 ;
        RECT -17.685 -78.570 -16.615 -78.400 ;
        RECT -17.685 -78.895 -17.515 -78.570 ;
        RECT -22.665 -79.065 -22.115 -78.895 ;
        RECT -18.065 -79.065 -17.515 -78.895 ;
        RECT -17.335 -79.135 -16.965 -78.795 ;
        RECT -16.785 -78.895 -16.615 -78.570 ;
        RECT -13.645 -78.570 -12.575 -78.400 ;
        RECT -13.645 -78.895 -13.475 -78.570 ;
        RECT -16.785 -79.075 -15.855 -78.895 ;
        RECT -14.405 -79.075 -13.475 -78.895 ;
        RECT -13.295 -79.135 -12.925 -78.795 ;
        RECT -12.745 -78.895 -12.575 -78.570 ;
        RECT -7.765 -78.570 -6.695 -78.400 ;
        RECT -7.765 -78.895 -7.595 -78.570 ;
        RECT -12.745 -79.065 -12.195 -78.895 ;
        RECT -8.145 -79.065 -7.595 -78.895 ;
        RECT -7.415 -79.135 -7.045 -78.795 ;
        RECT -6.865 -78.895 -6.695 -78.570 ;
        RECT -3.725 -78.570 -2.655 -78.400 ;
        RECT -3.725 -78.895 -3.555 -78.570 ;
        RECT -6.865 -79.075 -5.935 -78.895 ;
        RECT -4.485 -79.075 -3.555 -78.895 ;
        RECT -3.375 -79.135 -3.005 -78.795 ;
        RECT -2.825 -78.895 -2.655 -78.570 ;
        RECT 2.155 -78.570 3.225 -78.400 ;
        RECT 2.155 -78.895 2.325 -78.570 ;
        RECT -2.825 -79.065 -2.275 -78.895 ;
        RECT 1.775 -79.065 2.325 -78.895 ;
        RECT 2.505 -79.135 2.875 -78.795 ;
        RECT 3.055 -78.895 3.225 -78.570 ;
        RECT 6.195 -78.570 7.265 -78.400 ;
        RECT 6.195 -78.895 6.365 -78.570 ;
        RECT 3.055 -79.075 3.985 -78.895 ;
        RECT 5.435 -79.075 6.365 -78.895 ;
        RECT 6.545 -79.135 6.915 -78.795 ;
        RECT 7.095 -78.895 7.265 -78.570 ;
        RECT 12.075 -78.570 13.145 -78.400 ;
        RECT 12.075 -78.895 12.245 -78.570 ;
        RECT 7.095 -79.065 7.645 -78.895 ;
        RECT 11.695 -79.065 12.245 -78.895 ;
        RECT 12.425 -79.135 12.795 -78.795 ;
        RECT 12.975 -78.895 13.145 -78.570 ;
        RECT 16.115 -78.570 17.185 -78.400 ;
        RECT 16.115 -78.895 16.285 -78.570 ;
        RECT 12.975 -79.075 13.905 -78.895 ;
        RECT 15.355 -79.075 16.285 -78.895 ;
        RECT 16.465 -79.135 16.835 -78.795 ;
        RECT 17.015 -78.895 17.185 -78.570 ;
        RECT 21.995 -78.570 23.065 -78.400 ;
        RECT 21.995 -78.895 22.165 -78.570 ;
        RECT 17.015 -79.065 17.565 -78.895 ;
        RECT 21.615 -79.065 22.165 -78.895 ;
        RECT 22.345 -79.135 22.715 -78.795 ;
        RECT 22.895 -78.895 23.065 -78.570 ;
        RECT 22.895 -79.075 23.825 -78.895 ;
        RECT -293.120 -79.755 -291.280 -79.585 ;
        RECT 22.940 -79.755 24.780 -79.585 ;
        RECT -293.035 -80.480 -292.745 -79.755 ;
        RECT -292.575 -80.555 -292.265 -79.755 ;
        RECT -292.060 -80.555 -291.365 -79.925 ;
        RECT -293.035 -82.305 -292.745 -81.140 ;
        RECT -292.060 -81.155 -291.890 -80.555 ;
        RECT -291.720 -80.995 -291.385 -80.745 ;
        RECT -289.025 -80.905 -288.695 -79.925 ;
        RECT -287.165 -80.905 -286.835 -79.925 ;
        RECT -284.495 -80.555 -283.800 -79.925 ;
        RECT -292.575 -82.305 -292.295 -81.165 ;
        RECT -292.125 -82.135 -291.795 -81.155 ;
        RECT -291.625 -82.305 -291.365 -81.165 ;
        RECT -289.435 -81.315 -289.100 -81.065 ;
        RECT -288.930 -81.505 -288.760 -80.905 ;
        RECT -289.455 -82.135 -288.760 -81.505 ;
        RECT -287.100 -81.505 -286.930 -80.905 ;
        RECT -284.475 -80.995 -284.140 -80.745 ;
        RECT -286.760 -81.315 -286.425 -81.065 ;
        RECT -283.970 -81.155 -283.800 -80.555 ;
        RECT -282.140 -80.555 -281.445 -79.925 ;
        RECT -282.140 -81.155 -281.970 -80.555 ;
        RECT -281.800 -80.995 -281.465 -80.745 ;
        RECT -279.105 -80.905 -278.775 -79.925 ;
        RECT -277.245 -80.905 -276.915 -79.925 ;
        RECT -274.575 -80.555 -273.880 -79.925 ;
        RECT -287.100 -82.135 -286.405 -81.505 ;
        RECT -284.065 -82.135 -283.735 -81.155 ;
        RECT -282.205 -82.135 -281.875 -81.155 ;
        RECT -279.515 -81.315 -279.180 -81.065 ;
        RECT -279.010 -81.505 -278.840 -80.905 ;
        RECT -279.535 -82.135 -278.840 -81.505 ;
        RECT -277.180 -81.505 -277.010 -80.905 ;
        RECT -274.555 -80.995 -274.220 -80.745 ;
        RECT -276.840 -81.315 -276.505 -81.065 ;
        RECT -274.050 -81.155 -273.880 -80.555 ;
        RECT -272.220 -80.555 -271.525 -79.925 ;
        RECT -272.220 -81.155 -272.050 -80.555 ;
        RECT -271.880 -80.995 -271.545 -80.745 ;
        RECT -269.185 -80.905 -268.855 -79.925 ;
        RECT -267.325 -80.905 -266.995 -79.925 ;
        RECT -264.655 -80.555 -263.960 -79.925 ;
        RECT -277.180 -82.135 -276.485 -81.505 ;
        RECT -274.145 -82.135 -273.815 -81.155 ;
        RECT -272.285 -82.135 -271.955 -81.155 ;
        RECT -269.595 -81.315 -269.260 -81.065 ;
        RECT -269.090 -81.505 -268.920 -80.905 ;
        RECT -269.615 -82.135 -268.920 -81.505 ;
        RECT -267.260 -81.505 -267.090 -80.905 ;
        RECT -264.635 -80.995 -264.300 -80.745 ;
        RECT -266.920 -81.315 -266.585 -81.065 ;
        RECT -264.130 -81.155 -263.960 -80.555 ;
        RECT -262.300 -80.555 -261.605 -79.925 ;
        RECT -262.300 -81.155 -262.130 -80.555 ;
        RECT -261.960 -80.995 -261.625 -80.745 ;
        RECT -259.265 -80.905 -258.935 -79.925 ;
        RECT -257.405 -80.905 -257.075 -79.925 ;
        RECT -254.735 -80.555 -254.040 -79.925 ;
        RECT -267.260 -82.135 -266.565 -81.505 ;
        RECT -264.225 -82.135 -263.895 -81.155 ;
        RECT -262.365 -82.135 -262.035 -81.155 ;
        RECT -259.675 -81.315 -259.340 -81.065 ;
        RECT -259.170 -81.505 -259.000 -80.905 ;
        RECT -259.695 -82.135 -259.000 -81.505 ;
        RECT -257.340 -81.505 -257.170 -80.905 ;
        RECT -254.715 -80.995 -254.380 -80.745 ;
        RECT -257.000 -81.315 -256.665 -81.065 ;
        RECT -254.210 -81.155 -254.040 -80.555 ;
        RECT -252.380 -80.555 -251.685 -79.925 ;
        RECT -252.380 -81.155 -252.210 -80.555 ;
        RECT -252.040 -80.995 -251.705 -80.745 ;
        RECT -249.345 -80.905 -249.015 -79.925 ;
        RECT -247.485 -80.905 -247.155 -79.925 ;
        RECT -244.815 -80.555 -244.120 -79.925 ;
        RECT -257.340 -82.135 -256.645 -81.505 ;
        RECT -254.305 -82.135 -253.975 -81.155 ;
        RECT -252.445 -82.135 -252.115 -81.155 ;
        RECT -249.755 -81.315 -249.420 -81.065 ;
        RECT -249.250 -81.505 -249.080 -80.905 ;
        RECT -249.775 -82.135 -249.080 -81.505 ;
        RECT -247.420 -81.505 -247.250 -80.905 ;
        RECT -244.795 -80.995 -244.460 -80.745 ;
        RECT -247.080 -81.315 -246.745 -81.065 ;
        RECT -244.290 -81.155 -244.120 -80.555 ;
        RECT -242.460 -80.555 -241.765 -79.925 ;
        RECT -242.460 -81.155 -242.290 -80.555 ;
        RECT -242.120 -80.995 -241.785 -80.745 ;
        RECT -239.425 -80.905 -239.095 -79.925 ;
        RECT -237.565 -80.905 -237.235 -79.925 ;
        RECT -234.895 -80.555 -234.200 -79.925 ;
        RECT -247.420 -82.135 -246.725 -81.505 ;
        RECT -244.385 -82.135 -244.055 -81.155 ;
        RECT -242.525 -82.135 -242.195 -81.155 ;
        RECT -239.835 -81.315 -239.500 -81.065 ;
        RECT -239.330 -81.505 -239.160 -80.905 ;
        RECT -239.855 -82.135 -239.160 -81.505 ;
        RECT -237.500 -81.505 -237.330 -80.905 ;
        RECT -234.875 -80.995 -234.540 -80.745 ;
        RECT -237.160 -81.315 -236.825 -81.065 ;
        RECT -234.370 -81.155 -234.200 -80.555 ;
        RECT -232.540 -80.555 -231.845 -79.925 ;
        RECT -232.540 -81.155 -232.370 -80.555 ;
        RECT -232.200 -80.995 -231.865 -80.745 ;
        RECT -229.505 -80.905 -229.175 -79.925 ;
        RECT -227.645 -80.905 -227.315 -79.925 ;
        RECT -224.975 -80.555 -224.280 -79.925 ;
        RECT -237.500 -82.135 -236.805 -81.505 ;
        RECT -234.465 -82.135 -234.135 -81.155 ;
        RECT -232.605 -82.135 -232.275 -81.155 ;
        RECT -229.915 -81.315 -229.580 -81.065 ;
        RECT -229.410 -81.505 -229.240 -80.905 ;
        RECT -229.935 -82.135 -229.240 -81.505 ;
        RECT -227.580 -81.505 -227.410 -80.905 ;
        RECT -224.955 -80.995 -224.620 -80.745 ;
        RECT -227.240 -81.315 -226.905 -81.065 ;
        RECT -224.450 -81.155 -224.280 -80.555 ;
        RECT -222.620 -80.555 -221.925 -79.925 ;
        RECT -222.620 -81.155 -222.450 -80.555 ;
        RECT -222.280 -80.995 -221.945 -80.745 ;
        RECT -219.585 -80.905 -219.255 -79.925 ;
        RECT -217.725 -80.905 -217.395 -79.925 ;
        RECT -215.055 -80.555 -214.360 -79.925 ;
        RECT -227.580 -82.135 -226.885 -81.505 ;
        RECT -224.545 -82.135 -224.215 -81.155 ;
        RECT -222.685 -82.135 -222.355 -81.155 ;
        RECT -219.995 -81.315 -219.660 -81.065 ;
        RECT -219.490 -81.505 -219.320 -80.905 ;
        RECT -220.015 -82.135 -219.320 -81.505 ;
        RECT -217.660 -81.505 -217.490 -80.905 ;
        RECT -215.035 -80.995 -214.700 -80.745 ;
        RECT -217.320 -81.315 -216.985 -81.065 ;
        RECT -214.530 -81.155 -214.360 -80.555 ;
        RECT -212.700 -80.555 -212.005 -79.925 ;
        RECT -212.700 -81.155 -212.530 -80.555 ;
        RECT -212.360 -80.995 -212.025 -80.745 ;
        RECT -209.665 -80.905 -209.335 -79.925 ;
        RECT -207.805 -80.905 -207.475 -79.925 ;
        RECT -205.135 -80.555 -204.440 -79.925 ;
        RECT -217.660 -82.135 -216.965 -81.505 ;
        RECT -214.625 -82.135 -214.295 -81.155 ;
        RECT -212.765 -82.135 -212.435 -81.155 ;
        RECT -210.075 -81.315 -209.740 -81.065 ;
        RECT -209.570 -81.505 -209.400 -80.905 ;
        RECT -210.095 -82.135 -209.400 -81.505 ;
        RECT -207.740 -81.505 -207.570 -80.905 ;
        RECT -205.115 -80.995 -204.780 -80.745 ;
        RECT -207.400 -81.315 -207.065 -81.065 ;
        RECT -204.610 -81.155 -204.440 -80.555 ;
        RECT -202.780 -80.555 -202.085 -79.925 ;
        RECT -202.780 -81.155 -202.610 -80.555 ;
        RECT -202.440 -80.995 -202.105 -80.745 ;
        RECT -199.745 -80.905 -199.415 -79.925 ;
        RECT -197.885 -80.905 -197.555 -79.925 ;
        RECT -195.215 -80.555 -194.520 -79.925 ;
        RECT -207.740 -82.135 -207.045 -81.505 ;
        RECT -204.705 -82.135 -204.375 -81.155 ;
        RECT -202.845 -82.135 -202.515 -81.155 ;
        RECT -200.155 -81.315 -199.820 -81.065 ;
        RECT -199.650 -81.505 -199.480 -80.905 ;
        RECT -200.175 -82.135 -199.480 -81.505 ;
        RECT -197.820 -81.505 -197.650 -80.905 ;
        RECT -195.195 -80.995 -194.860 -80.745 ;
        RECT -197.480 -81.315 -197.145 -81.065 ;
        RECT -194.690 -81.155 -194.520 -80.555 ;
        RECT -192.860 -80.555 -192.165 -79.925 ;
        RECT -192.860 -81.155 -192.690 -80.555 ;
        RECT -192.520 -80.995 -192.185 -80.745 ;
        RECT -189.825 -80.905 -189.495 -79.925 ;
        RECT -187.965 -80.905 -187.635 -79.925 ;
        RECT -185.295 -80.555 -184.600 -79.925 ;
        RECT -197.820 -82.135 -197.125 -81.505 ;
        RECT -194.785 -82.135 -194.455 -81.155 ;
        RECT -192.925 -82.135 -192.595 -81.155 ;
        RECT -190.235 -81.315 -189.900 -81.065 ;
        RECT -189.730 -81.505 -189.560 -80.905 ;
        RECT -190.255 -82.135 -189.560 -81.505 ;
        RECT -187.900 -81.505 -187.730 -80.905 ;
        RECT -185.275 -80.995 -184.940 -80.745 ;
        RECT -187.560 -81.315 -187.225 -81.065 ;
        RECT -184.770 -81.155 -184.600 -80.555 ;
        RECT -182.940 -80.555 -182.245 -79.925 ;
        RECT -182.940 -81.155 -182.770 -80.555 ;
        RECT -182.600 -80.995 -182.265 -80.745 ;
        RECT -179.905 -80.905 -179.575 -79.925 ;
        RECT -178.045 -80.905 -177.715 -79.925 ;
        RECT -175.375 -80.555 -174.680 -79.925 ;
        RECT -187.900 -82.135 -187.205 -81.505 ;
        RECT -184.865 -82.135 -184.535 -81.155 ;
        RECT -183.005 -82.135 -182.675 -81.155 ;
        RECT -180.315 -81.315 -179.980 -81.065 ;
        RECT -179.810 -81.505 -179.640 -80.905 ;
        RECT -180.335 -82.135 -179.640 -81.505 ;
        RECT -177.980 -81.505 -177.810 -80.905 ;
        RECT -175.355 -80.995 -175.020 -80.745 ;
        RECT -177.640 -81.315 -177.305 -81.065 ;
        RECT -174.850 -81.155 -174.680 -80.555 ;
        RECT -173.020 -80.555 -172.325 -79.925 ;
        RECT -173.020 -81.155 -172.850 -80.555 ;
        RECT -172.680 -80.995 -172.345 -80.745 ;
        RECT -169.985 -80.905 -169.655 -79.925 ;
        RECT -168.125 -80.905 -167.795 -79.925 ;
        RECT -165.455 -80.555 -164.760 -79.925 ;
        RECT -177.980 -82.135 -177.285 -81.505 ;
        RECT -174.945 -82.135 -174.615 -81.155 ;
        RECT -173.085 -82.135 -172.755 -81.155 ;
        RECT -170.395 -81.315 -170.060 -81.065 ;
        RECT -169.890 -81.505 -169.720 -80.905 ;
        RECT -170.415 -82.135 -169.720 -81.505 ;
        RECT -168.060 -81.505 -167.890 -80.905 ;
        RECT -165.435 -80.995 -165.100 -80.745 ;
        RECT -167.720 -81.315 -167.385 -81.065 ;
        RECT -164.930 -81.155 -164.760 -80.555 ;
        RECT -163.100 -80.555 -162.405 -79.925 ;
        RECT -163.100 -81.155 -162.930 -80.555 ;
        RECT -162.760 -80.995 -162.425 -80.745 ;
        RECT -160.065 -80.905 -159.735 -79.925 ;
        RECT -158.205 -80.905 -157.875 -79.925 ;
        RECT -155.535 -80.555 -154.840 -79.925 ;
        RECT -168.060 -82.135 -167.365 -81.505 ;
        RECT -165.025 -82.135 -164.695 -81.155 ;
        RECT -163.165 -82.135 -162.835 -81.155 ;
        RECT -160.475 -81.315 -160.140 -81.065 ;
        RECT -159.970 -81.505 -159.800 -80.905 ;
        RECT -160.495 -82.135 -159.800 -81.505 ;
        RECT -158.140 -81.505 -157.970 -80.905 ;
        RECT -155.515 -80.995 -155.180 -80.745 ;
        RECT -157.800 -81.315 -157.465 -81.065 ;
        RECT -155.010 -81.155 -154.840 -80.555 ;
        RECT -153.180 -80.555 -152.485 -79.925 ;
        RECT -153.180 -81.155 -153.010 -80.555 ;
        RECT -152.840 -80.995 -152.505 -80.745 ;
        RECT -150.145 -80.905 -149.815 -79.925 ;
        RECT -148.285 -80.905 -147.955 -79.925 ;
        RECT -145.615 -80.555 -144.920 -79.925 ;
        RECT -158.140 -82.135 -157.445 -81.505 ;
        RECT -155.105 -82.135 -154.775 -81.155 ;
        RECT -153.245 -82.135 -152.915 -81.155 ;
        RECT -150.555 -81.315 -150.220 -81.065 ;
        RECT -150.050 -81.505 -149.880 -80.905 ;
        RECT -150.575 -82.135 -149.880 -81.505 ;
        RECT -148.220 -81.505 -148.050 -80.905 ;
        RECT -145.595 -80.995 -145.260 -80.745 ;
        RECT -147.880 -81.315 -147.545 -81.065 ;
        RECT -145.090 -81.155 -144.920 -80.555 ;
        RECT -143.260 -80.555 -142.565 -79.925 ;
        RECT -143.260 -81.155 -143.090 -80.555 ;
        RECT -142.920 -80.995 -142.585 -80.745 ;
        RECT -140.225 -80.905 -139.895 -79.925 ;
        RECT -138.365 -80.905 -138.035 -79.925 ;
        RECT -135.695 -80.555 -135.000 -79.925 ;
        RECT -148.220 -82.135 -147.525 -81.505 ;
        RECT -145.185 -82.135 -144.855 -81.155 ;
        RECT -143.325 -82.135 -142.995 -81.155 ;
        RECT -140.635 -81.315 -140.300 -81.065 ;
        RECT -140.130 -81.505 -139.960 -80.905 ;
        RECT -140.655 -82.135 -139.960 -81.505 ;
        RECT -138.300 -81.505 -138.130 -80.905 ;
        RECT -135.675 -80.995 -135.340 -80.745 ;
        RECT -137.960 -81.315 -137.625 -81.065 ;
        RECT -135.170 -81.155 -135.000 -80.555 ;
        RECT -133.340 -80.555 -132.645 -79.925 ;
        RECT -133.340 -81.155 -133.170 -80.555 ;
        RECT -133.000 -80.995 -132.665 -80.745 ;
        RECT -130.305 -80.905 -129.975 -79.925 ;
        RECT -128.445 -80.905 -128.115 -79.925 ;
        RECT -125.775 -80.555 -125.080 -79.925 ;
        RECT -138.300 -82.135 -137.605 -81.505 ;
        RECT -135.265 -82.135 -134.935 -81.155 ;
        RECT -133.405 -82.135 -133.075 -81.155 ;
        RECT -130.715 -81.315 -130.380 -81.065 ;
        RECT -130.210 -81.505 -130.040 -80.905 ;
        RECT -130.735 -82.135 -130.040 -81.505 ;
        RECT -128.380 -81.505 -128.210 -80.905 ;
        RECT -125.755 -80.995 -125.420 -80.745 ;
        RECT -128.040 -81.315 -127.705 -81.065 ;
        RECT -125.250 -81.155 -125.080 -80.555 ;
        RECT -123.420 -80.555 -122.725 -79.925 ;
        RECT -123.420 -81.155 -123.250 -80.555 ;
        RECT -123.080 -80.995 -122.745 -80.745 ;
        RECT -120.385 -80.905 -120.055 -79.925 ;
        RECT -118.525 -80.905 -118.195 -79.925 ;
        RECT -115.855 -80.555 -115.160 -79.925 ;
        RECT -128.380 -82.135 -127.685 -81.505 ;
        RECT -125.345 -82.135 -125.015 -81.155 ;
        RECT -123.485 -82.135 -123.155 -81.155 ;
        RECT -120.795 -81.315 -120.460 -81.065 ;
        RECT -120.290 -81.505 -120.120 -80.905 ;
        RECT -120.815 -82.135 -120.120 -81.505 ;
        RECT -118.460 -81.505 -118.290 -80.905 ;
        RECT -115.835 -80.995 -115.500 -80.745 ;
        RECT -118.120 -81.315 -117.785 -81.065 ;
        RECT -115.330 -81.155 -115.160 -80.555 ;
        RECT -113.500 -80.555 -112.805 -79.925 ;
        RECT -113.500 -81.155 -113.330 -80.555 ;
        RECT -113.160 -80.995 -112.825 -80.745 ;
        RECT -110.465 -80.905 -110.135 -79.925 ;
        RECT -108.605 -80.905 -108.275 -79.925 ;
        RECT -105.935 -80.555 -105.240 -79.925 ;
        RECT -118.460 -82.135 -117.765 -81.505 ;
        RECT -115.425 -82.135 -115.095 -81.155 ;
        RECT -113.565 -82.135 -113.235 -81.155 ;
        RECT -110.875 -81.315 -110.540 -81.065 ;
        RECT -110.370 -81.505 -110.200 -80.905 ;
        RECT -110.895 -82.135 -110.200 -81.505 ;
        RECT -108.540 -81.505 -108.370 -80.905 ;
        RECT -105.915 -80.995 -105.580 -80.745 ;
        RECT -108.200 -81.315 -107.865 -81.065 ;
        RECT -105.410 -81.155 -105.240 -80.555 ;
        RECT -103.580 -80.555 -102.885 -79.925 ;
        RECT -103.580 -81.155 -103.410 -80.555 ;
        RECT -103.240 -80.995 -102.905 -80.745 ;
        RECT -100.545 -80.905 -100.215 -79.925 ;
        RECT -98.685 -80.905 -98.355 -79.925 ;
        RECT -96.015 -80.555 -95.320 -79.925 ;
        RECT -108.540 -82.135 -107.845 -81.505 ;
        RECT -105.505 -82.135 -105.175 -81.155 ;
        RECT -103.645 -82.135 -103.315 -81.155 ;
        RECT -100.955 -81.315 -100.620 -81.065 ;
        RECT -100.450 -81.505 -100.280 -80.905 ;
        RECT -100.975 -82.135 -100.280 -81.505 ;
        RECT -98.620 -81.505 -98.450 -80.905 ;
        RECT -95.995 -80.995 -95.660 -80.745 ;
        RECT -98.280 -81.315 -97.945 -81.065 ;
        RECT -95.490 -81.155 -95.320 -80.555 ;
        RECT -93.660 -80.555 -92.965 -79.925 ;
        RECT -93.660 -81.155 -93.490 -80.555 ;
        RECT -93.320 -80.995 -92.985 -80.745 ;
        RECT -90.625 -80.905 -90.295 -79.925 ;
        RECT -88.765 -80.905 -88.435 -79.925 ;
        RECT -86.095 -80.555 -85.400 -79.925 ;
        RECT -98.620 -82.135 -97.925 -81.505 ;
        RECT -95.585 -82.135 -95.255 -81.155 ;
        RECT -93.725 -82.135 -93.395 -81.155 ;
        RECT -91.035 -81.315 -90.700 -81.065 ;
        RECT -90.530 -81.505 -90.360 -80.905 ;
        RECT -91.055 -82.135 -90.360 -81.505 ;
        RECT -88.700 -81.505 -88.530 -80.905 ;
        RECT -86.075 -80.995 -85.740 -80.745 ;
        RECT -88.360 -81.315 -88.025 -81.065 ;
        RECT -85.570 -81.155 -85.400 -80.555 ;
        RECT -83.740 -80.555 -83.045 -79.925 ;
        RECT -83.740 -81.155 -83.570 -80.555 ;
        RECT -83.400 -80.995 -83.065 -80.745 ;
        RECT -80.705 -80.905 -80.375 -79.925 ;
        RECT -78.845 -80.905 -78.515 -79.925 ;
        RECT -76.175 -80.555 -75.480 -79.925 ;
        RECT -88.700 -82.135 -88.005 -81.505 ;
        RECT -85.665 -82.135 -85.335 -81.155 ;
        RECT -83.805 -82.135 -83.475 -81.155 ;
        RECT -81.115 -81.315 -80.780 -81.065 ;
        RECT -80.610 -81.505 -80.440 -80.905 ;
        RECT -81.135 -82.135 -80.440 -81.505 ;
        RECT -78.780 -81.505 -78.610 -80.905 ;
        RECT -76.155 -80.995 -75.820 -80.745 ;
        RECT -78.440 -81.315 -78.105 -81.065 ;
        RECT -75.650 -81.155 -75.480 -80.555 ;
        RECT -73.820 -80.555 -73.125 -79.925 ;
        RECT -73.820 -81.155 -73.650 -80.555 ;
        RECT -73.480 -80.995 -73.145 -80.745 ;
        RECT -70.785 -80.905 -70.455 -79.925 ;
        RECT -68.925 -80.905 -68.595 -79.925 ;
        RECT -66.255 -80.555 -65.560 -79.925 ;
        RECT -78.780 -82.135 -78.085 -81.505 ;
        RECT -75.745 -82.135 -75.415 -81.155 ;
        RECT -73.885 -82.135 -73.555 -81.155 ;
        RECT -71.195 -81.315 -70.860 -81.065 ;
        RECT -70.690 -81.505 -70.520 -80.905 ;
        RECT -71.215 -82.135 -70.520 -81.505 ;
        RECT -68.860 -81.505 -68.690 -80.905 ;
        RECT -66.235 -80.995 -65.900 -80.745 ;
        RECT -68.520 -81.315 -68.185 -81.065 ;
        RECT -65.730 -81.155 -65.560 -80.555 ;
        RECT -63.900 -80.555 -63.205 -79.925 ;
        RECT -63.900 -81.155 -63.730 -80.555 ;
        RECT -63.560 -80.995 -63.225 -80.745 ;
        RECT -60.865 -80.905 -60.535 -79.925 ;
        RECT -59.005 -80.905 -58.675 -79.925 ;
        RECT -56.335 -80.555 -55.640 -79.925 ;
        RECT -68.860 -82.135 -68.165 -81.505 ;
        RECT -65.825 -82.135 -65.495 -81.155 ;
        RECT -63.965 -82.135 -63.635 -81.155 ;
        RECT -61.275 -81.315 -60.940 -81.065 ;
        RECT -60.770 -81.505 -60.600 -80.905 ;
        RECT -61.295 -82.135 -60.600 -81.505 ;
        RECT -58.940 -81.505 -58.770 -80.905 ;
        RECT -56.315 -80.995 -55.980 -80.745 ;
        RECT -58.600 -81.315 -58.265 -81.065 ;
        RECT -55.810 -81.155 -55.640 -80.555 ;
        RECT -53.980 -80.555 -53.285 -79.925 ;
        RECT -53.980 -81.155 -53.810 -80.555 ;
        RECT -53.640 -80.995 -53.305 -80.745 ;
        RECT -50.945 -80.905 -50.615 -79.925 ;
        RECT -49.085 -80.905 -48.755 -79.925 ;
        RECT -46.415 -80.555 -45.720 -79.925 ;
        RECT -58.940 -82.135 -58.245 -81.505 ;
        RECT -55.905 -82.135 -55.575 -81.155 ;
        RECT -54.045 -82.135 -53.715 -81.155 ;
        RECT -51.355 -81.315 -51.020 -81.065 ;
        RECT -50.850 -81.505 -50.680 -80.905 ;
        RECT -51.375 -82.135 -50.680 -81.505 ;
        RECT -49.020 -81.505 -48.850 -80.905 ;
        RECT -46.395 -80.995 -46.060 -80.745 ;
        RECT -48.680 -81.315 -48.345 -81.065 ;
        RECT -45.890 -81.155 -45.720 -80.555 ;
        RECT -44.060 -80.555 -43.365 -79.925 ;
        RECT -44.060 -81.155 -43.890 -80.555 ;
        RECT -43.720 -80.995 -43.385 -80.745 ;
        RECT -41.025 -80.905 -40.695 -79.925 ;
        RECT -39.165 -80.905 -38.835 -79.925 ;
        RECT -36.495 -80.555 -35.800 -79.925 ;
        RECT -49.020 -82.135 -48.325 -81.505 ;
        RECT -45.985 -82.135 -45.655 -81.155 ;
        RECT -44.125 -82.135 -43.795 -81.155 ;
        RECT -41.435 -81.315 -41.100 -81.065 ;
        RECT -40.930 -81.505 -40.760 -80.905 ;
        RECT -41.455 -82.135 -40.760 -81.505 ;
        RECT -39.100 -81.505 -38.930 -80.905 ;
        RECT -36.475 -80.995 -36.140 -80.745 ;
        RECT -38.760 -81.315 -38.425 -81.065 ;
        RECT -35.970 -81.155 -35.800 -80.555 ;
        RECT -34.140 -80.555 -33.445 -79.925 ;
        RECT -34.140 -81.155 -33.970 -80.555 ;
        RECT -33.800 -80.995 -33.465 -80.745 ;
        RECT -31.105 -80.905 -30.775 -79.925 ;
        RECT -29.245 -80.905 -28.915 -79.925 ;
        RECT -26.575 -80.555 -25.880 -79.925 ;
        RECT -39.100 -82.135 -38.405 -81.505 ;
        RECT -36.065 -82.135 -35.735 -81.155 ;
        RECT -34.205 -82.135 -33.875 -81.155 ;
        RECT -31.515 -81.315 -31.180 -81.065 ;
        RECT -31.010 -81.505 -30.840 -80.905 ;
        RECT -31.535 -82.135 -30.840 -81.505 ;
        RECT -29.180 -81.505 -29.010 -80.905 ;
        RECT -26.555 -80.995 -26.220 -80.745 ;
        RECT -28.840 -81.315 -28.505 -81.065 ;
        RECT -26.050 -81.155 -25.880 -80.555 ;
        RECT -24.220 -80.555 -23.525 -79.925 ;
        RECT -24.220 -81.155 -24.050 -80.555 ;
        RECT -23.880 -80.995 -23.545 -80.745 ;
        RECT -21.185 -80.905 -20.855 -79.925 ;
        RECT -19.325 -80.905 -18.995 -79.925 ;
        RECT -16.655 -80.555 -15.960 -79.925 ;
        RECT -29.180 -82.135 -28.485 -81.505 ;
        RECT -26.145 -82.135 -25.815 -81.155 ;
        RECT -24.285 -82.135 -23.955 -81.155 ;
        RECT -21.595 -81.315 -21.260 -81.065 ;
        RECT -21.090 -81.505 -20.920 -80.905 ;
        RECT -21.615 -82.135 -20.920 -81.505 ;
        RECT -19.260 -81.505 -19.090 -80.905 ;
        RECT -16.635 -80.995 -16.300 -80.745 ;
        RECT -18.920 -81.315 -18.585 -81.065 ;
        RECT -16.130 -81.155 -15.960 -80.555 ;
        RECT -14.300 -80.555 -13.605 -79.925 ;
        RECT -14.300 -81.155 -14.130 -80.555 ;
        RECT -13.960 -80.995 -13.625 -80.745 ;
        RECT -11.265 -80.905 -10.935 -79.925 ;
        RECT -9.405 -80.905 -9.075 -79.925 ;
        RECT -6.735 -80.555 -6.040 -79.925 ;
        RECT -19.260 -82.135 -18.565 -81.505 ;
        RECT -16.225 -82.135 -15.895 -81.155 ;
        RECT -14.365 -82.135 -14.035 -81.155 ;
        RECT -11.675 -81.315 -11.340 -81.065 ;
        RECT -11.170 -81.505 -11.000 -80.905 ;
        RECT -11.695 -82.135 -11.000 -81.505 ;
        RECT -9.340 -81.505 -9.170 -80.905 ;
        RECT -6.715 -80.995 -6.380 -80.745 ;
        RECT -9.000 -81.315 -8.665 -81.065 ;
        RECT -6.210 -81.155 -6.040 -80.555 ;
        RECT -4.380 -80.555 -3.685 -79.925 ;
        RECT -4.380 -81.155 -4.210 -80.555 ;
        RECT -4.040 -80.995 -3.705 -80.745 ;
        RECT -1.345 -80.905 -1.015 -79.925 ;
        RECT 0.515 -80.905 0.845 -79.925 ;
        RECT 3.185 -80.555 3.880 -79.925 ;
        RECT -9.340 -82.135 -8.645 -81.505 ;
        RECT -6.305 -82.135 -5.975 -81.155 ;
        RECT -4.445 -82.135 -4.115 -81.155 ;
        RECT -1.755 -81.315 -1.420 -81.065 ;
        RECT -1.250 -81.505 -1.080 -80.905 ;
        RECT -1.775 -82.135 -1.080 -81.505 ;
        RECT 0.580 -81.505 0.750 -80.905 ;
        RECT 3.205 -80.995 3.540 -80.745 ;
        RECT 0.920 -81.315 1.255 -81.065 ;
        RECT 3.710 -81.155 3.880 -80.555 ;
        RECT 5.540 -80.555 6.235 -79.925 ;
        RECT 5.540 -81.155 5.710 -80.555 ;
        RECT 5.880 -80.995 6.215 -80.745 ;
        RECT 8.575 -80.905 8.905 -79.925 ;
        RECT 10.435 -80.905 10.765 -79.925 ;
        RECT 13.105 -80.555 13.800 -79.925 ;
        RECT 0.580 -82.135 1.275 -81.505 ;
        RECT 3.615 -82.135 3.945 -81.155 ;
        RECT 5.475 -82.135 5.805 -81.155 ;
        RECT 8.165 -81.315 8.500 -81.065 ;
        RECT 8.670 -81.505 8.840 -80.905 ;
        RECT 8.145 -82.135 8.840 -81.505 ;
        RECT 10.500 -81.505 10.670 -80.905 ;
        RECT 13.125 -80.995 13.460 -80.745 ;
        RECT 10.840 -81.315 11.175 -81.065 ;
        RECT 13.630 -81.155 13.800 -80.555 ;
        RECT 15.460 -80.555 16.155 -79.925 ;
        RECT 15.460 -81.155 15.630 -80.555 ;
        RECT 15.800 -80.995 16.135 -80.745 ;
        RECT 18.495 -80.905 18.825 -79.925 ;
        RECT 20.355 -80.905 20.685 -79.925 ;
        RECT 23.025 -80.555 23.720 -79.925 ;
        RECT 23.925 -80.555 24.235 -79.755 ;
        RECT 24.405 -80.480 24.695 -79.755 ;
        RECT 10.500 -82.135 11.195 -81.505 ;
        RECT 13.535 -82.135 13.865 -81.155 ;
        RECT 15.395 -82.135 15.725 -81.155 ;
        RECT 18.085 -81.315 18.420 -81.065 ;
        RECT 18.590 -81.505 18.760 -80.905 ;
        RECT 18.065 -82.135 18.760 -81.505 ;
        RECT 20.420 -81.505 20.590 -80.905 ;
        RECT 23.045 -80.995 23.380 -80.745 ;
        RECT 20.760 -81.315 21.095 -81.065 ;
        RECT 23.550 -81.155 23.720 -80.555 ;
        RECT 20.420 -82.135 21.115 -81.505 ;
        RECT 23.455 -82.135 23.785 -81.155 ;
        RECT -293.120 -82.475 -291.280 -82.305 ;
        RECT -291.735 -83.860 -291.445 -83.150 ;
        RECT -291.205 -83.345 -291.035 -82.820 ;
        RECT -290.865 -83.165 -290.315 -82.995 ;
        RECT -291.205 -83.675 -290.655 -83.345 ;
        RECT -290.485 -83.490 -290.315 -83.165 ;
        RECT -290.135 -83.265 -289.765 -82.925 ;
        RECT -289.585 -83.165 -288.655 -82.985 ;
        RECT -287.205 -83.165 -286.275 -82.985 ;
        RECT -289.585 -83.490 -289.415 -83.165 ;
        RECT -290.485 -83.660 -289.415 -83.490 ;
        RECT -286.445 -83.490 -286.275 -83.165 ;
        RECT -286.095 -83.265 -285.725 -82.925 ;
        RECT -285.545 -83.165 -284.995 -82.995 ;
        RECT -280.945 -83.165 -280.395 -82.995 ;
        RECT -285.545 -83.490 -285.375 -83.165 ;
        RECT -286.445 -83.660 -285.375 -83.490 ;
        RECT -280.565 -83.490 -280.395 -83.165 ;
        RECT -280.215 -83.265 -279.845 -82.925 ;
        RECT -279.665 -83.165 -278.735 -82.985 ;
        RECT -277.285 -83.165 -276.355 -82.985 ;
        RECT -279.665 -83.490 -279.495 -83.165 ;
        RECT -280.565 -83.660 -279.495 -83.490 ;
        RECT -276.525 -83.490 -276.355 -83.165 ;
        RECT -276.175 -83.265 -275.805 -82.925 ;
        RECT -275.625 -83.165 -275.075 -82.995 ;
        RECT -271.025 -83.165 -270.475 -82.995 ;
        RECT -275.625 -83.490 -275.455 -83.165 ;
        RECT -276.525 -83.660 -275.455 -83.490 ;
        RECT -270.645 -83.490 -270.475 -83.165 ;
        RECT -270.295 -83.265 -269.925 -82.925 ;
        RECT -269.745 -83.165 -268.815 -82.985 ;
        RECT -267.365 -83.165 -266.435 -82.985 ;
        RECT -269.745 -83.490 -269.575 -83.165 ;
        RECT -270.645 -83.660 -269.575 -83.490 ;
        RECT -266.605 -83.490 -266.435 -83.165 ;
        RECT -266.255 -83.265 -265.885 -82.925 ;
        RECT -265.705 -83.165 -265.155 -82.995 ;
        RECT -261.105 -83.165 -260.555 -82.995 ;
        RECT -265.705 -83.490 -265.535 -83.165 ;
        RECT -266.605 -83.660 -265.535 -83.490 ;
        RECT -260.725 -83.490 -260.555 -83.165 ;
        RECT -260.375 -83.265 -260.005 -82.925 ;
        RECT -259.825 -83.165 -258.895 -82.985 ;
        RECT -257.445 -83.165 -256.515 -82.985 ;
        RECT -259.825 -83.490 -259.655 -83.165 ;
        RECT -260.725 -83.660 -259.655 -83.490 ;
        RECT -256.685 -83.490 -256.515 -83.165 ;
        RECT -256.335 -83.265 -255.965 -82.925 ;
        RECT -255.785 -83.165 -255.235 -82.995 ;
        RECT -251.185 -83.165 -250.635 -82.995 ;
        RECT -255.785 -83.490 -255.615 -83.165 ;
        RECT -256.685 -83.660 -255.615 -83.490 ;
        RECT -250.805 -83.490 -250.635 -83.165 ;
        RECT -250.455 -83.265 -250.085 -82.925 ;
        RECT -249.905 -83.165 -248.975 -82.985 ;
        RECT -247.525 -83.165 -246.595 -82.985 ;
        RECT -249.905 -83.490 -249.735 -83.165 ;
        RECT -250.805 -83.660 -249.735 -83.490 ;
        RECT -246.765 -83.490 -246.595 -83.165 ;
        RECT -246.415 -83.265 -246.045 -82.925 ;
        RECT -245.865 -83.165 -245.315 -82.995 ;
        RECT -241.265 -83.165 -240.715 -82.995 ;
        RECT -245.865 -83.490 -245.695 -83.165 ;
        RECT -246.765 -83.660 -245.695 -83.490 ;
        RECT -240.885 -83.490 -240.715 -83.165 ;
        RECT -240.535 -83.265 -240.165 -82.925 ;
        RECT -239.985 -83.165 -239.055 -82.985 ;
        RECT -237.605 -83.165 -236.675 -82.985 ;
        RECT -239.985 -83.490 -239.815 -83.165 ;
        RECT -240.885 -83.660 -239.815 -83.490 ;
        RECT -236.845 -83.490 -236.675 -83.165 ;
        RECT -236.495 -83.265 -236.125 -82.925 ;
        RECT -235.945 -83.165 -235.395 -82.995 ;
        RECT -231.345 -83.165 -230.795 -82.995 ;
        RECT -235.945 -83.490 -235.775 -83.165 ;
        RECT -236.845 -83.660 -235.775 -83.490 ;
        RECT -230.965 -83.490 -230.795 -83.165 ;
        RECT -230.615 -83.265 -230.245 -82.925 ;
        RECT -230.065 -83.165 -229.135 -82.985 ;
        RECT -227.685 -83.165 -226.755 -82.985 ;
        RECT -230.065 -83.490 -229.895 -83.165 ;
        RECT -230.965 -83.660 -229.895 -83.490 ;
        RECT -226.925 -83.490 -226.755 -83.165 ;
        RECT -226.575 -83.265 -226.205 -82.925 ;
        RECT -226.025 -83.165 -225.475 -82.995 ;
        RECT -221.425 -83.165 -220.875 -82.995 ;
        RECT -226.025 -83.490 -225.855 -83.165 ;
        RECT -226.925 -83.660 -225.855 -83.490 ;
        RECT -221.045 -83.490 -220.875 -83.165 ;
        RECT -220.695 -83.265 -220.325 -82.925 ;
        RECT -220.145 -83.165 -219.215 -82.985 ;
        RECT -217.765 -83.165 -216.835 -82.985 ;
        RECT -220.145 -83.490 -219.975 -83.165 ;
        RECT -221.045 -83.660 -219.975 -83.490 ;
        RECT -217.005 -83.490 -216.835 -83.165 ;
        RECT -216.655 -83.265 -216.285 -82.925 ;
        RECT -216.105 -83.165 -215.555 -82.995 ;
        RECT -211.505 -83.165 -210.955 -82.995 ;
        RECT -216.105 -83.490 -215.935 -83.165 ;
        RECT -217.005 -83.660 -215.935 -83.490 ;
        RECT -211.125 -83.490 -210.955 -83.165 ;
        RECT -210.775 -83.265 -210.405 -82.925 ;
        RECT -210.225 -83.165 -209.295 -82.985 ;
        RECT -207.845 -83.165 -206.915 -82.985 ;
        RECT -210.225 -83.490 -210.055 -83.165 ;
        RECT -211.125 -83.660 -210.055 -83.490 ;
        RECT -207.085 -83.490 -206.915 -83.165 ;
        RECT -206.735 -83.265 -206.365 -82.925 ;
        RECT -206.185 -83.165 -205.635 -82.995 ;
        RECT -201.585 -83.165 -201.035 -82.995 ;
        RECT -206.185 -83.490 -206.015 -83.165 ;
        RECT -207.085 -83.660 -206.015 -83.490 ;
        RECT -201.205 -83.490 -201.035 -83.165 ;
        RECT -200.855 -83.265 -200.485 -82.925 ;
        RECT -200.305 -83.165 -199.375 -82.985 ;
        RECT -197.925 -83.165 -196.995 -82.985 ;
        RECT -200.305 -83.490 -200.135 -83.165 ;
        RECT -201.205 -83.660 -200.135 -83.490 ;
        RECT -197.165 -83.490 -196.995 -83.165 ;
        RECT -196.815 -83.265 -196.445 -82.925 ;
        RECT -196.265 -83.165 -195.715 -82.995 ;
        RECT -191.665 -83.165 -191.115 -82.995 ;
        RECT -196.265 -83.490 -196.095 -83.165 ;
        RECT -197.165 -83.660 -196.095 -83.490 ;
        RECT -191.285 -83.490 -191.115 -83.165 ;
        RECT -190.935 -83.265 -190.565 -82.925 ;
        RECT -190.385 -83.165 -189.455 -82.985 ;
        RECT -188.005 -83.165 -187.075 -82.985 ;
        RECT -190.385 -83.490 -190.215 -83.165 ;
        RECT -191.285 -83.660 -190.215 -83.490 ;
        RECT -187.245 -83.490 -187.075 -83.165 ;
        RECT -186.895 -83.265 -186.525 -82.925 ;
        RECT -186.345 -83.165 -185.795 -82.995 ;
        RECT -181.745 -83.165 -181.195 -82.995 ;
        RECT -186.345 -83.490 -186.175 -83.165 ;
        RECT -187.245 -83.660 -186.175 -83.490 ;
        RECT -181.365 -83.490 -181.195 -83.165 ;
        RECT -181.015 -83.265 -180.645 -82.925 ;
        RECT -180.465 -83.165 -179.535 -82.985 ;
        RECT -178.085 -83.165 -177.155 -82.985 ;
        RECT -180.465 -83.490 -180.295 -83.165 ;
        RECT -181.365 -83.660 -180.295 -83.490 ;
        RECT -177.325 -83.490 -177.155 -83.165 ;
        RECT -176.975 -83.265 -176.605 -82.925 ;
        RECT -176.425 -83.165 -175.875 -82.995 ;
        RECT -171.825 -83.165 -171.275 -82.995 ;
        RECT -176.425 -83.490 -176.255 -83.165 ;
        RECT -177.325 -83.660 -176.255 -83.490 ;
        RECT -171.445 -83.490 -171.275 -83.165 ;
        RECT -171.095 -83.265 -170.725 -82.925 ;
        RECT -170.545 -83.165 -169.615 -82.985 ;
        RECT -168.165 -83.165 -167.235 -82.985 ;
        RECT -170.545 -83.490 -170.375 -83.165 ;
        RECT -171.445 -83.660 -170.375 -83.490 ;
        RECT -167.405 -83.490 -167.235 -83.165 ;
        RECT -167.055 -83.265 -166.685 -82.925 ;
        RECT -166.505 -83.165 -165.955 -82.995 ;
        RECT -161.905 -83.165 -161.355 -82.995 ;
        RECT -166.505 -83.490 -166.335 -83.165 ;
        RECT -167.405 -83.660 -166.335 -83.490 ;
        RECT -161.525 -83.490 -161.355 -83.165 ;
        RECT -161.175 -83.265 -160.805 -82.925 ;
        RECT -160.625 -83.165 -159.695 -82.985 ;
        RECT -158.245 -83.165 -157.315 -82.985 ;
        RECT -160.625 -83.490 -160.455 -83.165 ;
        RECT -161.525 -83.660 -160.455 -83.490 ;
        RECT -157.485 -83.490 -157.315 -83.165 ;
        RECT -157.135 -83.265 -156.765 -82.925 ;
        RECT -156.585 -83.165 -156.035 -82.995 ;
        RECT -151.985 -83.165 -151.435 -82.995 ;
        RECT -156.585 -83.490 -156.415 -83.165 ;
        RECT -157.485 -83.660 -156.415 -83.490 ;
        RECT -151.605 -83.490 -151.435 -83.165 ;
        RECT -151.255 -83.265 -150.885 -82.925 ;
        RECT -150.705 -83.165 -149.775 -82.985 ;
        RECT -148.325 -83.165 -147.395 -82.985 ;
        RECT -150.705 -83.490 -150.535 -83.165 ;
        RECT -151.605 -83.660 -150.535 -83.490 ;
        RECT -147.565 -83.490 -147.395 -83.165 ;
        RECT -147.215 -83.265 -146.845 -82.925 ;
        RECT -146.665 -83.165 -146.115 -82.995 ;
        RECT -142.065 -83.165 -141.515 -82.995 ;
        RECT -146.665 -83.490 -146.495 -83.165 ;
        RECT -147.565 -83.660 -146.495 -83.490 ;
        RECT -141.685 -83.490 -141.515 -83.165 ;
        RECT -141.335 -83.265 -140.965 -82.925 ;
        RECT -140.785 -83.165 -139.855 -82.985 ;
        RECT -138.405 -83.165 -137.475 -82.985 ;
        RECT -140.785 -83.490 -140.615 -83.165 ;
        RECT -141.685 -83.660 -140.615 -83.490 ;
        RECT -137.645 -83.490 -137.475 -83.165 ;
        RECT -137.295 -83.265 -136.925 -82.925 ;
        RECT -136.745 -83.165 -136.195 -82.995 ;
        RECT -132.145 -83.165 -131.595 -82.995 ;
        RECT -136.745 -83.490 -136.575 -83.165 ;
        RECT -137.645 -83.660 -136.575 -83.490 ;
        RECT -131.765 -83.490 -131.595 -83.165 ;
        RECT -131.415 -83.265 -131.045 -82.925 ;
        RECT -130.865 -83.165 -129.935 -82.985 ;
        RECT -128.485 -83.165 -127.555 -82.985 ;
        RECT -130.865 -83.490 -130.695 -83.165 ;
        RECT -131.765 -83.660 -130.695 -83.490 ;
        RECT -127.725 -83.490 -127.555 -83.165 ;
        RECT -127.375 -83.265 -127.005 -82.925 ;
        RECT -126.825 -83.165 -126.275 -82.995 ;
        RECT -122.225 -83.165 -121.675 -82.995 ;
        RECT -126.825 -83.490 -126.655 -83.165 ;
        RECT -127.725 -83.660 -126.655 -83.490 ;
        RECT -121.845 -83.490 -121.675 -83.165 ;
        RECT -121.495 -83.265 -121.125 -82.925 ;
        RECT -120.945 -83.165 -120.015 -82.985 ;
        RECT -118.565 -83.165 -117.635 -82.985 ;
        RECT -120.945 -83.490 -120.775 -83.165 ;
        RECT -121.845 -83.660 -120.775 -83.490 ;
        RECT -117.805 -83.490 -117.635 -83.165 ;
        RECT -117.455 -83.265 -117.085 -82.925 ;
        RECT -116.905 -83.165 -116.355 -82.995 ;
        RECT -112.305 -83.165 -111.755 -82.995 ;
        RECT -116.905 -83.490 -116.735 -83.165 ;
        RECT -117.805 -83.660 -116.735 -83.490 ;
        RECT -111.925 -83.490 -111.755 -83.165 ;
        RECT -111.575 -83.265 -111.205 -82.925 ;
        RECT -111.025 -83.165 -110.095 -82.985 ;
        RECT -108.645 -83.165 -107.715 -82.985 ;
        RECT -111.025 -83.490 -110.855 -83.165 ;
        RECT -111.925 -83.660 -110.855 -83.490 ;
        RECT -107.885 -83.490 -107.715 -83.165 ;
        RECT -107.535 -83.265 -107.165 -82.925 ;
        RECT -106.985 -83.165 -106.435 -82.995 ;
        RECT -102.385 -83.165 -101.835 -82.995 ;
        RECT -106.985 -83.490 -106.815 -83.165 ;
        RECT -107.885 -83.660 -106.815 -83.490 ;
        RECT -102.005 -83.490 -101.835 -83.165 ;
        RECT -101.655 -83.265 -101.285 -82.925 ;
        RECT -101.105 -83.165 -100.175 -82.985 ;
        RECT -98.725 -83.165 -97.795 -82.985 ;
        RECT -101.105 -83.490 -100.935 -83.165 ;
        RECT -102.005 -83.660 -100.935 -83.490 ;
        RECT -97.965 -83.490 -97.795 -83.165 ;
        RECT -97.615 -83.265 -97.245 -82.925 ;
        RECT -97.065 -83.165 -96.515 -82.995 ;
        RECT -92.465 -83.165 -91.915 -82.995 ;
        RECT -97.065 -83.490 -96.895 -83.165 ;
        RECT -97.965 -83.660 -96.895 -83.490 ;
        RECT -92.085 -83.490 -91.915 -83.165 ;
        RECT -91.735 -83.265 -91.365 -82.925 ;
        RECT -91.185 -83.165 -90.255 -82.985 ;
        RECT -88.805 -83.165 -87.875 -82.985 ;
        RECT -91.185 -83.490 -91.015 -83.165 ;
        RECT -92.085 -83.660 -91.015 -83.490 ;
        RECT -88.045 -83.490 -87.875 -83.165 ;
        RECT -87.695 -83.265 -87.325 -82.925 ;
        RECT -87.145 -83.165 -86.595 -82.995 ;
        RECT -82.545 -83.165 -81.995 -82.995 ;
        RECT -87.145 -83.490 -86.975 -83.165 ;
        RECT -88.045 -83.660 -86.975 -83.490 ;
        RECT -82.165 -83.490 -81.995 -83.165 ;
        RECT -81.815 -83.265 -81.445 -82.925 ;
        RECT -81.265 -83.165 -80.335 -82.985 ;
        RECT -78.885 -83.165 -77.955 -82.985 ;
        RECT -81.265 -83.490 -81.095 -83.165 ;
        RECT -82.165 -83.660 -81.095 -83.490 ;
        RECT -78.125 -83.490 -77.955 -83.165 ;
        RECT -77.775 -83.265 -77.405 -82.925 ;
        RECT -77.225 -83.165 -76.675 -82.995 ;
        RECT -72.625 -83.165 -72.075 -82.995 ;
        RECT -77.225 -83.490 -77.055 -83.165 ;
        RECT -78.125 -83.660 -77.055 -83.490 ;
        RECT -72.245 -83.490 -72.075 -83.165 ;
        RECT -71.895 -83.265 -71.525 -82.925 ;
        RECT -71.345 -83.165 -70.415 -82.985 ;
        RECT -68.965 -83.165 -68.035 -82.985 ;
        RECT -71.345 -83.490 -71.175 -83.165 ;
        RECT -72.245 -83.660 -71.175 -83.490 ;
        RECT -68.205 -83.490 -68.035 -83.165 ;
        RECT -67.855 -83.265 -67.485 -82.925 ;
        RECT -67.305 -83.165 -66.755 -82.995 ;
        RECT -62.705 -83.165 -62.155 -82.995 ;
        RECT -67.305 -83.490 -67.135 -83.165 ;
        RECT -68.205 -83.660 -67.135 -83.490 ;
        RECT -62.325 -83.490 -62.155 -83.165 ;
        RECT -61.975 -83.265 -61.605 -82.925 ;
        RECT -61.425 -83.165 -60.495 -82.985 ;
        RECT -59.045 -83.165 -58.115 -82.985 ;
        RECT -61.425 -83.490 -61.255 -83.165 ;
        RECT -62.325 -83.660 -61.255 -83.490 ;
        RECT -58.285 -83.490 -58.115 -83.165 ;
        RECT -57.935 -83.265 -57.565 -82.925 ;
        RECT -57.385 -83.165 -56.835 -82.995 ;
        RECT -52.785 -83.165 -52.235 -82.995 ;
        RECT -57.385 -83.490 -57.215 -83.165 ;
        RECT -58.285 -83.660 -57.215 -83.490 ;
        RECT -52.405 -83.490 -52.235 -83.165 ;
        RECT -52.055 -83.265 -51.685 -82.925 ;
        RECT -51.505 -83.165 -50.575 -82.985 ;
        RECT -49.125 -83.165 -48.195 -82.985 ;
        RECT -51.505 -83.490 -51.335 -83.165 ;
        RECT -52.405 -83.660 -51.335 -83.490 ;
        RECT -48.365 -83.490 -48.195 -83.165 ;
        RECT -48.015 -83.265 -47.645 -82.925 ;
        RECT -47.465 -83.165 -46.915 -82.995 ;
        RECT -42.865 -83.165 -42.315 -82.995 ;
        RECT -47.465 -83.490 -47.295 -83.165 ;
        RECT -48.365 -83.660 -47.295 -83.490 ;
        RECT -42.485 -83.490 -42.315 -83.165 ;
        RECT -42.135 -83.265 -41.765 -82.925 ;
        RECT -41.585 -83.165 -40.655 -82.985 ;
        RECT -39.205 -83.165 -38.275 -82.985 ;
        RECT -41.585 -83.490 -41.415 -83.165 ;
        RECT -42.485 -83.660 -41.415 -83.490 ;
        RECT -38.445 -83.490 -38.275 -83.165 ;
        RECT -38.095 -83.265 -37.725 -82.925 ;
        RECT -37.545 -83.165 -36.995 -82.995 ;
        RECT -32.945 -83.165 -32.395 -82.995 ;
        RECT -37.545 -83.490 -37.375 -83.165 ;
        RECT -38.445 -83.660 -37.375 -83.490 ;
        RECT -32.565 -83.490 -32.395 -83.165 ;
        RECT -32.215 -83.265 -31.845 -82.925 ;
        RECT -31.665 -83.165 -30.735 -82.985 ;
        RECT -29.285 -83.165 -28.355 -82.985 ;
        RECT -31.665 -83.490 -31.495 -83.165 ;
        RECT -32.565 -83.660 -31.495 -83.490 ;
        RECT -28.525 -83.490 -28.355 -83.165 ;
        RECT -28.175 -83.265 -27.805 -82.925 ;
        RECT -27.625 -83.165 -27.075 -82.995 ;
        RECT -23.025 -83.165 -22.475 -82.995 ;
        RECT -27.625 -83.490 -27.455 -83.165 ;
        RECT -28.525 -83.660 -27.455 -83.490 ;
        RECT -22.645 -83.490 -22.475 -83.165 ;
        RECT -22.295 -83.265 -21.925 -82.925 ;
        RECT -21.745 -83.165 -20.815 -82.985 ;
        RECT -19.365 -83.165 -18.435 -82.985 ;
        RECT -21.745 -83.490 -21.575 -83.165 ;
        RECT -22.645 -83.660 -21.575 -83.490 ;
        RECT -18.605 -83.490 -18.435 -83.165 ;
        RECT -18.255 -83.265 -17.885 -82.925 ;
        RECT -17.705 -83.165 -17.155 -82.995 ;
        RECT -13.105 -83.165 -12.555 -82.995 ;
        RECT -17.705 -83.490 -17.535 -83.165 ;
        RECT -18.605 -83.660 -17.535 -83.490 ;
        RECT -12.725 -83.490 -12.555 -83.165 ;
        RECT -12.375 -83.265 -12.005 -82.925 ;
        RECT -11.825 -83.165 -10.895 -82.985 ;
        RECT -9.445 -83.165 -8.515 -82.985 ;
        RECT -11.825 -83.490 -11.655 -83.165 ;
        RECT -12.725 -83.660 -11.655 -83.490 ;
        RECT -8.685 -83.490 -8.515 -83.165 ;
        RECT -8.335 -83.265 -7.965 -82.925 ;
        RECT -7.785 -83.165 -7.235 -82.995 ;
        RECT -3.185 -83.165 -2.635 -82.995 ;
        RECT -7.785 -83.490 -7.615 -83.165 ;
        RECT -8.685 -83.660 -7.615 -83.490 ;
        RECT -2.805 -83.490 -2.635 -83.165 ;
        RECT -2.455 -83.265 -2.085 -82.925 ;
        RECT -1.905 -83.165 -0.975 -82.985 ;
        RECT 0.475 -83.165 1.405 -82.985 ;
        RECT -1.905 -83.490 -1.735 -83.165 ;
        RECT -2.805 -83.660 -1.735 -83.490 ;
        RECT 1.235 -83.490 1.405 -83.165 ;
        RECT 1.585 -83.265 1.955 -82.925 ;
        RECT 2.135 -83.165 2.685 -82.995 ;
        RECT 6.735 -83.165 7.285 -82.995 ;
        RECT 2.135 -83.490 2.305 -83.165 ;
        RECT 1.235 -83.660 2.305 -83.490 ;
        RECT 7.115 -83.490 7.285 -83.165 ;
        RECT 7.465 -83.265 7.835 -82.925 ;
        RECT 8.015 -83.165 8.945 -82.985 ;
        RECT 10.395 -83.165 11.325 -82.985 ;
        RECT 8.015 -83.490 8.185 -83.165 ;
        RECT 7.115 -83.660 8.185 -83.490 ;
        RECT 11.155 -83.490 11.325 -83.165 ;
        RECT 11.505 -83.265 11.875 -82.925 ;
        RECT 12.055 -83.165 12.605 -82.995 ;
        RECT 16.655 -83.165 17.205 -82.995 ;
        RECT 12.055 -83.490 12.225 -83.165 ;
        RECT 11.155 -83.660 12.225 -83.490 ;
        RECT 17.035 -83.490 17.205 -83.165 ;
        RECT 17.385 -83.265 17.755 -82.925 ;
        RECT 17.935 -83.165 18.865 -82.985 ;
        RECT 20.315 -83.165 21.245 -82.985 ;
        RECT 17.935 -83.490 18.105 -83.165 ;
        RECT 17.035 -83.660 18.105 -83.490 ;
        RECT 21.075 -83.490 21.245 -83.165 ;
        RECT 21.425 -83.265 21.795 -82.925 ;
        RECT 21.975 -83.165 22.525 -82.995 ;
        RECT 21.975 -83.490 22.145 -83.165 ;
        RECT 22.695 -83.345 22.865 -82.820 ;
        RECT 21.075 -83.660 22.145 -83.490 ;
        RECT -291.205 -83.860 -291.035 -83.675 ;
        RECT -290.060 -83.765 -289.730 -83.660 ;
        RECT -286.130 -83.765 -285.800 -83.660 ;
        RECT -280.140 -83.765 -279.810 -83.660 ;
        RECT -276.210 -83.765 -275.880 -83.660 ;
        RECT -270.220 -83.765 -269.890 -83.660 ;
        RECT -266.290 -83.765 -265.960 -83.660 ;
        RECT -260.300 -83.765 -259.970 -83.660 ;
        RECT -256.370 -83.765 -256.040 -83.660 ;
        RECT -250.380 -83.765 -250.050 -83.660 ;
        RECT -246.450 -83.765 -246.120 -83.660 ;
        RECT -240.460 -83.765 -240.130 -83.660 ;
        RECT -236.530 -83.765 -236.200 -83.660 ;
        RECT -230.540 -83.765 -230.210 -83.660 ;
        RECT -226.610 -83.765 -226.280 -83.660 ;
        RECT -220.620 -83.765 -220.290 -83.660 ;
        RECT -216.690 -83.765 -216.360 -83.660 ;
        RECT -210.700 -83.765 -210.370 -83.660 ;
        RECT -206.770 -83.765 -206.440 -83.660 ;
        RECT -200.780 -83.765 -200.450 -83.660 ;
        RECT -196.850 -83.765 -196.520 -83.660 ;
        RECT -190.860 -83.765 -190.530 -83.660 ;
        RECT -186.930 -83.765 -186.600 -83.660 ;
        RECT -180.940 -83.765 -180.610 -83.660 ;
        RECT -177.010 -83.765 -176.680 -83.660 ;
        RECT -171.020 -83.765 -170.690 -83.660 ;
        RECT -167.090 -83.765 -166.760 -83.660 ;
        RECT -161.100 -83.765 -160.770 -83.660 ;
        RECT -157.170 -83.765 -156.840 -83.660 ;
        RECT -151.180 -83.765 -150.850 -83.660 ;
        RECT -147.250 -83.765 -146.920 -83.660 ;
        RECT -141.260 -83.765 -140.930 -83.660 ;
        RECT -137.330 -83.765 -137.000 -83.660 ;
        RECT -131.340 -83.765 -131.010 -83.660 ;
        RECT -127.410 -83.765 -127.080 -83.660 ;
        RECT -121.420 -83.765 -121.090 -83.660 ;
        RECT -117.490 -83.765 -117.160 -83.660 ;
        RECT -111.500 -83.765 -111.170 -83.660 ;
        RECT -107.570 -83.765 -107.240 -83.660 ;
        RECT -101.580 -83.765 -101.250 -83.660 ;
        RECT -97.650 -83.765 -97.320 -83.660 ;
        RECT -91.660 -83.765 -91.330 -83.660 ;
        RECT -87.730 -83.765 -87.400 -83.660 ;
        RECT -81.740 -83.765 -81.410 -83.660 ;
        RECT -77.810 -83.765 -77.480 -83.660 ;
        RECT -71.820 -83.765 -71.490 -83.660 ;
        RECT -67.890 -83.765 -67.560 -83.660 ;
        RECT -61.900 -83.765 -61.570 -83.660 ;
        RECT -57.970 -83.765 -57.640 -83.660 ;
        RECT -51.980 -83.765 -51.650 -83.660 ;
        RECT -48.050 -83.765 -47.720 -83.660 ;
        RECT -42.060 -83.765 -41.730 -83.660 ;
        RECT -38.130 -83.765 -37.800 -83.660 ;
        RECT -32.140 -83.765 -31.810 -83.660 ;
        RECT -28.210 -83.765 -27.880 -83.660 ;
        RECT -22.220 -83.765 -21.890 -83.660 ;
        RECT -18.290 -83.765 -17.960 -83.660 ;
        RECT -12.300 -83.765 -11.970 -83.660 ;
        RECT -8.370 -83.765 -8.040 -83.660 ;
        RECT -2.380 -83.765 -2.050 -83.660 ;
        RECT 1.550 -83.765 1.880 -83.660 ;
        RECT 7.540 -83.765 7.870 -83.660 ;
        RECT 11.470 -83.765 11.800 -83.660 ;
        RECT 17.460 -83.765 17.790 -83.660 ;
        RECT 21.390 -83.765 21.720 -83.660 ;
        RECT 22.315 -83.675 22.865 -83.345 ;
        RECT -291.735 -83.875 -291.035 -83.860 ;
        RECT -291.820 -84.045 -291.035 -83.875 ;
        RECT -291.500 -84.050 -291.035 -84.045 ;
        RECT -291.205 -84.200 -291.035 -84.050 ;
        RECT -287.205 -83.935 -286.300 -83.845 ;
        RECT -285.500 -83.935 -284.995 -83.855 ;
        RECT -287.205 -84.115 -284.995 -83.935 ;
        RECT -277.285 -83.935 -276.380 -83.845 ;
        RECT -275.580 -83.935 -275.075 -83.855 ;
        RECT -277.285 -84.115 -275.075 -83.935 ;
        RECT -267.365 -83.935 -266.460 -83.845 ;
        RECT -265.660 -83.935 -265.155 -83.855 ;
        RECT -267.365 -84.115 -265.155 -83.935 ;
        RECT -257.445 -83.935 -256.540 -83.845 ;
        RECT -255.740 -83.935 -255.235 -83.855 ;
        RECT -257.445 -84.115 -255.235 -83.935 ;
        RECT -247.525 -83.935 -246.620 -83.845 ;
        RECT -245.820 -83.935 -245.315 -83.855 ;
        RECT -247.525 -84.115 -245.315 -83.935 ;
        RECT -237.605 -83.935 -236.700 -83.845 ;
        RECT -235.900 -83.935 -235.395 -83.855 ;
        RECT -237.605 -84.115 -235.395 -83.935 ;
        RECT -227.685 -83.935 -226.780 -83.845 ;
        RECT -225.980 -83.935 -225.475 -83.855 ;
        RECT -227.685 -84.115 -225.475 -83.935 ;
        RECT -217.765 -83.935 -216.860 -83.845 ;
        RECT -216.060 -83.935 -215.555 -83.855 ;
        RECT -217.765 -84.115 -215.555 -83.935 ;
        RECT -207.845 -83.935 -206.940 -83.845 ;
        RECT -206.140 -83.935 -205.635 -83.855 ;
        RECT -207.845 -84.115 -205.635 -83.935 ;
        RECT -197.925 -83.935 -197.020 -83.845 ;
        RECT -196.220 -83.935 -195.715 -83.855 ;
        RECT -197.925 -84.115 -195.715 -83.935 ;
        RECT -188.005 -83.935 -187.100 -83.845 ;
        RECT -186.300 -83.935 -185.795 -83.855 ;
        RECT -188.005 -84.115 -185.795 -83.935 ;
        RECT -178.085 -83.935 -177.180 -83.845 ;
        RECT -176.380 -83.935 -175.875 -83.855 ;
        RECT -178.085 -84.115 -175.875 -83.935 ;
        RECT -168.165 -83.935 -167.260 -83.845 ;
        RECT -166.460 -83.935 -165.955 -83.855 ;
        RECT -168.165 -84.115 -165.955 -83.935 ;
        RECT -158.245 -83.935 -157.340 -83.845 ;
        RECT -156.540 -83.935 -156.035 -83.855 ;
        RECT -158.245 -84.115 -156.035 -83.935 ;
        RECT -148.325 -83.935 -147.420 -83.845 ;
        RECT -146.620 -83.935 -146.115 -83.855 ;
        RECT -148.325 -84.115 -146.115 -83.935 ;
        RECT -138.405 -83.935 -137.500 -83.845 ;
        RECT -136.700 -83.935 -136.195 -83.855 ;
        RECT -138.405 -84.115 -136.195 -83.935 ;
        RECT -128.485 -83.935 -127.580 -83.845 ;
        RECT -126.780 -83.935 -126.275 -83.855 ;
        RECT -128.485 -84.115 -126.275 -83.935 ;
        RECT -118.565 -83.935 -117.660 -83.845 ;
        RECT -116.860 -83.935 -116.355 -83.855 ;
        RECT -118.565 -84.115 -116.355 -83.935 ;
        RECT -108.645 -83.935 -107.740 -83.845 ;
        RECT -106.940 -83.935 -106.435 -83.855 ;
        RECT -108.645 -84.115 -106.435 -83.935 ;
        RECT -98.725 -83.935 -97.820 -83.845 ;
        RECT -97.020 -83.935 -96.515 -83.855 ;
        RECT -98.725 -84.115 -96.515 -83.935 ;
        RECT -88.805 -83.935 -87.900 -83.845 ;
        RECT -87.100 -83.935 -86.595 -83.855 ;
        RECT -88.805 -84.115 -86.595 -83.935 ;
        RECT -78.885 -83.935 -77.980 -83.845 ;
        RECT -77.180 -83.935 -76.675 -83.855 ;
        RECT -78.885 -84.115 -76.675 -83.935 ;
        RECT -68.965 -83.935 -68.060 -83.845 ;
        RECT -67.260 -83.935 -66.755 -83.855 ;
        RECT -68.965 -84.115 -66.755 -83.935 ;
        RECT -59.045 -83.935 -58.140 -83.845 ;
        RECT -57.340 -83.935 -56.835 -83.855 ;
        RECT -59.045 -84.115 -56.835 -83.935 ;
        RECT -49.125 -83.935 -48.220 -83.845 ;
        RECT -47.420 -83.935 -46.915 -83.855 ;
        RECT -49.125 -84.115 -46.915 -83.935 ;
        RECT -39.205 -83.935 -38.300 -83.845 ;
        RECT -37.500 -83.935 -36.995 -83.855 ;
        RECT -39.205 -84.115 -36.995 -83.935 ;
        RECT -29.285 -83.935 -28.380 -83.845 ;
        RECT -27.580 -83.935 -27.075 -83.855 ;
        RECT -29.285 -84.115 -27.075 -83.935 ;
        RECT -19.365 -83.935 -18.460 -83.845 ;
        RECT -17.660 -83.935 -17.155 -83.855 ;
        RECT -19.365 -84.115 -17.155 -83.935 ;
        RECT -9.445 -83.935 -8.540 -83.845 ;
        RECT -7.740 -83.935 -7.235 -83.855 ;
        RECT -9.445 -84.115 -7.235 -83.935 ;
        RECT 0.475 -83.935 1.380 -83.845 ;
        RECT 2.180 -83.935 2.685 -83.855 ;
        RECT 0.475 -84.115 2.685 -83.935 ;
        RECT 10.395 -83.935 11.300 -83.845 ;
        RECT 12.100 -83.935 12.605 -83.855 ;
        RECT 10.395 -84.115 12.605 -83.935 ;
        RECT 20.315 -83.935 21.220 -83.845 ;
        RECT 22.020 -83.935 22.525 -83.855 ;
        RECT 20.315 -84.115 22.525 -83.935 ;
        RECT 22.695 -83.870 22.865 -83.675 ;
        RECT 23.105 -83.870 23.395 -83.150 ;
        RECT 22.695 -83.875 23.395 -83.870 ;
        RECT 22.695 -84.045 23.480 -83.875 ;
        RECT 22.695 -84.050 23.160 -84.045 ;
        RECT 22.695 -84.200 22.865 -84.050 ;
        RECT -294.265 -172.590 -294.095 -172.440 ;
        RECT -294.880 -172.760 -294.095 -172.590 ;
        RECT -294.795 -173.925 -294.505 -172.760 ;
        RECT -294.265 -172.965 -294.095 -172.760 ;
        RECT -293.925 -172.705 -291.715 -172.525 ;
        RECT -293.925 -172.795 -293.020 -172.705 ;
        RECT -292.220 -172.785 -291.715 -172.705 ;
        RECT -284.005 -172.705 -281.795 -172.525 ;
        RECT -284.005 -172.795 -283.100 -172.705 ;
        RECT -282.300 -172.785 -281.795 -172.705 ;
        RECT -274.085 -172.705 -271.875 -172.525 ;
        RECT -274.085 -172.795 -273.180 -172.705 ;
        RECT -272.380 -172.785 -271.875 -172.705 ;
        RECT -264.165 -172.705 -261.955 -172.525 ;
        RECT -264.165 -172.795 -263.260 -172.705 ;
        RECT -262.460 -172.785 -261.955 -172.705 ;
        RECT -254.245 -172.705 -252.035 -172.525 ;
        RECT -254.245 -172.795 -253.340 -172.705 ;
        RECT -252.540 -172.785 -252.035 -172.705 ;
        RECT -244.325 -172.705 -242.115 -172.525 ;
        RECT -244.325 -172.795 -243.420 -172.705 ;
        RECT -242.620 -172.785 -242.115 -172.705 ;
        RECT -234.405 -172.705 -232.195 -172.525 ;
        RECT -234.405 -172.795 -233.500 -172.705 ;
        RECT -232.700 -172.785 -232.195 -172.705 ;
        RECT -224.485 -172.705 -222.275 -172.525 ;
        RECT -224.485 -172.795 -223.580 -172.705 ;
        RECT -222.780 -172.785 -222.275 -172.705 ;
        RECT -214.565 -172.705 -212.355 -172.525 ;
        RECT -214.565 -172.795 -213.660 -172.705 ;
        RECT -212.860 -172.785 -212.355 -172.705 ;
        RECT -204.645 -172.705 -202.435 -172.525 ;
        RECT -204.645 -172.795 -203.740 -172.705 ;
        RECT -202.940 -172.785 -202.435 -172.705 ;
        RECT -194.725 -172.705 -192.515 -172.525 ;
        RECT -194.725 -172.795 -193.820 -172.705 ;
        RECT -193.020 -172.785 -192.515 -172.705 ;
        RECT -184.805 -172.705 -182.595 -172.525 ;
        RECT -184.805 -172.795 -183.900 -172.705 ;
        RECT -183.100 -172.785 -182.595 -172.705 ;
        RECT -174.885 -172.705 -172.675 -172.525 ;
        RECT -174.885 -172.795 -173.980 -172.705 ;
        RECT -173.180 -172.785 -172.675 -172.705 ;
        RECT -164.965 -172.705 -162.755 -172.525 ;
        RECT -164.965 -172.795 -164.060 -172.705 ;
        RECT -163.260 -172.785 -162.755 -172.705 ;
        RECT -155.045 -172.705 -152.835 -172.525 ;
        RECT -155.045 -172.795 -154.140 -172.705 ;
        RECT -153.340 -172.785 -152.835 -172.705 ;
        RECT -145.125 -172.705 -142.915 -172.525 ;
        RECT -145.125 -172.795 -144.220 -172.705 ;
        RECT -143.420 -172.785 -142.915 -172.705 ;
        RECT -135.205 -172.705 -132.995 -172.525 ;
        RECT -135.205 -172.795 -134.300 -172.705 ;
        RECT -133.500 -172.785 -132.995 -172.705 ;
        RECT -125.285 -172.705 -123.075 -172.525 ;
        RECT -125.285 -172.795 -124.380 -172.705 ;
        RECT -123.580 -172.785 -123.075 -172.705 ;
        RECT -115.365 -172.705 -113.155 -172.525 ;
        RECT -115.365 -172.795 -114.460 -172.705 ;
        RECT -113.660 -172.785 -113.155 -172.705 ;
        RECT -105.445 -172.705 -103.235 -172.525 ;
        RECT -105.445 -172.795 -104.540 -172.705 ;
        RECT -103.740 -172.785 -103.235 -172.705 ;
        RECT -95.525 -172.705 -93.315 -172.525 ;
        RECT -95.525 -172.795 -94.620 -172.705 ;
        RECT -93.820 -172.785 -93.315 -172.705 ;
        RECT -85.605 -172.705 -83.395 -172.525 ;
        RECT -85.605 -172.795 -84.700 -172.705 ;
        RECT -83.900 -172.785 -83.395 -172.705 ;
        RECT -75.685 -172.705 -73.475 -172.525 ;
        RECT -75.685 -172.795 -74.780 -172.705 ;
        RECT -73.980 -172.785 -73.475 -172.705 ;
        RECT -65.765 -172.705 -63.555 -172.525 ;
        RECT -65.765 -172.795 -64.860 -172.705 ;
        RECT -64.060 -172.785 -63.555 -172.705 ;
        RECT -55.845 -172.705 -53.635 -172.525 ;
        RECT -55.845 -172.795 -54.940 -172.705 ;
        RECT -54.140 -172.785 -53.635 -172.705 ;
        RECT -45.925 -172.705 -43.715 -172.525 ;
        RECT -45.925 -172.795 -45.020 -172.705 ;
        RECT -44.220 -172.785 -43.715 -172.705 ;
        RECT -36.005 -172.705 -33.795 -172.525 ;
        RECT -36.005 -172.795 -35.100 -172.705 ;
        RECT -34.300 -172.785 -33.795 -172.705 ;
        RECT -26.085 -172.705 -23.875 -172.525 ;
        RECT -26.085 -172.795 -25.180 -172.705 ;
        RECT -24.380 -172.785 -23.875 -172.705 ;
        RECT -16.165 -172.705 -13.955 -172.525 ;
        RECT -16.165 -172.795 -15.260 -172.705 ;
        RECT -14.460 -172.785 -13.955 -172.705 ;
        RECT -6.245 -172.705 -4.035 -172.525 ;
        RECT -6.245 -172.795 -5.340 -172.705 ;
        RECT -4.540 -172.785 -4.035 -172.705 ;
        RECT 3.675 -172.705 5.885 -172.525 ;
        RECT 3.675 -172.795 4.580 -172.705 ;
        RECT 5.380 -172.785 5.885 -172.705 ;
        RECT 13.595 -172.705 15.805 -172.525 ;
        RECT 13.595 -172.795 14.500 -172.705 ;
        RECT 15.300 -172.785 15.805 -172.705 ;
        RECT -294.265 -173.295 -293.335 -172.965 ;
        RECT -292.850 -172.980 -292.520 -172.875 ;
        RECT -286.860 -172.980 -286.530 -172.875 ;
        RECT -282.930 -172.980 -282.600 -172.875 ;
        RECT -276.940 -172.980 -276.610 -172.875 ;
        RECT -273.010 -172.980 -272.680 -172.875 ;
        RECT -267.020 -172.980 -266.690 -172.875 ;
        RECT -263.090 -172.980 -262.760 -172.875 ;
        RECT -257.100 -172.980 -256.770 -172.875 ;
        RECT -253.170 -172.980 -252.840 -172.875 ;
        RECT -247.180 -172.980 -246.850 -172.875 ;
        RECT -243.250 -172.980 -242.920 -172.875 ;
        RECT -237.260 -172.980 -236.930 -172.875 ;
        RECT -233.330 -172.980 -233.000 -172.875 ;
        RECT -227.340 -172.980 -227.010 -172.875 ;
        RECT -223.410 -172.980 -223.080 -172.875 ;
        RECT -217.420 -172.980 -217.090 -172.875 ;
        RECT -213.490 -172.980 -213.160 -172.875 ;
        RECT -207.500 -172.980 -207.170 -172.875 ;
        RECT -203.570 -172.980 -203.240 -172.875 ;
        RECT -197.580 -172.980 -197.250 -172.875 ;
        RECT -193.650 -172.980 -193.320 -172.875 ;
        RECT -187.660 -172.980 -187.330 -172.875 ;
        RECT -183.730 -172.980 -183.400 -172.875 ;
        RECT -177.740 -172.980 -177.410 -172.875 ;
        RECT -173.810 -172.980 -173.480 -172.875 ;
        RECT -167.820 -172.980 -167.490 -172.875 ;
        RECT -163.890 -172.980 -163.560 -172.875 ;
        RECT -157.900 -172.980 -157.570 -172.875 ;
        RECT -153.970 -172.980 -153.640 -172.875 ;
        RECT -147.980 -172.980 -147.650 -172.875 ;
        RECT -144.050 -172.980 -143.720 -172.875 ;
        RECT -138.060 -172.980 -137.730 -172.875 ;
        RECT -134.130 -172.980 -133.800 -172.875 ;
        RECT -128.140 -172.980 -127.810 -172.875 ;
        RECT -124.210 -172.980 -123.880 -172.875 ;
        RECT -118.220 -172.980 -117.890 -172.875 ;
        RECT -114.290 -172.980 -113.960 -172.875 ;
        RECT -108.300 -172.980 -107.970 -172.875 ;
        RECT -104.370 -172.980 -104.040 -172.875 ;
        RECT -98.380 -172.980 -98.050 -172.875 ;
        RECT -94.450 -172.980 -94.120 -172.875 ;
        RECT -88.460 -172.980 -88.130 -172.875 ;
        RECT -84.530 -172.980 -84.200 -172.875 ;
        RECT -78.540 -172.980 -78.210 -172.875 ;
        RECT -74.610 -172.980 -74.280 -172.875 ;
        RECT -68.620 -172.980 -68.290 -172.875 ;
        RECT -64.690 -172.980 -64.360 -172.875 ;
        RECT -58.700 -172.980 -58.370 -172.875 ;
        RECT -54.770 -172.980 -54.440 -172.875 ;
        RECT -48.780 -172.980 -48.450 -172.875 ;
        RECT -44.850 -172.980 -44.520 -172.875 ;
        RECT -38.860 -172.980 -38.530 -172.875 ;
        RECT -34.930 -172.980 -34.600 -172.875 ;
        RECT -28.940 -172.980 -28.610 -172.875 ;
        RECT -25.010 -172.980 -24.680 -172.875 ;
        RECT -19.020 -172.980 -18.690 -172.875 ;
        RECT -15.090 -172.980 -14.760 -172.875 ;
        RECT -9.100 -172.980 -8.770 -172.875 ;
        RECT -5.170 -172.980 -4.840 -172.875 ;
        RECT 0.820 -172.980 1.150 -172.875 ;
        RECT 4.750 -172.980 5.080 -172.875 ;
        RECT 10.740 -172.980 11.070 -172.875 ;
        RECT 14.670 -172.980 15.000 -172.875 ;
        RECT 20.660 -172.980 20.990 -172.875 ;
        RECT -293.165 -173.150 -292.095 -172.980 ;
        RECT -294.265 -173.820 -294.095 -173.295 ;
        RECT -293.165 -173.475 -292.995 -173.150 ;
        RECT -293.925 -173.655 -292.995 -173.475 ;
        RECT -292.815 -173.715 -292.445 -173.375 ;
        RECT -292.265 -173.475 -292.095 -173.150 ;
        RECT -287.285 -173.150 -286.215 -172.980 ;
        RECT -287.285 -173.475 -287.115 -173.150 ;
        RECT -292.265 -173.645 -291.715 -173.475 ;
        RECT -287.665 -173.645 -287.115 -173.475 ;
        RECT -286.935 -173.715 -286.565 -173.375 ;
        RECT -286.385 -173.475 -286.215 -173.150 ;
        RECT -283.245 -173.150 -282.175 -172.980 ;
        RECT -283.245 -173.475 -283.075 -173.150 ;
        RECT -286.385 -173.655 -285.455 -173.475 ;
        RECT -284.005 -173.655 -283.075 -173.475 ;
        RECT -282.895 -173.715 -282.525 -173.375 ;
        RECT -282.345 -173.475 -282.175 -173.150 ;
        RECT -277.365 -173.150 -276.295 -172.980 ;
        RECT -277.365 -173.475 -277.195 -173.150 ;
        RECT -282.345 -173.645 -281.795 -173.475 ;
        RECT -277.745 -173.645 -277.195 -173.475 ;
        RECT -277.015 -173.715 -276.645 -173.375 ;
        RECT -276.465 -173.475 -276.295 -173.150 ;
        RECT -273.325 -173.150 -272.255 -172.980 ;
        RECT -273.325 -173.475 -273.155 -173.150 ;
        RECT -276.465 -173.655 -275.535 -173.475 ;
        RECT -274.085 -173.655 -273.155 -173.475 ;
        RECT -272.975 -173.715 -272.605 -173.375 ;
        RECT -272.425 -173.475 -272.255 -173.150 ;
        RECT -267.445 -173.150 -266.375 -172.980 ;
        RECT -267.445 -173.475 -267.275 -173.150 ;
        RECT -272.425 -173.645 -271.875 -173.475 ;
        RECT -267.825 -173.645 -267.275 -173.475 ;
        RECT -267.095 -173.715 -266.725 -173.375 ;
        RECT -266.545 -173.475 -266.375 -173.150 ;
        RECT -263.405 -173.150 -262.335 -172.980 ;
        RECT -263.405 -173.475 -263.235 -173.150 ;
        RECT -266.545 -173.655 -265.615 -173.475 ;
        RECT -264.165 -173.655 -263.235 -173.475 ;
        RECT -263.055 -173.715 -262.685 -173.375 ;
        RECT -262.505 -173.475 -262.335 -173.150 ;
        RECT -257.525 -173.150 -256.455 -172.980 ;
        RECT -257.525 -173.475 -257.355 -173.150 ;
        RECT -262.505 -173.645 -261.955 -173.475 ;
        RECT -257.905 -173.645 -257.355 -173.475 ;
        RECT -257.175 -173.715 -256.805 -173.375 ;
        RECT -256.625 -173.475 -256.455 -173.150 ;
        RECT -253.485 -173.150 -252.415 -172.980 ;
        RECT -253.485 -173.475 -253.315 -173.150 ;
        RECT -256.625 -173.655 -255.695 -173.475 ;
        RECT -254.245 -173.655 -253.315 -173.475 ;
        RECT -253.135 -173.715 -252.765 -173.375 ;
        RECT -252.585 -173.475 -252.415 -173.150 ;
        RECT -247.605 -173.150 -246.535 -172.980 ;
        RECT -247.605 -173.475 -247.435 -173.150 ;
        RECT -252.585 -173.645 -252.035 -173.475 ;
        RECT -247.985 -173.645 -247.435 -173.475 ;
        RECT -247.255 -173.715 -246.885 -173.375 ;
        RECT -246.705 -173.475 -246.535 -173.150 ;
        RECT -243.565 -173.150 -242.495 -172.980 ;
        RECT -243.565 -173.475 -243.395 -173.150 ;
        RECT -246.705 -173.655 -245.775 -173.475 ;
        RECT -244.325 -173.655 -243.395 -173.475 ;
        RECT -243.215 -173.715 -242.845 -173.375 ;
        RECT -242.665 -173.475 -242.495 -173.150 ;
        RECT -237.685 -173.150 -236.615 -172.980 ;
        RECT -237.685 -173.475 -237.515 -173.150 ;
        RECT -242.665 -173.645 -242.115 -173.475 ;
        RECT -238.065 -173.645 -237.515 -173.475 ;
        RECT -237.335 -173.715 -236.965 -173.375 ;
        RECT -236.785 -173.475 -236.615 -173.150 ;
        RECT -233.645 -173.150 -232.575 -172.980 ;
        RECT -233.645 -173.475 -233.475 -173.150 ;
        RECT -236.785 -173.655 -235.855 -173.475 ;
        RECT -234.405 -173.655 -233.475 -173.475 ;
        RECT -233.295 -173.715 -232.925 -173.375 ;
        RECT -232.745 -173.475 -232.575 -173.150 ;
        RECT -227.765 -173.150 -226.695 -172.980 ;
        RECT -227.765 -173.475 -227.595 -173.150 ;
        RECT -232.745 -173.645 -232.195 -173.475 ;
        RECT -228.145 -173.645 -227.595 -173.475 ;
        RECT -227.415 -173.715 -227.045 -173.375 ;
        RECT -226.865 -173.475 -226.695 -173.150 ;
        RECT -223.725 -173.150 -222.655 -172.980 ;
        RECT -223.725 -173.475 -223.555 -173.150 ;
        RECT -226.865 -173.655 -225.935 -173.475 ;
        RECT -224.485 -173.655 -223.555 -173.475 ;
        RECT -223.375 -173.715 -223.005 -173.375 ;
        RECT -222.825 -173.475 -222.655 -173.150 ;
        RECT -217.845 -173.150 -216.775 -172.980 ;
        RECT -217.845 -173.475 -217.675 -173.150 ;
        RECT -222.825 -173.645 -222.275 -173.475 ;
        RECT -218.225 -173.645 -217.675 -173.475 ;
        RECT -217.495 -173.715 -217.125 -173.375 ;
        RECT -216.945 -173.475 -216.775 -173.150 ;
        RECT -213.805 -173.150 -212.735 -172.980 ;
        RECT -213.805 -173.475 -213.635 -173.150 ;
        RECT -216.945 -173.655 -216.015 -173.475 ;
        RECT -214.565 -173.655 -213.635 -173.475 ;
        RECT -213.455 -173.715 -213.085 -173.375 ;
        RECT -212.905 -173.475 -212.735 -173.150 ;
        RECT -207.925 -173.150 -206.855 -172.980 ;
        RECT -207.925 -173.475 -207.755 -173.150 ;
        RECT -212.905 -173.645 -212.355 -173.475 ;
        RECT -208.305 -173.645 -207.755 -173.475 ;
        RECT -207.575 -173.715 -207.205 -173.375 ;
        RECT -207.025 -173.475 -206.855 -173.150 ;
        RECT -203.885 -173.150 -202.815 -172.980 ;
        RECT -203.885 -173.475 -203.715 -173.150 ;
        RECT -207.025 -173.655 -206.095 -173.475 ;
        RECT -204.645 -173.655 -203.715 -173.475 ;
        RECT -203.535 -173.715 -203.165 -173.375 ;
        RECT -202.985 -173.475 -202.815 -173.150 ;
        RECT -198.005 -173.150 -196.935 -172.980 ;
        RECT -198.005 -173.475 -197.835 -173.150 ;
        RECT -202.985 -173.645 -202.435 -173.475 ;
        RECT -198.385 -173.645 -197.835 -173.475 ;
        RECT -197.655 -173.715 -197.285 -173.375 ;
        RECT -197.105 -173.475 -196.935 -173.150 ;
        RECT -193.965 -173.150 -192.895 -172.980 ;
        RECT -193.965 -173.475 -193.795 -173.150 ;
        RECT -197.105 -173.655 -196.175 -173.475 ;
        RECT -194.725 -173.655 -193.795 -173.475 ;
        RECT -193.615 -173.715 -193.245 -173.375 ;
        RECT -193.065 -173.475 -192.895 -173.150 ;
        RECT -188.085 -173.150 -187.015 -172.980 ;
        RECT -188.085 -173.475 -187.915 -173.150 ;
        RECT -193.065 -173.645 -192.515 -173.475 ;
        RECT -188.465 -173.645 -187.915 -173.475 ;
        RECT -187.735 -173.715 -187.365 -173.375 ;
        RECT -187.185 -173.475 -187.015 -173.150 ;
        RECT -184.045 -173.150 -182.975 -172.980 ;
        RECT -184.045 -173.475 -183.875 -173.150 ;
        RECT -187.185 -173.655 -186.255 -173.475 ;
        RECT -184.805 -173.655 -183.875 -173.475 ;
        RECT -183.695 -173.715 -183.325 -173.375 ;
        RECT -183.145 -173.475 -182.975 -173.150 ;
        RECT -178.165 -173.150 -177.095 -172.980 ;
        RECT -178.165 -173.475 -177.995 -173.150 ;
        RECT -183.145 -173.645 -182.595 -173.475 ;
        RECT -178.545 -173.645 -177.995 -173.475 ;
        RECT -177.815 -173.715 -177.445 -173.375 ;
        RECT -177.265 -173.475 -177.095 -173.150 ;
        RECT -174.125 -173.150 -173.055 -172.980 ;
        RECT -174.125 -173.475 -173.955 -173.150 ;
        RECT -177.265 -173.655 -176.335 -173.475 ;
        RECT -174.885 -173.655 -173.955 -173.475 ;
        RECT -173.775 -173.715 -173.405 -173.375 ;
        RECT -173.225 -173.475 -173.055 -173.150 ;
        RECT -168.245 -173.150 -167.175 -172.980 ;
        RECT -168.245 -173.475 -168.075 -173.150 ;
        RECT -173.225 -173.645 -172.675 -173.475 ;
        RECT -168.625 -173.645 -168.075 -173.475 ;
        RECT -167.895 -173.715 -167.525 -173.375 ;
        RECT -167.345 -173.475 -167.175 -173.150 ;
        RECT -164.205 -173.150 -163.135 -172.980 ;
        RECT -164.205 -173.475 -164.035 -173.150 ;
        RECT -167.345 -173.655 -166.415 -173.475 ;
        RECT -164.965 -173.655 -164.035 -173.475 ;
        RECT -163.855 -173.715 -163.485 -173.375 ;
        RECT -163.305 -173.475 -163.135 -173.150 ;
        RECT -158.325 -173.150 -157.255 -172.980 ;
        RECT -158.325 -173.475 -158.155 -173.150 ;
        RECT -163.305 -173.645 -162.755 -173.475 ;
        RECT -158.705 -173.645 -158.155 -173.475 ;
        RECT -157.975 -173.715 -157.605 -173.375 ;
        RECT -157.425 -173.475 -157.255 -173.150 ;
        RECT -154.285 -173.150 -153.215 -172.980 ;
        RECT -154.285 -173.475 -154.115 -173.150 ;
        RECT -157.425 -173.655 -156.495 -173.475 ;
        RECT -155.045 -173.655 -154.115 -173.475 ;
        RECT -153.935 -173.715 -153.565 -173.375 ;
        RECT -153.385 -173.475 -153.215 -173.150 ;
        RECT -148.405 -173.150 -147.335 -172.980 ;
        RECT -148.405 -173.475 -148.235 -173.150 ;
        RECT -153.385 -173.645 -152.835 -173.475 ;
        RECT -148.785 -173.645 -148.235 -173.475 ;
        RECT -148.055 -173.715 -147.685 -173.375 ;
        RECT -147.505 -173.475 -147.335 -173.150 ;
        RECT -144.365 -173.150 -143.295 -172.980 ;
        RECT -144.365 -173.475 -144.195 -173.150 ;
        RECT -147.505 -173.655 -146.575 -173.475 ;
        RECT -145.125 -173.655 -144.195 -173.475 ;
        RECT -144.015 -173.715 -143.645 -173.375 ;
        RECT -143.465 -173.475 -143.295 -173.150 ;
        RECT -138.485 -173.150 -137.415 -172.980 ;
        RECT -138.485 -173.475 -138.315 -173.150 ;
        RECT -143.465 -173.645 -142.915 -173.475 ;
        RECT -138.865 -173.645 -138.315 -173.475 ;
        RECT -138.135 -173.715 -137.765 -173.375 ;
        RECT -137.585 -173.475 -137.415 -173.150 ;
        RECT -134.445 -173.150 -133.375 -172.980 ;
        RECT -134.445 -173.475 -134.275 -173.150 ;
        RECT -137.585 -173.655 -136.655 -173.475 ;
        RECT -135.205 -173.655 -134.275 -173.475 ;
        RECT -134.095 -173.715 -133.725 -173.375 ;
        RECT -133.545 -173.475 -133.375 -173.150 ;
        RECT -128.565 -173.150 -127.495 -172.980 ;
        RECT -128.565 -173.475 -128.395 -173.150 ;
        RECT -133.545 -173.645 -132.995 -173.475 ;
        RECT -128.945 -173.645 -128.395 -173.475 ;
        RECT -128.215 -173.715 -127.845 -173.375 ;
        RECT -127.665 -173.475 -127.495 -173.150 ;
        RECT -124.525 -173.150 -123.455 -172.980 ;
        RECT -124.525 -173.475 -124.355 -173.150 ;
        RECT -127.665 -173.655 -126.735 -173.475 ;
        RECT -125.285 -173.655 -124.355 -173.475 ;
        RECT -124.175 -173.715 -123.805 -173.375 ;
        RECT -123.625 -173.475 -123.455 -173.150 ;
        RECT -118.645 -173.150 -117.575 -172.980 ;
        RECT -118.645 -173.475 -118.475 -173.150 ;
        RECT -123.625 -173.645 -123.075 -173.475 ;
        RECT -119.025 -173.645 -118.475 -173.475 ;
        RECT -118.295 -173.715 -117.925 -173.375 ;
        RECT -117.745 -173.475 -117.575 -173.150 ;
        RECT -114.605 -173.150 -113.535 -172.980 ;
        RECT -114.605 -173.475 -114.435 -173.150 ;
        RECT -117.745 -173.655 -116.815 -173.475 ;
        RECT -115.365 -173.655 -114.435 -173.475 ;
        RECT -114.255 -173.715 -113.885 -173.375 ;
        RECT -113.705 -173.475 -113.535 -173.150 ;
        RECT -108.725 -173.150 -107.655 -172.980 ;
        RECT -108.725 -173.475 -108.555 -173.150 ;
        RECT -113.705 -173.645 -113.155 -173.475 ;
        RECT -109.105 -173.645 -108.555 -173.475 ;
        RECT -108.375 -173.715 -108.005 -173.375 ;
        RECT -107.825 -173.475 -107.655 -173.150 ;
        RECT -104.685 -173.150 -103.615 -172.980 ;
        RECT -104.685 -173.475 -104.515 -173.150 ;
        RECT -107.825 -173.655 -106.895 -173.475 ;
        RECT -105.445 -173.655 -104.515 -173.475 ;
        RECT -104.335 -173.715 -103.965 -173.375 ;
        RECT -103.785 -173.475 -103.615 -173.150 ;
        RECT -98.805 -173.150 -97.735 -172.980 ;
        RECT -98.805 -173.475 -98.635 -173.150 ;
        RECT -103.785 -173.645 -103.235 -173.475 ;
        RECT -99.185 -173.645 -98.635 -173.475 ;
        RECT -98.455 -173.715 -98.085 -173.375 ;
        RECT -97.905 -173.475 -97.735 -173.150 ;
        RECT -94.765 -173.150 -93.695 -172.980 ;
        RECT -94.765 -173.475 -94.595 -173.150 ;
        RECT -97.905 -173.655 -96.975 -173.475 ;
        RECT -95.525 -173.655 -94.595 -173.475 ;
        RECT -94.415 -173.715 -94.045 -173.375 ;
        RECT -93.865 -173.475 -93.695 -173.150 ;
        RECT -88.885 -173.150 -87.815 -172.980 ;
        RECT -88.885 -173.475 -88.715 -173.150 ;
        RECT -93.865 -173.645 -93.315 -173.475 ;
        RECT -89.265 -173.645 -88.715 -173.475 ;
        RECT -88.535 -173.715 -88.165 -173.375 ;
        RECT -87.985 -173.475 -87.815 -173.150 ;
        RECT -84.845 -173.150 -83.775 -172.980 ;
        RECT -84.845 -173.475 -84.675 -173.150 ;
        RECT -87.985 -173.655 -87.055 -173.475 ;
        RECT -85.605 -173.655 -84.675 -173.475 ;
        RECT -84.495 -173.715 -84.125 -173.375 ;
        RECT -83.945 -173.475 -83.775 -173.150 ;
        RECT -78.965 -173.150 -77.895 -172.980 ;
        RECT -78.965 -173.475 -78.795 -173.150 ;
        RECT -83.945 -173.645 -83.395 -173.475 ;
        RECT -79.345 -173.645 -78.795 -173.475 ;
        RECT -78.615 -173.715 -78.245 -173.375 ;
        RECT -78.065 -173.475 -77.895 -173.150 ;
        RECT -74.925 -173.150 -73.855 -172.980 ;
        RECT -74.925 -173.475 -74.755 -173.150 ;
        RECT -78.065 -173.655 -77.135 -173.475 ;
        RECT -75.685 -173.655 -74.755 -173.475 ;
        RECT -74.575 -173.715 -74.205 -173.375 ;
        RECT -74.025 -173.475 -73.855 -173.150 ;
        RECT -69.045 -173.150 -67.975 -172.980 ;
        RECT -69.045 -173.475 -68.875 -173.150 ;
        RECT -74.025 -173.645 -73.475 -173.475 ;
        RECT -69.425 -173.645 -68.875 -173.475 ;
        RECT -68.695 -173.715 -68.325 -173.375 ;
        RECT -68.145 -173.475 -67.975 -173.150 ;
        RECT -65.005 -173.150 -63.935 -172.980 ;
        RECT -65.005 -173.475 -64.835 -173.150 ;
        RECT -68.145 -173.655 -67.215 -173.475 ;
        RECT -65.765 -173.655 -64.835 -173.475 ;
        RECT -64.655 -173.715 -64.285 -173.375 ;
        RECT -64.105 -173.475 -63.935 -173.150 ;
        RECT -59.125 -173.150 -58.055 -172.980 ;
        RECT -59.125 -173.475 -58.955 -173.150 ;
        RECT -64.105 -173.645 -63.555 -173.475 ;
        RECT -59.505 -173.645 -58.955 -173.475 ;
        RECT -58.775 -173.715 -58.405 -173.375 ;
        RECT -58.225 -173.475 -58.055 -173.150 ;
        RECT -55.085 -173.150 -54.015 -172.980 ;
        RECT -55.085 -173.475 -54.915 -173.150 ;
        RECT -58.225 -173.655 -57.295 -173.475 ;
        RECT -55.845 -173.655 -54.915 -173.475 ;
        RECT -54.735 -173.715 -54.365 -173.375 ;
        RECT -54.185 -173.475 -54.015 -173.150 ;
        RECT -49.205 -173.150 -48.135 -172.980 ;
        RECT -49.205 -173.475 -49.035 -173.150 ;
        RECT -54.185 -173.645 -53.635 -173.475 ;
        RECT -49.585 -173.645 -49.035 -173.475 ;
        RECT -48.855 -173.715 -48.485 -173.375 ;
        RECT -48.305 -173.475 -48.135 -173.150 ;
        RECT -45.165 -173.150 -44.095 -172.980 ;
        RECT -45.165 -173.475 -44.995 -173.150 ;
        RECT -48.305 -173.655 -47.375 -173.475 ;
        RECT -45.925 -173.655 -44.995 -173.475 ;
        RECT -44.815 -173.715 -44.445 -173.375 ;
        RECT -44.265 -173.475 -44.095 -173.150 ;
        RECT -39.285 -173.150 -38.215 -172.980 ;
        RECT -39.285 -173.475 -39.115 -173.150 ;
        RECT -44.265 -173.645 -43.715 -173.475 ;
        RECT -39.665 -173.645 -39.115 -173.475 ;
        RECT -38.935 -173.715 -38.565 -173.375 ;
        RECT -38.385 -173.475 -38.215 -173.150 ;
        RECT -35.245 -173.150 -34.175 -172.980 ;
        RECT -35.245 -173.475 -35.075 -173.150 ;
        RECT -38.385 -173.655 -37.455 -173.475 ;
        RECT -36.005 -173.655 -35.075 -173.475 ;
        RECT -34.895 -173.715 -34.525 -173.375 ;
        RECT -34.345 -173.475 -34.175 -173.150 ;
        RECT -29.365 -173.150 -28.295 -172.980 ;
        RECT -29.365 -173.475 -29.195 -173.150 ;
        RECT -34.345 -173.645 -33.795 -173.475 ;
        RECT -29.745 -173.645 -29.195 -173.475 ;
        RECT -29.015 -173.715 -28.645 -173.375 ;
        RECT -28.465 -173.475 -28.295 -173.150 ;
        RECT -25.325 -173.150 -24.255 -172.980 ;
        RECT -25.325 -173.475 -25.155 -173.150 ;
        RECT -28.465 -173.655 -27.535 -173.475 ;
        RECT -26.085 -173.655 -25.155 -173.475 ;
        RECT -24.975 -173.715 -24.605 -173.375 ;
        RECT -24.425 -173.475 -24.255 -173.150 ;
        RECT -19.445 -173.150 -18.375 -172.980 ;
        RECT -19.445 -173.475 -19.275 -173.150 ;
        RECT -24.425 -173.645 -23.875 -173.475 ;
        RECT -19.825 -173.645 -19.275 -173.475 ;
        RECT -19.095 -173.715 -18.725 -173.375 ;
        RECT -18.545 -173.475 -18.375 -173.150 ;
        RECT -15.405 -173.150 -14.335 -172.980 ;
        RECT -15.405 -173.475 -15.235 -173.150 ;
        RECT -18.545 -173.655 -17.615 -173.475 ;
        RECT -16.165 -173.655 -15.235 -173.475 ;
        RECT -15.055 -173.715 -14.685 -173.375 ;
        RECT -14.505 -173.475 -14.335 -173.150 ;
        RECT -9.525 -173.150 -8.455 -172.980 ;
        RECT -9.525 -173.475 -9.355 -173.150 ;
        RECT -14.505 -173.645 -13.955 -173.475 ;
        RECT -9.905 -173.645 -9.355 -173.475 ;
        RECT -9.175 -173.715 -8.805 -173.375 ;
        RECT -8.625 -173.475 -8.455 -173.150 ;
        RECT -5.485 -173.150 -4.415 -172.980 ;
        RECT -5.485 -173.475 -5.315 -173.150 ;
        RECT -8.625 -173.655 -7.695 -173.475 ;
        RECT -6.245 -173.655 -5.315 -173.475 ;
        RECT -5.135 -173.715 -4.765 -173.375 ;
        RECT -4.585 -173.475 -4.415 -173.150 ;
        RECT 0.395 -173.150 1.465 -172.980 ;
        RECT 0.395 -173.475 0.565 -173.150 ;
        RECT -4.585 -173.645 -4.035 -173.475 ;
        RECT 0.015 -173.645 0.565 -173.475 ;
        RECT 0.745 -173.715 1.115 -173.375 ;
        RECT 1.295 -173.475 1.465 -173.150 ;
        RECT 4.435 -173.150 5.505 -172.980 ;
        RECT 4.435 -173.475 4.605 -173.150 ;
        RECT 1.295 -173.655 2.225 -173.475 ;
        RECT 3.675 -173.655 4.605 -173.475 ;
        RECT 4.785 -173.715 5.155 -173.375 ;
        RECT 5.335 -173.475 5.505 -173.150 ;
        RECT 10.315 -173.150 11.385 -172.980 ;
        RECT 10.315 -173.475 10.485 -173.150 ;
        RECT 5.335 -173.645 5.885 -173.475 ;
        RECT 9.935 -173.645 10.485 -173.475 ;
        RECT 10.665 -173.715 11.035 -173.375 ;
        RECT 11.215 -173.475 11.385 -173.150 ;
        RECT 14.355 -173.150 15.425 -172.980 ;
        RECT 14.355 -173.475 14.525 -173.150 ;
        RECT 11.215 -173.655 12.145 -173.475 ;
        RECT 13.595 -173.655 14.525 -173.475 ;
        RECT 14.705 -173.715 15.075 -173.375 ;
        RECT 15.255 -173.475 15.425 -173.150 ;
        RECT 20.235 -173.150 21.305 -172.980 ;
        RECT 20.235 -173.475 20.405 -173.150 ;
        RECT 15.255 -173.645 15.805 -173.475 ;
        RECT 19.855 -173.645 20.405 -173.475 ;
        RECT 20.585 -173.715 20.955 -173.375 ;
        RECT 21.135 -173.475 21.305 -173.150 ;
        RECT 21.135 -173.655 22.065 -173.475 ;
        RECT -294.880 -174.335 -293.040 -174.165 ;
        RECT 21.180 -174.335 23.020 -174.165 ;
        RECT -294.795 -175.060 -294.505 -174.335 ;
        RECT -294.335 -175.135 -294.025 -174.335 ;
        RECT -293.820 -175.135 -293.125 -174.505 ;
        RECT -294.795 -176.885 -294.505 -175.720 ;
        RECT -293.820 -175.735 -293.650 -175.135 ;
        RECT -293.480 -175.575 -293.145 -175.325 ;
        RECT -290.785 -175.485 -290.455 -174.505 ;
        RECT -288.925 -175.485 -288.595 -174.505 ;
        RECT -286.255 -175.135 -285.560 -174.505 ;
        RECT -294.335 -176.885 -294.055 -175.745 ;
        RECT -293.885 -176.715 -293.555 -175.735 ;
        RECT -293.385 -176.885 -293.125 -175.745 ;
        RECT -291.195 -175.895 -290.860 -175.645 ;
        RECT -290.690 -176.085 -290.520 -175.485 ;
        RECT -291.215 -176.715 -290.520 -176.085 ;
        RECT -288.860 -176.085 -288.690 -175.485 ;
        RECT -286.235 -175.575 -285.900 -175.325 ;
        RECT -288.520 -175.895 -288.185 -175.645 ;
        RECT -285.730 -175.735 -285.560 -175.135 ;
        RECT -283.900 -175.135 -283.205 -174.505 ;
        RECT -283.900 -175.735 -283.730 -175.135 ;
        RECT -283.560 -175.575 -283.225 -175.325 ;
        RECT -280.865 -175.485 -280.535 -174.505 ;
        RECT -279.005 -175.485 -278.675 -174.505 ;
        RECT -276.335 -175.135 -275.640 -174.505 ;
        RECT -288.860 -176.715 -288.165 -176.085 ;
        RECT -285.825 -176.715 -285.495 -175.735 ;
        RECT -283.965 -176.715 -283.635 -175.735 ;
        RECT -281.275 -175.895 -280.940 -175.645 ;
        RECT -280.770 -176.085 -280.600 -175.485 ;
        RECT -281.295 -176.715 -280.600 -176.085 ;
        RECT -278.940 -176.085 -278.770 -175.485 ;
        RECT -276.315 -175.575 -275.980 -175.325 ;
        RECT -278.600 -175.895 -278.265 -175.645 ;
        RECT -275.810 -175.735 -275.640 -175.135 ;
        RECT -273.980 -175.135 -273.285 -174.505 ;
        RECT -273.980 -175.735 -273.810 -175.135 ;
        RECT -273.640 -175.575 -273.305 -175.325 ;
        RECT -270.945 -175.485 -270.615 -174.505 ;
        RECT -269.085 -175.485 -268.755 -174.505 ;
        RECT -266.415 -175.135 -265.720 -174.505 ;
        RECT -278.940 -176.715 -278.245 -176.085 ;
        RECT -275.905 -176.715 -275.575 -175.735 ;
        RECT -274.045 -176.715 -273.715 -175.735 ;
        RECT -271.355 -175.895 -271.020 -175.645 ;
        RECT -270.850 -176.085 -270.680 -175.485 ;
        RECT -271.375 -176.715 -270.680 -176.085 ;
        RECT -269.020 -176.085 -268.850 -175.485 ;
        RECT -266.395 -175.575 -266.060 -175.325 ;
        RECT -268.680 -175.895 -268.345 -175.645 ;
        RECT -265.890 -175.735 -265.720 -175.135 ;
        RECT -264.060 -175.135 -263.365 -174.505 ;
        RECT -264.060 -175.735 -263.890 -175.135 ;
        RECT -263.720 -175.575 -263.385 -175.325 ;
        RECT -261.025 -175.485 -260.695 -174.505 ;
        RECT -259.165 -175.485 -258.835 -174.505 ;
        RECT -256.495 -175.135 -255.800 -174.505 ;
        RECT -269.020 -176.715 -268.325 -176.085 ;
        RECT -265.985 -176.715 -265.655 -175.735 ;
        RECT -264.125 -176.715 -263.795 -175.735 ;
        RECT -261.435 -175.895 -261.100 -175.645 ;
        RECT -260.930 -176.085 -260.760 -175.485 ;
        RECT -261.455 -176.715 -260.760 -176.085 ;
        RECT -259.100 -176.085 -258.930 -175.485 ;
        RECT -256.475 -175.575 -256.140 -175.325 ;
        RECT -258.760 -175.895 -258.425 -175.645 ;
        RECT -255.970 -175.735 -255.800 -175.135 ;
        RECT -254.140 -175.135 -253.445 -174.505 ;
        RECT -254.140 -175.735 -253.970 -175.135 ;
        RECT -253.800 -175.575 -253.465 -175.325 ;
        RECT -251.105 -175.485 -250.775 -174.505 ;
        RECT -249.245 -175.485 -248.915 -174.505 ;
        RECT -246.575 -175.135 -245.880 -174.505 ;
        RECT -259.100 -176.715 -258.405 -176.085 ;
        RECT -256.065 -176.715 -255.735 -175.735 ;
        RECT -254.205 -176.715 -253.875 -175.735 ;
        RECT -251.515 -175.895 -251.180 -175.645 ;
        RECT -251.010 -176.085 -250.840 -175.485 ;
        RECT -251.535 -176.715 -250.840 -176.085 ;
        RECT -249.180 -176.085 -249.010 -175.485 ;
        RECT -246.555 -175.575 -246.220 -175.325 ;
        RECT -248.840 -175.895 -248.505 -175.645 ;
        RECT -246.050 -175.735 -245.880 -175.135 ;
        RECT -244.220 -175.135 -243.525 -174.505 ;
        RECT -244.220 -175.735 -244.050 -175.135 ;
        RECT -243.880 -175.575 -243.545 -175.325 ;
        RECT -241.185 -175.485 -240.855 -174.505 ;
        RECT -239.325 -175.485 -238.995 -174.505 ;
        RECT -236.655 -175.135 -235.960 -174.505 ;
        RECT -249.180 -176.715 -248.485 -176.085 ;
        RECT -246.145 -176.715 -245.815 -175.735 ;
        RECT -244.285 -176.715 -243.955 -175.735 ;
        RECT -241.595 -175.895 -241.260 -175.645 ;
        RECT -241.090 -176.085 -240.920 -175.485 ;
        RECT -241.615 -176.715 -240.920 -176.085 ;
        RECT -239.260 -176.085 -239.090 -175.485 ;
        RECT -236.635 -175.575 -236.300 -175.325 ;
        RECT -238.920 -175.895 -238.585 -175.645 ;
        RECT -236.130 -175.735 -235.960 -175.135 ;
        RECT -234.300 -175.135 -233.605 -174.505 ;
        RECT -234.300 -175.735 -234.130 -175.135 ;
        RECT -233.960 -175.575 -233.625 -175.325 ;
        RECT -231.265 -175.485 -230.935 -174.505 ;
        RECT -229.405 -175.485 -229.075 -174.505 ;
        RECT -226.735 -175.135 -226.040 -174.505 ;
        RECT -239.260 -176.715 -238.565 -176.085 ;
        RECT -236.225 -176.715 -235.895 -175.735 ;
        RECT -234.365 -176.715 -234.035 -175.735 ;
        RECT -231.675 -175.895 -231.340 -175.645 ;
        RECT -231.170 -176.085 -231.000 -175.485 ;
        RECT -231.695 -176.715 -231.000 -176.085 ;
        RECT -229.340 -176.085 -229.170 -175.485 ;
        RECT -226.715 -175.575 -226.380 -175.325 ;
        RECT -229.000 -175.895 -228.665 -175.645 ;
        RECT -226.210 -175.735 -226.040 -175.135 ;
        RECT -224.380 -175.135 -223.685 -174.505 ;
        RECT -224.380 -175.735 -224.210 -175.135 ;
        RECT -224.040 -175.575 -223.705 -175.325 ;
        RECT -221.345 -175.485 -221.015 -174.505 ;
        RECT -219.485 -175.485 -219.155 -174.505 ;
        RECT -216.815 -175.135 -216.120 -174.505 ;
        RECT -229.340 -176.715 -228.645 -176.085 ;
        RECT -226.305 -176.715 -225.975 -175.735 ;
        RECT -224.445 -176.715 -224.115 -175.735 ;
        RECT -221.755 -175.895 -221.420 -175.645 ;
        RECT -221.250 -176.085 -221.080 -175.485 ;
        RECT -221.775 -176.715 -221.080 -176.085 ;
        RECT -219.420 -176.085 -219.250 -175.485 ;
        RECT -216.795 -175.575 -216.460 -175.325 ;
        RECT -219.080 -175.895 -218.745 -175.645 ;
        RECT -216.290 -175.735 -216.120 -175.135 ;
        RECT -214.460 -175.135 -213.765 -174.505 ;
        RECT -214.460 -175.735 -214.290 -175.135 ;
        RECT -214.120 -175.575 -213.785 -175.325 ;
        RECT -211.425 -175.485 -211.095 -174.505 ;
        RECT -209.565 -175.485 -209.235 -174.505 ;
        RECT -206.895 -175.135 -206.200 -174.505 ;
        RECT -219.420 -176.715 -218.725 -176.085 ;
        RECT -216.385 -176.715 -216.055 -175.735 ;
        RECT -214.525 -176.715 -214.195 -175.735 ;
        RECT -211.835 -175.895 -211.500 -175.645 ;
        RECT -211.330 -176.085 -211.160 -175.485 ;
        RECT -211.855 -176.715 -211.160 -176.085 ;
        RECT -209.500 -176.085 -209.330 -175.485 ;
        RECT -206.875 -175.575 -206.540 -175.325 ;
        RECT -209.160 -175.895 -208.825 -175.645 ;
        RECT -206.370 -175.735 -206.200 -175.135 ;
        RECT -204.540 -175.135 -203.845 -174.505 ;
        RECT -204.540 -175.735 -204.370 -175.135 ;
        RECT -204.200 -175.575 -203.865 -175.325 ;
        RECT -201.505 -175.485 -201.175 -174.505 ;
        RECT -199.645 -175.485 -199.315 -174.505 ;
        RECT -196.975 -175.135 -196.280 -174.505 ;
        RECT -209.500 -176.715 -208.805 -176.085 ;
        RECT -206.465 -176.715 -206.135 -175.735 ;
        RECT -204.605 -176.715 -204.275 -175.735 ;
        RECT -201.915 -175.895 -201.580 -175.645 ;
        RECT -201.410 -176.085 -201.240 -175.485 ;
        RECT -201.935 -176.715 -201.240 -176.085 ;
        RECT -199.580 -176.085 -199.410 -175.485 ;
        RECT -196.955 -175.575 -196.620 -175.325 ;
        RECT -199.240 -175.895 -198.905 -175.645 ;
        RECT -196.450 -175.735 -196.280 -175.135 ;
        RECT -194.620 -175.135 -193.925 -174.505 ;
        RECT -194.620 -175.735 -194.450 -175.135 ;
        RECT -194.280 -175.575 -193.945 -175.325 ;
        RECT -191.585 -175.485 -191.255 -174.505 ;
        RECT -189.725 -175.485 -189.395 -174.505 ;
        RECT -187.055 -175.135 -186.360 -174.505 ;
        RECT -199.580 -176.715 -198.885 -176.085 ;
        RECT -196.545 -176.715 -196.215 -175.735 ;
        RECT -194.685 -176.715 -194.355 -175.735 ;
        RECT -191.995 -175.895 -191.660 -175.645 ;
        RECT -191.490 -176.085 -191.320 -175.485 ;
        RECT -192.015 -176.715 -191.320 -176.085 ;
        RECT -189.660 -176.085 -189.490 -175.485 ;
        RECT -187.035 -175.575 -186.700 -175.325 ;
        RECT -189.320 -175.895 -188.985 -175.645 ;
        RECT -186.530 -175.735 -186.360 -175.135 ;
        RECT -184.700 -175.135 -184.005 -174.505 ;
        RECT -184.700 -175.735 -184.530 -175.135 ;
        RECT -184.360 -175.575 -184.025 -175.325 ;
        RECT -181.665 -175.485 -181.335 -174.505 ;
        RECT -179.805 -175.485 -179.475 -174.505 ;
        RECT -177.135 -175.135 -176.440 -174.505 ;
        RECT -189.660 -176.715 -188.965 -176.085 ;
        RECT -186.625 -176.715 -186.295 -175.735 ;
        RECT -184.765 -176.715 -184.435 -175.735 ;
        RECT -182.075 -175.895 -181.740 -175.645 ;
        RECT -181.570 -176.085 -181.400 -175.485 ;
        RECT -182.095 -176.715 -181.400 -176.085 ;
        RECT -179.740 -176.085 -179.570 -175.485 ;
        RECT -177.115 -175.575 -176.780 -175.325 ;
        RECT -179.400 -175.895 -179.065 -175.645 ;
        RECT -176.610 -175.735 -176.440 -175.135 ;
        RECT -174.780 -175.135 -174.085 -174.505 ;
        RECT -174.780 -175.735 -174.610 -175.135 ;
        RECT -174.440 -175.575 -174.105 -175.325 ;
        RECT -171.745 -175.485 -171.415 -174.505 ;
        RECT -169.885 -175.485 -169.555 -174.505 ;
        RECT -167.215 -175.135 -166.520 -174.505 ;
        RECT -179.740 -176.715 -179.045 -176.085 ;
        RECT -176.705 -176.715 -176.375 -175.735 ;
        RECT -174.845 -176.715 -174.515 -175.735 ;
        RECT -172.155 -175.895 -171.820 -175.645 ;
        RECT -171.650 -176.085 -171.480 -175.485 ;
        RECT -172.175 -176.715 -171.480 -176.085 ;
        RECT -169.820 -176.085 -169.650 -175.485 ;
        RECT -167.195 -175.575 -166.860 -175.325 ;
        RECT -169.480 -175.895 -169.145 -175.645 ;
        RECT -166.690 -175.735 -166.520 -175.135 ;
        RECT -164.860 -175.135 -164.165 -174.505 ;
        RECT -164.860 -175.735 -164.690 -175.135 ;
        RECT -164.520 -175.575 -164.185 -175.325 ;
        RECT -161.825 -175.485 -161.495 -174.505 ;
        RECT -159.965 -175.485 -159.635 -174.505 ;
        RECT -157.295 -175.135 -156.600 -174.505 ;
        RECT -169.820 -176.715 -169.125 -176.085 ;
        RECT -166.785 -176.715 -166.455 -175.735 ;
        RECT -164.925 -176.715 -164.595 -175.735 ;
        RECT -162.235 -175.895 -161.900 -175.645 ;
        RECT -161.730 -176.085 -161.560 -175.485 ;
        RECT -162.255 -176.715 -161.560 -176.085 ;
        RECT -159.900 -176.085 -159.730 -175.485 ;
        RECT -157.275 -175.575 -156.940 -175.325 ;
        RECT -159.560 -175.895 -159.225 -175.645 ;
        RECT -156.770 -175.735 -156.600 -175.135 ;
        RECT -154.940 -175.135 -154.245 -174.505 ;
        RECT -154.940 -175.735 -154.770 -175.135 ;
        RECT -154.600 -175.575 -154.265 -175.325 ;
        RECT -151.905 -175.485 -151.575 -174.505 ;
        RECT -150.045 -175.485 -149.715 -174.505 ;
        RECT -147.375 -175.135 -146.680 -174.505 ;
        RECT -159.900 -176.715 -159.205 -176.085 ;
        RECT -156.865 -176.715 -156.535 -175.735 ;
        RECT -155.005 -176.715 -154.675 -175.735 ;
        RECT -152.315 -175.895 -151.980 -175.645 ;
        RECT -151.810 -176.085 -151.640 -175.485 ;
        RECT -152.335 -176.715 -151.640 -176.085 ;
        RECT -149.980 -176.085 -149.810 -175.485 ;
        RECT -147.355 -175.575 -147.020 -175.325 ;
        RECT -149.640 -175.895 -149.305 -175.645 ;
        RECT -146.850 -175.735 -146.680 -175.135 ;
        RECT -145.020 -175.135 -144.325 -174.505 ;
        RECT -145.020 -175.735 -144.850 -175.135 ;
        RECT -144.680 -175.575 -144.345 -175.325 ;
        RECT -141.985 -175.485 -141.655 -174.505 ;
        RECT -140.125 -175.485 -139.795 -174.505 ;
        RECT -137.455 -175.135 -136.760 -174.505 ;
        RECT -149.980 -176.715 -149.285 -176.085 ;
        RECT -146.945 -176.715 -146.615 -175.735 ;
        RECT -145.085 -176.715 -144.755 -175.735 ;
        RECT -142.395 -175.895 -142.060 -175.645 ;
        RECT -141.890 -176.085 -141.720 -175.485 ;
        RECT -142.415 -176.715 -141.720 -176.085 ;
        RECT -140.060 -176.085 -139.890 -175.485 ;
        RECT -137.435 -175.575 -137.100 -175.325 ;
        RECT -139.720 -175.895 -139.385 -175.645 ;
        RECT -136.930 -175.735 -136.760 -175.135 ;
        RECT -135.100 -175.135 -134.405 -174.505 ;
        RECT -135.100 -175.735 -134.930 -175.135 ;
        RECT -134.760 -175.575 -134.425 -175.325 ;
        RECT -132.065 -175.485 -131.735 -174.505 ;
        RECT -130.205 -175.485 -129.875 -174.505 ;
        RECT -127.535 -175.135 -126.840 -174.505 ;
        RECT -140.060 -176.715 -139.365 -176.085 ;
        RECT -137.025 -176.715 -136.695 -175.735 ;
        RECT -135.165 -176.715 -134.835 -175.735 ;
        RECT -132.475 -175.895 -132.140 -175.645 ;
        RECT -131.970 -176.085 -131.800 -175.485 ;
        RECT -132.495 -176.715 -131.800 -176.085 ;
        RECT -130.140 -176.085 -129.970 -175.485 ;
        RECT -127.515 -175.575 -127.180 -175.325 ;
        RECT -129.800 -175.895 -129.465 -175.645 ;
        RECT -127.010 -175.735 -126.840 -175.135 ;
        RECT -125.180 -175.135 -124.485 -174.505 ;
        RECT -125.180 -175.735 -125.010 -175.135 ;
        RECT -124.840 -175.575 -124.505 -175.325 ;
        RECT -122.145 -175.485 -121.815 -174.505 ;
        RECT -120.285 -175.485 -119.955 -174.505 ;
        RECT -117.615 -175.135 -116.920 -174.505 ;
        RECT -130.140 -176.715 -129.445 -176.085 ;
        RECT -127.105 -176.715 -126.775 -175.735 ;
        RECT -125.245 -176.715 -124.915 -175.735 ;
        RECT -122.555 -175.895 -122.220 -175.645 ;
        RECT -122.050 -176.085 -121.880 -175.485 ;
        RECT -122.575 -176.715 -121.880 -176.085 ;
        RECT -120.220 -176.085 -120.050 -175.485 ;
        RECT -117.595 -175.575 -117.260 -175.325 ;
        RECT -119.880 -175.895 -119.545 -175.645 ;
        RECT -117.090 -175.735 -116.920 -175.135 ;
        RECT -115.260 -175.135 -114.565 -174.505 ;
        RECT -115.260 -175.735 -115.090 -175.135 ;
        RECT -114.920 -175.575 -114.585 -175.325 ;
        RECT -112.225 -175.485 -111.895 -174.505 ;
        RECT -110.365 -175.485 -110.035 -174.505 ;
        RECT -107.695 -175.135 -107.000 -174.505 ;
        RECT -120.220 -176.715 -119.525 -176.085 ;
        RECT -117.185 -176.715 -116.855 -175.735 ;
        RECT -115.325 -176.715 -114.995 -175.735 ;
        RECT -112.635 -175.895 -112.300 -175.645 ;
        RECT -112.130 -176.085 -111.960 -175.485 ;
        RECT -112.655 -176.715 -111.960 -176.085 ;
        RECT -110.300 -176.085 -110.130 -175.485 ;
        RECT -107.675 -175.575 -107.340 -175.325 ;
        RECT -109.960 -175.895 -109.625 -175.645 ;
        RECT -107.170 -175.735 -107.000 -175.135 ;
        RECT -105.340 -175.135 -104.645 -174.505 ;
        RECT -105.340 -175.735 -105.170 -175.135 ;
        RECT -105.000 -175.575 -104.665 -175.325 ;
        RECT -102.305 -175.485 -101.975 -174.505 ;
        RECT -100.445 -175.485 -100.115 -174.505 ;
        RECT -97.775 -175.135 -97.080 -174.505 ;
        RECT -110.300 -176.715 -109.605 -176.085 ;
        RECT -107.265 -176.715 -106.935 -175.735 ;
        RECT -105.405 -176.715 -105.075 -175.735 ;
        RECT -102.715 -175.895 -102.380 -175.645 ;
        RECT -102.210 -176.085 -102.040 -175.485 ;
        RECT -102.735 -176.715 -102.040 -176.085 ;
        RECT -100.380 -176.085 -100.210 -175.485 ;
        RECT -97.755 -175.575 -97.420 -175.325 ;
        RECT -100.040 -175.895 -99.705 -175.645 ;
        RECT -97.250 -175.735 -97.080 -175.135 ;
        RECT -95.420 -175.135 -94.725 -174.505 ;
        RECT -95.420 -175.735 -95.250 -175.135 ;
        RECT -95.080 -175.575 -94.745 -175.325 ;
        RECT -92.385 -175.485 -92.055 -174.505 ;
        RECT -90.525 -175.485 -90.195 -174.505 ;
        RECT -87.855 -175.135 -87.160 -174.505 ;
        RECT -100.380 -176.715 -99.685 -176.085 ;
        RECT -97.345 -176.715 -97.015 -175.735 ;
        RECT -95.485 -176.715 -95.155 -175.735 ;
        RECT -92.795 -175.895 -92.460 -175.645 ;
        RECT -92.290 -176.085 -92.120 -175.485 ;
        RECT -92.815 -176.715 -92.120 -176.085 ;
        RECT -90.460 -176.085 -90.290 -175.485 ;
        RECT -87.835 -175.575 -87.500 -175.325 ;
        RECT -90.120 -175.895 -89.785 -175.645 ;
        RECT -87.330 -175.735 -87.160 -175.135 ;
        RECT -85.500 -175.135 -84.805 -174.505 ;
        RECT -85.500 -175.735 -85.330 -175.135 ;
        RECT -85.160 -175.575 -84.825 -175.325 ;
        RECT -82.465 -175.485 -82.135 -174.505 ;
        RECT -80.605 -175.485 -80.275 -174.505 ;
        RECT -77.935 -175.135 -77.240 -174.505 ;
        RECT -90.460 -176.715 -89.765 -176.085 ;
        RECT -87.425 -176.715 -87.095 -175.735 ;
        RECT -85.565 -176.715 -85.235 -175.735 ;
        RECT -82.875 -175.895 -82.540 -175.645 ;
        RECT -82.370 -176.085 -82.200 -175.485 ;
        RECT -82.895 -176.715 -82.200 -176.085 ;
        RECT -80.540 -176.085 -80.370 -175.485 ;
        RECT -77.915 -175.575 -77.580 -175.325 ;
        RECT -80.200 -175.895 -79.865 -175.645 ;
        RECT -77.410 -175.735 -77.240 -175.135 ;
        RECT -75.580 -175.135 -74.885 -174.505 ;
        RECT -75.580 -175.735 -75.410 -175.135 ;
        RECT -75.240 -175.575 -74.905 -175.325 ;
        RECT -72.545 -175.485 -72.215 -174.505 ;
        RECT -70.685 -175.485 -70.355 -174.505 ;
        RECT -68.015 -175.135 -67.320 -174.505 ;
        RECT -80.540 -176.715 -79.845 -176.085 ;
        RECT -77.505 -176.715 -77.175 -175.735 ;
        RECT -75.645 -176.715 -75.315 -175.735 ;
        RECT -72.955 -175.895 -72.620 -175.645 ;
        RECT -72.450 -176.085 -72.280 -175.485 ;
        RECT -72.975 -176.715 -72.280 -176.085 ;
        RECT -70.620 -176.085 -70.450 -175.485 ;
        RECT -67.995 -175.575 -67.660 -175.325 ;
        RECT -70.280 -175.895 -69.945 -175.645 ;
        RECT -67.490 -175.735 -67.320 -175.135 ;
        RECT -65.660 -175.135 -64.965 -174.505 ;
        RECT -65.660 -175.735 -65.490 -175.135 ;
        RECT -65.320 -175.575 -64.985 -175.325 ;
        RECT -62.625 -175.485 -62.295 -174.505 ;
        RECT -60.765 -175.485 -60.435 -174.505 ;
        RECT -58.095 -175.135 -57.400 -174.505 ;
        RECT -70.620 -176.715 -69.925 -176.085 ;
        RECT -67.585 -176.715 -67.255 -175.735 ;
        RECT -65.725 -176.715 -65.395 -175.735 ;
        RECT -63.035 -175.895 -62.700 -175.645 ;
        RECT -62.530 -176.085 -62.360 -175.485 ;
        RECT -63.055 -176.715 -62.360 -176.085 ;
        RECT -60.700 -176.085 -60.530 -175.485 ;
        RECT -58.075 -175.575 -57.740 -175.325 ;
        RECT -60.360 -175.895 -60.025 -175.645 ;
        RECT -57.570 -175.735 -57.400 -175.135 ;
        RECT -55.740 -175.135 -55.045 -174.505 ;
        RECT -55.740 -175.735 -55.570 -175.135 ;
        RECT -55.400 -175.575 -55.065 -175.325 ;
        RECT -52.705 -175.485 -52.375 -174.505 ;
        RECT -50.845 -175.485 -50.515 -174.505 ;
        RECT -48.175 -175.135 -47.480 -174.505 ;
        RECT -60.700 -176.715 -60.005 -176.085 ;
        RECT -57.665 -176.715 -57.335 -175.735 ;
        RECT -55.805 -176.715 -55.475 -175.735 ;
        RECT -53.115 -175.895 -52.780 -175.645 ;
        RECT -52.610 -176.085 -52.440 -175.485 ;
        RECT -53.135 -176.715 -52.440 -176.085 ;
        RECT -50.780 -176.085 -50.610 -175.485 ;
        RECT -48.155 -175.575 -47.820 -175.325 ;
        RECT -50.440 -175.895 -50.105 -175.645 ;
        RECT -47.650 -175.735 -47.480 -175.135 ;
        RECT -45.820 -175.135 -45.125 -174.505 ;
        RECT -45.820 -175.735 -45.650 -175.135 ;
        RECT -45.480 -175.575 -45.145 -175.325 ;
        RECT -42.785 -175.485 -42.455 -174.505 ;
        RECT -40.925 -175.485 -40.595 -174.505 ;
        RECT -38.255 -175.135 -37.560 -174.505 ;
        RECT -50.780 -176.715 -50.085 -176.085 ;
        RECT -47.745 -176.715 -47.415 -175.735 ;
        RECT -45.885 -176.715 -45.555 -175.735 ;
        RECT -43.195 -175.895 -42.860 -175.645 ;
        RECT -42.690 -176.085 -42.520 -175.485 ;
        RECT -43.215 -176.715 -42.520 -176.085 ;
        RECT -40.860 -176.085 -40.690 -175.485 ;
        RECT -38.235 -175.575 -37.900 -175.325 ;
        RECT -40.520 -175.895 -40.185 -175.645 ;
        RECT -37.730 -175.735 -37.560 -175.135 ;
        RECT -35.900 -175.135 -35.205 -174.505 ;
        RECT -35.900 -175.735 -35.730 -175.135 ;
        RECT -35.560 -175.575 -35.225 -175.325 ;
        RECT -32.865 -175.485 -32.535 -174.505 ;
        RECT -31.005 -175.485 -30.675 -174.505 ;
        RECT -28.335 -175.135 -27.640 -174.505 ;
        RECT -40.860 -176.715 -40.165 -176.085 ;
        RECT -37.825 -176.715 -37.495 -175.735 ;
        RECT -35.965 -176.715 -35.635 -175.735 ;
        RECT -33.275 -175.895 -32.940 -175.645 ;
        RECT -32.770 -176.085 -32.600 -175.485 ;
        RECT -33.295 -176.715 -32.600 -176.085 ;
        RECT -30.940 -176.085 -30.770 -175.485 ;
        RECT -28.315 -175.575 -27.980 -175.325 ;
        RECT -30.600 -175.895 -30.265 -175.645 ;
        RECT -27.810 -175.735 -27.640 -175.135 ;
        RECT -25.980 -175.135 -25.285 -174.505 ;
        RECT -25.980 -175.735 -25.810 -175.135 ;
        RECT -25.640 -175.575 -25.305 -175.325 ;
        RECT -22.945 -175.485 -22.615 -174.505 ;
        RECT -21.085 -175.485 -20.755 -174.505 ;
        RECT -18.415 -175.135 -17.720 -174.505 ;
        RECT -30.940 -176.715 -30.245 -176.085 ;
        RECT -27.905 -176.715 -27.575 -175.735 ;
        RECT -26.045 -176.715 -25.715 -175.735 ;
        RECT -23.355 -175.895 -23.020 -175.645 ;
        RECT -22.850 -176.085 -22.680 -175.485 ;
        RECT -23.375 -176.715 -22.680 -176.085 ;
        RECT -21.020 -176.085 -20.850 -175.485 ;
        RECT -18.395 -175.575 -18.060 -175.325 ;
        RECT -20.680 -175.895 -20.345 -175.645 ;
        RECT -17.890 -175.735 -17.720 -175.135 ;
        RECT -16.060 -175.135 -15.365 -174.505 ;
        RECT -16.060 -175.735 -15.890 -175.135 ;
        RECT -15.720 -175.575 -15.385 -175.325 ;
        RECT -13.025 -175.485 -12.695 -174.505 ;
        RECT -11.165 -175.485 -10.835 -174.505 ;
        RECT -8.495 -175.135 -7.800 -174.505 ;
        RECT -21.020 -176.715 -20.325 -176.085 ;
        RECT -17.985 -176.715 -17.655 -175.735 ;
        RECT -16.125 -176.715 -15.795 -175.735 ;
        RECT -13.435 -175.895 -13.100 -175.645 ;
        RECT -12.930 -176.085 -12.760 -175.485 ;
        RECT -13.455 -176.715 -12.760 -176.085 ;
        RECT -11.100 -176.085 -10.930 -175.485 ;
        RECT -8.475 -175.575 -8.140 -175.325 ;
        RECT -10.760 -175.895 -10.425 -175.645 ;
        RECT -7.970 -175.735 -7.800 -175.135 ;
        RECT -6.140 -175.135 -5.445 -174.505 ;
        RECT -6.140 -175.735 -5.970 -175.135 ;
        RECT -5.800 -175.575 -5.465 -175.325 ;
        RECT -3.105 -175.485 -2.775 -174.505 ;
        RECT -1.245 -175.485 -0.915 -174.505 ;
        RECT 1.425 -175.135 2.120 -174.505 ;
        RECT -11.100 -176.715 -10.405 -176.085 ;
        RECT -8.065 -176.715 -7.735 -175.735 ;
        RECT -6.205 -176.715 -5.875 -175.735 ;
        RECT -3.515 -175.895 -3.180 -175.645 ;
        RECT -3.010 -176.085 -2.840 -175.485 ;
        RECT -3.535 -176.715 -2.840 -176.085 ;
        RECT -1.180 -176.085 -1.010 -175.485 ;
        RECT 1.445 -175.575 1.780 -175.325 ;
        RECT -0.840 -175.895 -0.505 -175.645 ;
        RECT 1.950 -175.735 2.120 -175.135 ;
        RECT 3.780 -175.135 4.475 -174.505 ;
        RECT 3.780 -175.735 3.950 -175.135 ;
        RECT 4.120 -175.575 4.455 -175.325 ;
        RECT 6.815 -175.485 7.145 -174.505 ;
        RECT 8.675 -175.485 9.005 -174.505 ;
        RECT 11.345 -175.135 12.040 -174.505 ;
        RECT -1.180 -176.715 -0.485 -176.085 ;
        RECT 1.855 -176.715 2.185 -175.735 ;
        RECT 3.715 -176.715 4.045 -175.735 ;
        RECT 6.405 -175.895 6.740 -175.645 ;
        RECT 6.910 -176.085 7.080 -175.485 ;
        RECT 6.385 -176.715 7.080 -176.085 ;
        RECT 8.740 -176.085 8.910 -175.485 ;
        RECT 11.365 -175.575 11.700 -175.325 ;
        RECT 9.080 -175.895 9.415 -175.645 ;
        RECT 11.870 -175.735 12.040 -175.135 ;
        RECT 13.700 -175.135 14.395 -174.505 ;
        RECT 13.700 -175.735 13.870 -175.135 ;
        RECT 14.040 -175.575 14.375 -175.325 ;
        RECT 16.735 -175.485 17.065 -174.505 ;
        RECT 18.595 -175.485 18.925 -174.505 ;
        RECT 21.265 -175.135 21.960 -174.505 ;
        RECT 22.165 -175.135 22.475 -174.335 ;
        RECT 22.645 -175.060 22.935 -174.335 ;
        RECT 8.740 -176.715 9.435 -176.085 ;
        RECT 11.775 -176.715 12.105 -175.735 ;
        RECT 13.635 -176.715 13.965 -175.735 ;
        RECT 16.325 -175.895 16.660 -175.645 ;
        RECT 16.830 -176.085 17.000 -175.485 ;
        RECT 16.305 -176.715 17.000 -176.085 ;
        RECT 18.660 -176.085 18.830 -175.485 ;
        RECT 21.285 -175.575 21.620 -175.325 ;
        RECT 19.000 -175.895 19.335 -175.645 ;
        RECT 21.790 -175.735 21.960 -175.135 ;
        RECT 18.660 -176.715 19.355 -176.085 ;
        RECT 21.695 -176.715 22.025 -175.735 ;
        RECT -294.880 -177.055 -293.040 -176.885 ;
        RECT -293.495 -178.440 -293.205 -177.730 ;
        RECT -292.965 -177.925 -292.795 -177.400 ;
        RECT -292.625 -177.745 -292.075 -177.575 ;
        RECT -292.965 -178.255 -292.415 -177.925 ;
        RECT -292.245 -178.070 -292.075 -177.745 ;
        RECT -291.895 -177.845 -291.525 -177.505 ;
        RECT -291.345 -177.745 -290.415 -177.565 ;
        RECT -288.965 -177.745 -288.035 -177.565 ;
        RECT -291.345 -178.070 -291.175 -177.745 ;
        RECT -292.245 -178.240 -291.175 -178.070 ;
        RECT -288.205 -178.070 -288.035 -177.745 ;
        RECT -287.855 -177.845 -287.485 -177.505 ;
        RECT -287.305 -177.745 -286.755 -177.575 ;
        RECT -282.705 -177.745 -282.155 -177.575 ;
        RECT -287.305 -178.070 -287.135 -177.745 ;
        RECT -288.205 -178.240 -287.135 -178.070 ;
        RECT -282.325 -178.070 -282.155 -177.745 ;
        RECT -281.975 -177.845 -281.605 -177.505 ;
        RECT -281.425 -177.745 -280.495 -177.565 ;
        RECT -279.045 -177.745 -278.115 -177.565 ;
        RECT -281.425 -178.070 -281.255 -177.745 ;
        RECT -282.325 -178.240 -281.255 -178.070 ;
        RECT -278.285 -178.070 -278.115 -177.745 ;
        RECT -277.935 -177.845 -277.565 -177.505 ;
        RECT -277.385 -177.745 -276.835 -177.575 ;
        RECT -272.785 -177.745 -272.235 -177.575 ;
        RECT -277.385 -178.070 -277.215 -177.745 ;
        RECT -278.285 -178.240 -277.215 -178.070 ;
        RECT -272.405 -178.070 -272.235 -177.745 ;
        RECT -272.055 -177.845 -271.685 -177.505 ;
        RECT -271.505 -177.745 -270.575 -177.565 ;
        RECT -269.125 -177.745 -268.195 -177.565 ;
        RECT -271.505 -178.070 -271.335 -177.745 ;
        RECT -272.405 -178.240 -271.335 -178.070 ;
        RECT -268.365 -178.070 -268.195 -177.745 ;
        RECT -268.015 -177.845 -267.645 -177.505 ;
        RECT -267.465 -177.745 -266.915 -177.575 ;
        RECT -262.865 -177.745 -262.315 -177.575 ;
        RECT -267.465 -178.070 -267.295 -177.745 ;
        RECT -268.365 -178.240 -267.295 -178.070 ;
        RECT -262.485 -178.070 -262.315 -177.745 ;
        RECT -262.135 -177.845 -261.765 -177.505 ;
        RECT -261.585 -177.745 -260.655 -177.565 ;
        RECT -259.205 -177.745 -258.275 -177.565 ;
        RECT -261.585 -178.070 -261.415 -177.745 ;
        RECT -262.485 -178.240 -261.415 -178.070 ;
        RECT -258.445 -178.070 -258.275 -177.745 ;
        RECT -258.095 -177.845 -257.725 -177.505 ;
        RECT -257.545 -177.745 -256.995 -177.575 ;
        RECT -252.945 -177.745 -252.395 -177.575 ;
        RECT -257.545 -178.070 -257.375 -177.745 ;
        RECT -258.445 -178.240 -257.375 -178.070 ;
        RECT -252.565 -178.070 -252.395 -177.745 ;
        RECT -252.215 -177.845 -251.845 -177.505 ;
        RECT -251.665 -177.745 -250.735 -177.565 ;
        RECT -249.285 -177.745 -248.355 -177.565 ;
        RECT -251.665 -178.070 -251.495 -177.745 ;
        RECT -252.565 -178.240 -251.495 -178.070 ;
        RECT -248.525 -178.070 -248.355 -177.745 ;
        RECT -248.175 -177.845 -247.805 -177.505 ;
        RECT -247.625 -177.745 -247.075 -177.575 ;
        RECT -243.025 -177.745 -242.475 -177.575 ;
        RECT -247.625 -178.070 -247.455 -177.745 ;
        RECT -248.525 -178.240 -247.455 -178.070 ;
        RECT -242.645 -178.070 -242.475 -177.745 ;
        RECT -242.295 -177.845 -241.925 -177.505 ;
        RECT -241.745 -177.745 -240.815 -177.565 ;
        RECT -239.365 -177.745 -238.435 -177.565 ;
        RECT -241.745 -178.070 -241.575 -177.745 ;
        RECT -242.645 -178.240 -241.575 -178.070 ;
        RECT -238.605 -178.070 -238.435 -177.745 ;
        RECT -238.255 -177.845 -237.885 -177.505 ;
        RECT -237.705 -177.745 -237.155 -177.575 ;
        RECT -233.105 -177.745 -232.555 -177.575 ;
        RECT -237.705 -178.070 -237.535 -177.745 ;
        RECT -238.605 -178.240 -237.535 -178.070 ;
        RECT -232.725 -178.070 -232.555 -177.745 ;
        RECT -232.375 -177.845 -232.005 -177.505 ;
        RECT -231.825 -177.745 -230.895 -177.565 ;
        RECT -229.445 -177.745 -228.515 -177.565 ;
        RECT -231.825 -178.070 -231.655 -177.745 ;
        RECT -232.725 -178.240 -231.655 -178.070 ;
        RECT -228.685 -178.070 -228.515 -177.745 ;
        RECT -228.335 -177.845 -227.965 -177.505 ;
        RECT -227.785 -177.745 -227.235 -177.575 ;
        RECT -223.185 -177.745 -222.635 -177.575 ;
        RECT -227.785 -178.070 -227.615 -177.745 ;
        RECT -228.685 -178.240 -227.615 -178.070 ;
        RECT -222.805 -178.070 -222.635 -177.745 ;
        RECT -222.455 -177.845 -222.085 -177.505 ;
        RECT -221.905 -177.745 -220.975 -177.565 ;
        RECT -219.525 -177.745 -218.595 -177.565 ;
        RECT -221.905 -178.070 -221.735 -177.745 ;
        RECT -222.805 -178.240 -221.735 -178.070 ;
        RECT -218.765 -178.070 -218.595 -177.745 ;
        RECT -218.415 -177.845 -218.045 -177.505 ;
        RECT -217.865 -177.745 -217.315 -177.575 ;
        RECT -213.265 -177.745 -212.715 -177.575 ;
        RECT -217.865 -178.070 -217.695 -177.745 ;
        RECT -218.765 -178.240 -217.695 -178.070 ;
        RECT -212.885 -178.070 -212.715 -177.745 ;
        RECT -212.535 -177.845 -212.165 -177.505 ;
        RECT -211.985 -177.745 -211.055 -177.565 ;
        RECT -209.605 -177.745 -208.675 -177.565 ;
        RECT -211.985 -178.070 -211.815 -177.745 ;
        RECT -212.885 -178.240 -211.815 -178.070 ;
        RECT -208.845 -178.070 -208.675 -177.745 ;
        RECT -208.495 -177.845 -208.125 -177.505 ;
        RECT -207.945 -177.745 -207.395 -177.575 ;
        RECT -203.345 -177.745 -202.795 -177.575 ;
        RECT -207.945 -178.070 -207.775 -177.745 ;
        RECT -208.845 -178.240 -207.775 -178.070 ;
        RECT -202.965 -178.070 -202.795 -177.745 ;
        RECT -202.615 -177.845 -202.245 -177.505 ;
        RECT -202.065 -177.745 -201.135 -177.565 ;
        RECT -199.685 -177.745 -198.755 -177.565 ;
        RECT -202.065 -178.070 -201.895 -177.745 ;
        RECT -202.965 -178.240 -201.895 -178.070 ;
        RECT -198.925 -178.070 -198.755 -177.745 ;
        RECT -198.575 -177.845 -198.205 -177.505 ;
        RECT -198.025 -177.745 -197.475 -177.575 ;
        RECT -193.425 -177.745 -192.875 -177.575 ;
        RECT -198.025 -178.070 -197.855 -177.745 ;
        RECT -198.925 -178.240 -197.855 -178.070 ;
        RECT -193.045 -178.070 -192.875 -177.745 ;
        RECT -192.695 -177.845 -192.325 -177.505 ;
        RECT -192.145 -177.745 -191.215 -177.565 ;
        RECT -189.765 -177.745 -188.835 -177.565 ;
        RECT -192.145 -178.070 -191.975 -177.745 ;
        RECT -193.045 -178.240 -191.975 -178.070 ;
        RECT -189.005 -178.070 -188.835 -177.745 ;
        RECT -188.655 -177.845 -188.285 -177.505 ;
        RECT -188.105 -177.745 -187.555 -177.575 ;
        RECT -183.505 -177.745 -182.955 -177.575 ;
        RECT -188.105 -178.070 -187.935 -177.745 ;
        RECT -189.005 -178.240 -187.935 -178.070 ;
        RECT -183.125 -178.070 -182.955 -177.745 ;
        RECT -182.775 -177.845 -182.405 -177.505 ;
        RECT -182.225 -177.745 -181.295 -177.565 ;
        RECT -179.845 -177.745 -178.915 -177.565 ;
        RECT -182.225 -178.070 -182.055 -177.745 ;
        RECT -183.125 -178.240 -182.055 -178.070 ;
        RECT -179.085 -178.070 -178.915 -177.745 ;
        RECT -178.735 -177.845 -178.365 -177.505 ;
        RECT -178.185 -177.745 -177.635 -177.575 ;
        RECT -173.585 -177.745 -173.035 -177.575 ;
        RECT -178.185 -178.070 -178.015 -177.745 ;
        RECT -179.085 -178.240 -178.015 -178.070 ;
        RECT -173.205 -178.070 -173.035 -177.745 ;
        RECT -172.855 -177.845 -172.485 -177.505 ;
        RECT -172.305 -177.745 -171.375 -177.565 ;
        RECT -169.925 -177.745 -168.995 -177.565 ;
        RECT -172.305 -178.070 -172.135 -177.745 ;
        RECT -173.205 -178.240 -172.135 -178.070 ;
        RECT -169.165 -178.070 -168.995 -177.745 ;
        RECT -168.815 -177.845 -168.445 -177.505 ;
        RECT -168.265 -177.745 -167.715 -177.575 ;
        RECT -163.665 -177.745 -163.115 -177.575 ;
        RECT -168.265 -178.070 -168.095 -177.745 ;
        RECT -169.165 -178.240 -168.095 -178.070 ;
        RECT -163.285 -178.070 -163.115 -177.745 ;
        RECT -162.935 -177.845 -162.565 -177.505 ;
        RECT -162.385 -177.745 -161.455 -177.565 ;
        RECT -160.005 -177.745 -159.075 -177.565 ;
        RECT -162.385 -178.070 -162.215 -177.745 ;
        RECT -163.285 -178.240 -162.215 -178.070 ;
        RECT -159.245 -178.070 -159.075 -177.745 ;
        RECT -158.895 -177.845 -158.525 -177.505 ;
        RECT -158.345 -177.745 -157.795 -177.575 ;
        RECT -153.745 -177.745 -153.195 -177.575 ;
        RECT -158.345 -178.070 -158.175 -177.745 ;
        RECT -159.245 -178.240 -158.175 -178.070 ;
        RECT -153.365 -178.070 -153.195 -177.745 ;
        RECT -153.015 -177.845 -152.645 -177.505 ;
        RECT -152.465 -177.745 -151.535 -177.565 ;
        RECT -150.085 -177.745 -149.155 -177.565 ;
        RECT -152.465 -178.070 -152.295 -177.745 ;
        RECT -153.365 -178.240 -152.295 -178.070 ;
        RECT -149.325 -178.070 -149.155 -177.745 ;
        RECT -148.975 -177.845 -148.605 -177.505 ;
        RECT -148.425 -177.745 -147.875 -177.575 ;
        RECT -143.825 -177.745 -143.275 -177.575 ;
        RECT -148.425 -178.070 -148.255 -177.745 ;
        RECT -149.325 -178.240 -148.255 -178.070 ;
        RECT -143.445 -178.070 -143.275 -177.745 ;
        RECT -143.095 -177.845 -142.725 -177.505 ;
        RECT -142.545 -177.745 -141.615 -177.565 ;
        RECT -140.165 -177.745 -139.235 -177.565 ;
        RECT -142.545 -178.070 -142.375 -177.745 ;
        RECT -143.445 -178.240 -142.375 -178.070 ;
        RECT -139.405 -178.070 -139.235 -177.745 ;
        RECT -139.055 -177.845 -138.685 -177.505 ;
        RECT -138.505 -177.745 -137.955 -177.575 ;
        RECT -133.905 -177.745 -133.355 -177.575 ;
        RECT -138.505 -178.070 -138.335 -177.745 ;
        RECT -139.405 -178.240 -138.335 -178.070 ;
        RECT -133.525 -178.070 -133.355 -177.745 ;
        RECT -133.175 -177.845 -132.805 -177.505 ;
        RECT -132.625 -177.745 -131.695 -177.565 ;
        RECT -130.245 -177.745 -129.315 -177.565 ;
        RECT -132.625 -178.070 -132.455 -177.745 ;
        RECT -133.525 -178.240 -132.455 -178.070 ;
        RECT -129.485 -178.070 -129.315 -177.745 ;
        RECT -129.135 -177.845 -128.765 -177.505 ;
        RECT -128.585 -177.745 -128.035 -177.575 ;
        RECT -123.985 -177.745 -123.435 -177.575 ;
        RECT -128.585 -178.070 -128.415 -177.745 ;
        RECT -129.485 -178.240 -128.415 -178.070 ;
        RECT -123.605 -178.070 -123.435 -177.745 ;
        RECT -123.255 -177.845 -122.885 -177.505 ;
        RECT -122.705 -177.745 -121.775 -177.565 ;
        RECT -120.325 -177.745 -119.395 -177.565 ;
        RECT -122.705 -178.070 -122.535 -177.745 ;
        RECT -123.605 -178.240 -122.535 -178.070 ;
        RECT -119.565 -178.070 -119.395 -177.745 ;
        RECT -119.215 -177.845 -118.845 -177.505 ;
        RECT -118.665 -177.745 -118.115 -177.575 ;
        RECT -114.065 -177.745 -113.515 -177.575 ;
        RECT -118.665 -178.070 -118.495 -177.745 ;
        RECT -119.565 -178.240 -118.495 -178.070 ;
        RECT -113.685 -178.070 -113.515 -177.745 ;
        RECT -113.335 -177.845 -112.965 -177.505 ;
        RECT -112.785 -177.745 -111.855 -177.565 ;
        RECT -110.405 -177.745 -109.475 -177.565 ;
        RECT -112.785 -178.070 -112.615 -177.745 ;
        RECT -113.685 -178.240 -112.615 -178.070 ;
        RECT -109.645 -178.070 -109.475 -177.745 ;
        RECT -109.295 -177.845 -108.925 -177.505 ;
        RECT -108.745 -177.745 -108.195 -177.575 ;
        RECT -104.145 -177.745 -103.595 -177.575 ;
        RECT -108.745 -178.070 -108.575 -177.745 ;
        RECT -109.645 -178.240 -108.575 -178.070 ;
        RECT -103.765 -178.070 -103.595 -177.745 ;
        RECT -103.415 -177.845 -103.045 -177.505 ;
        RECT -102.865 -177.745 -101.935 -177.565 ;
        RECT -100.485 -177.745 -99.555 -177.565 ;
        RECT -102.865 -178.070 -102.695 -177.745 ;
        RECT -103.765 -178.240 -102.695 -178.070 ;
        RECT -99.725 -178.070 -99.555 -177.745 ;
        RECT -99.375 -177.845 -99.005 -177.505 ;
        RECT -98.825 -177.745 -98.275 -177.575 ;
        RECT -94.225 -177.745 -93.675 -177.575 ;
        RECT -98.825 -178.070 -98.655 -177.745 ;
        RECT -99.725 -178.240 -98.655 -178.070 ;
        RECT -93.845 -178.070 -93.675 -177.745 ;
        RECT -93.495 -177.845 -93.125 -177.505 ;
        RECT -92.945 -177.745 -92.015 -177.565 ;
        RECT -90.565 -177.745 -89.635 -177.565 ;
        RECT -92.945 -178.070 -92.775 -177.745 ;
        RECT -93.845 -178.240 -92.775 -178.070 ;
        RECT -89.805 -178.070 -89.635 -177.745 ;
        RECT -89.455 -177.845 -89.085 -177.505 ;
        RECT -88.905 -177.745 -88.355 -177.575 ;
        RECT -84.305 -177.745 -83.755 -177.575 ;
        RECT -88.905 -178.070 -88.735 -177.745 ;
        RECT -89.805 -178.240 -88.735 -178.070 ;
        RECT -83.925 -178.070 -83.755 -177.745 ;
        RECT -83.575 -177.845 -83.205 -177.505 ;
        RECT -83.025 -177.745 -82.095 -177.565 ;
        RECT -80.645 -177.745 -79.715 -177.565 ;
        RECT -83.025 -178.070 -82.855 -177.745 ;
        RECT -83.925 -178.240 -82.855 -178.070 ;
        RECT -79.885 -178.070 -79.715 -177.745 ;
        RECT -79.535 -177.845 -79.165 -177.505 ;
        RECT -78.985 -177.745 -78.435 -177.575 ;
        RECT -74.385 -177.745 -73.835 -177.575 ;
        RECT -78.985 -178.070 -78.815 -177.745 ;
        RECT -79.885 -178.240 -78.815 -178.070 ;
        RECT -74.005 -178.070 -73.835 -177.745 ;
        RECT -73.655 -177.845 -73.285 -177.505 ;
        RECT -73.105 -177.745 -72.175 -177.565 ;
        RECT -70.725 -177.745 -69.795 -177.565 ;
        RECT -73.105 -178.070 -72.935 -177.745 ;
        RECT -74.005 -178.240 -72.935 -178.070 ;
        RECT -69.965 -178.070 -69.795 -177.745 ;
        RECT -69.615 -177.845 -69.245 -177.505 ;
        RECT -69.065 -177.745 -68.515 -177.575 ;
        RECT -64.465 -177.745 -63.915 -177.575 ;
        RECT -69.065 -178.070 -68.895 -177.745 ;
        RECT -69.965 -178.240 -68.895 -178.070 ;
        RECT -64.085 -178.070 -63.915 -177.745 ;
        RECT -63.735 -177.845 -63.365 -177.505 ;
        RECT -63.185 -177.745 -62.255 -177.565 ;
        RECT -60.805 -177.745 -59.875 -177.565 ;
        RECT -63.185 -178.070 -63.015 -177.745 ;
        RECT -64.085 -178.240 -63.015 -178.070 ;
        RECT -60.045 -178.070 -59.875 -177.745 ;
        RECT -59.695 -177.845 -59.325 -177.505 ;
        RECT -59.145 -177.745 -58.595 -177.575 ;
        RECT -54.545 -177.745 -53.995 -177.575 ;
        RECT -59.145 -178.070 -58.975 -177.745 ;
        RECT -60.045 -178.240 -58.975 -178.070 ;
        RECT -54.165 -178.070 -53.995 -177.745 ;
        RECT -53.815 -177.845 -53.445 -177.505 ;
        RECT -53.265 -177.745 -52.335 -177.565 ;
        RECT -50.885 -177.745 -49.955 -177.565 ;
        RECT -53.265 -178.070 -53.095 -177.745 ;
        RECT -54.165 -178.240 -53.095 -178.070 ;
        RECT -50.125 -178.070 -49.955 -177.745 ;
        RECT -49.775 -177.845 -49.405 -177.505 ;
        RECT -49.225 -177.745 -48.675 -177.575 ;
        RECT -44.625 -177.745 -44.075 -177.575 ;
        RECT -49.225 -178.070 -49.055 -177.745 ;
        RECT -50.125 -178.240 -49.055 -178.070 ;
        RECT -44.245 -178.070 -44.075 -177.745 ;
        RECT -43.895 -177.845 -43.525 -177.505 ;
        RECT -43.345 -177.745 -42.415 -177.565 ;
        RECT -40.965 -177.745 -40.035 -177.565 ;
        RECT -43.345 -178.070 -43.175 -177.745 ;
        RECT -44.245 -178.240 -43.175 -178.070 ;
        RECT -40.205 -178.070 -40.035 -177.745 ;
        RECT -39.855 -177.845 -39.485 -177.505 ;
        RECT -39.305 -177.745 -38.755 -177.575 ;
        RECT -34.705 -177.745 -34.155 -177.575 ;
        RECT -39.305 -178.070 -39.135 -177.745 ;
        RECT -40.205 -178.240 -39.135 -178.070 ;
        RECT -34.325 -178.070 -34.155 -177.745 ;
        RECT -33.975 -177.845 -33.605 -177.505 ;
        RECT -33.425 -177.745 -32.495 -177.565 ;
        RECT -31.045 -177.745 -30.115 -177.565 ;
        RECT -33.425 -178.070 -33.255 -177.745 ;
        RECT -34.325 -178.240 -33.255 -178.070 ;
        RECT -30.285 -178.070 -30.115 -177.745 ;
        RECT -29.935 -177.845 -29.565 -177.505 ;
        RECT -29.385 -177.745 -28.835 -177.575 ;
        RECT -24.785 -177.745 -24.235 -177.575 ;
        RECT -29.385 -178.070 -29.215 -177.745 ;
        RECT -30.285 -178.240 -29.215 -178.070 ;
        RECT -24.405 -178.070 -24.235 -177.745 ;
        RECT -24.055 -177.845 -23.685 -177.505 ;
        RECT -23.505 -177.745 -22.575 -177.565 ;
        RECT -21.125 -177.745 -20.195 -177.565 ;
        RECT -23.505 -178.070 -23.335 -177.745 ;
        RECT -24.405 -178.240 -23.335 -178.070 ;
        RECT -20.365 -178.070 -20.195 -177.745 ;
        RECT -20.015 -177.845 -19.645 -177.505 ;
        RECT -19.465 -177.745 -18.915 -177.575 ;
        RECT -14.865 -177.745 -14.315 -177.575 ;
        RECT -19.465 -178.070 -19.295 -177.745 ;
        RECT -20.365 -178.240 -19.295 -178.070 ;
        RECT -14.485 -178.070 -14.315 -177.745 ;
        RECT -14.135 -177.845 -13.765 -177.505 ;
        RECT -13.585 -177.745 -12.655 -177.565 ;
        RECT -11.205 -177.745 -10.275 -177.565 ;
        RECT -13.585 -178.070 -13.415 -177.745 ;
        RECT -14.485 -178.240 -13.415 -178.070 ;
        RECT -10.445 -178.070 -10.275 -177.745 ;
        RECT -10.095 -177.845 -9.725 -177.505 ;
        RECT -9.545 -177.745 -8.995 -177.575 ;
        RECT -4.945 -177.745 -4.395 -177.575 ;
        RECT -9.545 -178.070 -9.375 -177.745 ;
        RECT -10.445 -178.240 -9.375 -178.070 ;
        RECT -4.565 -178.070 -4.395 -177.745 ;
        RECT -4.215 -177.845 -3.845 -177.505 ;
        RECT -3.665 -177.745 -2.735 -177.565 ;
        RECT -1.285 -177.745 -0.355 -177.565 ;
        RECT -3.665 -178.070 -3.495 -177.745 ;
        RECT -4.565 -178.240 -3.495 -178.070 ;
        RECT -0.525 -178.070 -0.355 -177.745 ;
        RECT -0.175 -177.845 0.195 -177.505 ;
        RECT 0.375 -177.745 0.925 -177.575 ;
        RECT 4.975 -177.745 5.525 -177.575 ;
        RECT 0.375 -178.070 0.545 -177.745 ;
        RECT -0.525 -178.240 0.545 -178.070 ;
        RECT 5.355 -178.070 5.525 -177.745 ;
        RECT 5.705 -177.845 6.075 -177.505 ;
        RECT 6.255 -177.745 7.185 -177.565 ;
        RECT 8.635 -177.745 9.565 -177.565 ;
        RECT 6.255 -178.070 6.425 -177.745 ;
        RECT 5.355 -178.240 6.425 -178.070 ;
        RECT 9.395 -178.070 9.565 -177.745 ;
        RECT 9.745 -177.845 10.115 -177.505 ;
        RECT 10.295 -177.745 10.845 -177.575 ;
        RECT 14.895 -177.745 15.445 -177.575 ;
        RECT 10.295 -178.070 10.465 -177.745 ;
        RECT 9.395 -178.240 10.465 -178.070 ;
        RECT 15.275 -178.070 15.445 -177.745 ;
        RECT 15.625 -177.845 15.995 -177.505 ;
        RECT 16.175 -177.745 17.105 -177.565 ;
        RECT 18.555 -177.745 19.485 -177.565 ;
        RECT 16.175 -178.070 16.345 -177.745 ;
        RECT 15.275 -178.240 16.345 -178.070 ;
        RECT 19.315 -178.070 19.485 -177.745 ;
        RECT 19.665 -177.845 20.035 -177.505 ;
        RECT 20.215 -177.745 20.765 -177.575 ;
        RECT 20.215 -178.070 20.385 -177.745 ;
        RECT 20.935 -177.925 21.105 -177.400 ;
        RECT 19.315 -178.240 20.385 -178.070 ;
        RECT -292.965 -178.440 -292.795 -178.255 ;
        RECT -291.820 -178.345 -291.490 -178.240 ;
        RECT -287.890 -178.345 -287.560 -178.240 ;
        RECT -281.900 -178.345 -281.570 -178.240 ;
        RECT -277.970 -178.345 -277.640 -178.240 ;
        RECT -271.980 -178.345 -271.650 -178.240 ;
        RECT -268.050 -178.345 -267.720 -178.240 ;
        RECT -262.060 -178.345 -261.730 -178.240 ;
        RECT -258.130 -178.345 -257.800 -178.240 ;
        RECT -252.140 -178.345 -251.810 -178.240 ;
        RECT -248.210 -178.345 -247.880 -178.240 ;
        RECT -242.220 -178.345 -241.890 -178.240 ;
        RECT -238.290 -178.345 -237.960 -178.240 ;
        RECT -232.300 -178.345 -231.970 -178.240 ;
        RECT -228.370 -178.345 -228.040 -178.240 ;
        RECT -222.380 -178.345 -222.050 -178.240 ;
        RECT -218.450 -178.345 -218.120 -178.240 ;
        RECT -212.460 -178.345 -212.130 -178.240 ;
        RECT -208.530 -178.345 -208.200 -178.240 ;
        RECT -202.540 -178.345 -202.210 -178.240 ;
        RECT -198.610 -178.345 -198.280 -178.240 ;
        RECT -192.620 -178.345 -192.290 -178.240 ;
        RECT -188.690 -178.345 -188.360 -178.240 ;
        RECT -182.700 -178.345 -182.370 -178.240 ;
        RECT -178.770 -178.345 -178.440 -178.240 ;
        RECT -172.780 -178.345 -172.450 -178.240 ;
        RECT -168.850 -178.345 -168.520 -178.240 ;
        RECT -162.860 -178.345 -162.530 -178.240 ;
        RECT -158.930 -178.345 -158.600 -178.240 ;
        RECT -152.940 -178.345 -152.610 -178.240 ;
        RECT -149.010 -178.345 -148.680 -178.240 ;
        RECT -143.020 -178.345 -142.690 -178.240 ;
        RECT -139.090 -178.345 -138.760 -178.240 ;
        RECT -133.100 -178.345 -132.770 -178.240 ;
        RECT -129.170 -178.345 -128.840 -178.240 ;
        RECT -123.180 -178.345 -122.850 -178.240 ;
        RECT -119.250 -178.345 -118.920 -178.240 ;
        RECT -113.260 -178.345 -112.930 -178.240 ;
        RECT -109.330 -178.345 -109.000 -178.240 ;
        RECT -103.340 -178.345 -103.010 -178.240 ;
        RECT -99.410 -178.345 -99.080 -178.240 ;
        RECT -93.420 -178.345 -93.090 -178.240 ;
        RECT -89.490 -178.345 -89.160 -178.240 ;
        RECT -83.500 -178.345 -83.170 -178.240 ;
        RECT -79.570 -178.345 -79.240 -178.240 ;
        RECT -73.580 -178.345 -73.250 -178.240 ;
        RECT -69.650 -178.345 -69.320 -178.240 ;
        RECT -63.660 -178.345 -63.330 -178.240 ;
        RECT -59.730 -178.345 -59.400 -178.240 ;
        RECT -53.740 -178.345 -53.410 -178.240 ;
        RECT -49.810 -178.345 -49.480 -178.240 ;
        RECT -43.820 -178.345 -43.490 -178.240 ;
        RECT -39.890 -178.345 -39.560 -178.240 ;
        RECT -33.900 -178.345 -33.570 -178.240 ;
        RECT -29.970 -178.345 -29.640 -178.240 ;
        RECT -23.980 -178.345 -23.650 -178.240 ;
        RECT -20.050 -178.345 -19.720 -178.240 ;
        RECT -14.060 -178.345 -13.730 -178.240 ;
        RECT -10.130 -178.345 -9.800 -178.240 ;
        RECT -4.140 -178.345 -3.810 -178.240 ;
        RECT -0.210 -178.345 0.120 -178.240 ;
        RECT 5.780 -178.345 6.110 -178.240 ;
        RECT 9.710 -178.345 10.040 -178.240 ;
        RECT 15.700 -178.345 16.030 -178.240 ;
        RECT 19.630 -178.345 19.960 -178.240 ;
        RECT 20.555 -178.255 21.105 -177.925 ;
        RECT -293.495 -178.455 -292.795 -178.440 ;
        RECT -293.580 -178.625 -292.795 -178.455 ;
        RECT -293.260 -178.630 -292.795 -178.625 ;
        RECT -292.965 -178.780 -292.795 -178.630 ;
        RECT -288.965 -178.515 -288.060 -178.425 ;
        RECT -287.260 -178.515 -286.755 -178.435 ;
        RECT -288.965 -178.695 -286.755 -178.515 ;
        RECT -279.045 -178.515 -278.140 -178.425 ;
        RECT -277.340 -178.515 -276.835 -178.435 ;
        RECT -279.045 -178.695 -276.835 -178.515 ;
        RECT -269.125 -178.515 -268.220 -178.425 ;
        RECT -267.420 -178.515 -266.915 -178.435 ;
        RECT -269.125 -178.695 -266.915 -178.515 ;
        RECT -259.205 -178.515 -258.300 -178.425 ;
        RECT -257.500 -178.515 -256.995 -178.435 ;
        RECT -259.205 -178.695 -256.995 -178.515 ;
        RECT -249.285 -178.515 -248.380 -178.425 ;
        RECT -247.580 -178.515 -247.075 -178.435 ;
        RECT -249.285 -178.695 -247.075 -178.515 ;
        RECT -239.365 -178.515 -238.460 -178.425 ;
        RECT -237.660 -178.515 -237.155 -178.435 ;
        RECT -239.365 -178.695 -237.155 -178.515 ;
        RECT -229.445 -178.515 -228.540 -178.425 ;
        RECT -227.740 -178.515 -227.235 -178.435 ;
        RECT -229.445 -178.695 -227.235 -178.515 ;
        RECT -219.525 -178.515 -218.620 -178.425 ;
        RECT -217.820 -178.515 -217.315 -178.435 ;
        RECT -219.525 -178.695 -217.315 -178.515 ;
        RECT -209.605 -178.515 -208.700 -178.425 ;
        RECT -207.900 -178.515 -207.395 -178.435 ;
        RECT -209.605 -178.695 -207.395 -178.515 ;
        RECT -199.685 -178.515 -198.780 -178.425 ;
        RECT -197.980 -178.515 -197.475 -178.435 ;
        RECT -199.685 -178.695 -197.475 -178.515 ;
        RECT -189.765 -178.515 -188.860 -178.425 ;
        RECT -188.060 -178.515 -187.555 -178.435 ;
        RECT -189.765 -178.695 -187.555 -178.515 ;
        RECT -179.845 -178.515 -178.940 -178.425 ;
        RECT -178.140 -178.515 -177.635 -178.435 ;
        RECT -179.845 -178.695 -177.635 -178.515 ;
        RECT -169.925 -178.515 -169.020 -178.425 ;
        RECT -168.220 -178.515 -167.715 -178.435 ;
        RECT -169.925 -178.695 -167.715 -178.515 ;
        RECT -160.005 -178.515 -159.100 -178.425 ;
        RECT -158.300 -178.515 -157.795 -178.435 ;
        RECT -160.005 -178.695 -157.795 -178.515 ;
        RECT -150.085 -178.515 -149.180 -178.425 ;
        RECT -148.380 -178.515 -147.875 -178.435 ;
        RECT -150.085 -178.695 -147.875 -178.515 ;
        RECT -140.165 -178.515 -139.260 -178.425 ;
        RECT -138.460 -178.515 -137.955 -178.435 ;
        RECT -140.165 -178.695 -137.955 -178.515 ;
        RECT -130.245 -178.515 -129.340 -178.425 ;
        RECT -128.540 -178.515 -128.035 -178.435 ;
        RECT -130.245 -178.695 -128.035 -178.515 ;
        RECT -120.325 -178.515 -119.420 -178.425 ;
        RECT -118.620 -178.515 -118.115 -178.435 ;
        RECT -120.325 -178.695 -118.115 -178.515 ;
        RECT -110.405 -178.515 -109.500 -178.425 ;
        RECT -108.700 -178.515 -108.195 -178.435 ;
        RECT -110.405 -178.695 -108.195 -178.515 ;
        RECT -100.485 -178.515 -99.580 -178.425 ;
        RECT -98.780 -178.515 -98.275 -178.435 ;
        RECT -100.485 -178.695 -98.275 -178.515 ;
        RECT -90.565 -178.515 -89.660 -178.425 ;
        RECT -88.860 -178.515 -88.355 -178.435 ;
        RECT -90.565 -178.695 -88.355 -178.515 ;
        RECT -80.645 -178.515 -79.740 -178.425 ;
        RECT -78.940 -178.515 -78.435 -178.435 ;
        RECT -80.645 -178.695 -78.435 -178.515 ;
        RECT -70.725 -178.515 -69.820 -178.425 ;
        RECT -69.020 -178.515 -68.515 -178.435 ;
        RECT -70.725 -178.695 -68.515 -178.515 ;
        RECT -60.805 -178.515 -59.900 -178.425 ;
        RECT -59.100 -178.515 -58.595 -178.435 ;
        RECT -60.805 -178.695 -58.595 -178.515 ;
        RECT -50.885 -178.515 -49.980 -178.425 ;
        RECT -49.180 -178.515 -48.675 -178.435 ;
        RECT -50.885 -178.695 -48.675 -178.515 ;
        RECT -40.965 -178.515 -40.060 -178.425 ;
        RECT -39.260 -178.515 -38.755 -178.435 ;
        RECT -40.965 -178.695 -38.755 -178.515 ;
        RECT -31.045 -178.515 -30.140 -178.425 ;
        RECT -29.340 -178.515 -28.835 -178.435 ;
        RECT -31.045 -178.695 -28.835 -178.515 ;
        RECT -21.125 -178.515 -20.220 -178.425 ;
        RECT -19.420 -178.515 -18.915 -178.435 ;
        RECT -21.125 -178.695 -18.915 -178.515 ;
        RECT -11.205 -178.515 -10.300 -178.425 ;
        RECT -9.500 -178.515 -8.995 -178.435 ;
        RECT -11.205 -178.695 -8.995 -178.515 ;
        RECT -1.285 -178.515 -0.380 -178.425 ;
        RECT 0.420 -178.515 0.925 -178.435 ;
        RECT -1.285 -178.695 0.925 -178.515 ;
        RECT 8.635 -178.515 9.540 -178.425 ;
        RECT 10.340 -178.515 10.845 -178.435 ;
        RECT 8.635 -178.695 10.845 -178.515 ;
        RECT 18.555 -178.515 19.460 -178.425 ;
        RECT 20.260 -178.515 20.765 -178.435 ;
        RECT 18.555 -178.695 20.765 -178.515 ;
        RECT 20.935 -178.450 21.105 -178.255 ;
        RECT 21.345 -178.450 21.635 -177.730 ;
        RECT 20.935 -178.455 21.635 -178.450 ;
        RECT 20.935 -178.625 21.720 -178.455 ;
        RECT 20.935 -178.630 21.400 -178.625 ;
        RECT 20.935 -178.780 21.105 -178.630 ;
      LAYER mcon ;
        RECT -291.315 94.820 -291.145 94.990 ;
        RECT -290.845 94.825 -290.675 94.995 ;
        RECT -290.020 94.795 -289.850 94.965 ;
        RECT -288.655 94.795 -288.485 94.965 ;
        RECT -280.100 94.795 -279.930 94.965 ;
        RECT -278.735 94.795 -278.565 94.965 ;
        RECT -270.180 94.795 -270.010 94.965 ;
        RECT -268.815 94.795 -268.645 94.965 ;
        RECT -260.260 94.795 -260.090 94.965 ;
        RECT -258.895 94.795 -258.725 94.965 ;
        RECT -250.340 94.795 -250.170 94.965 ;
        RECT -248.975 94.795 -248.805 94.965 ;
        RECT -240.420 94.795 -240.250 94.965 ;
        RECT -239.055 94.795 -238.885 94.965 ;
        RECT -230.500 94.795 -230.330 94.965 ;
        RECT -229.135 94.795 -228.965 94.965 ;
        RECT -220.580 94.795 -220.410 94.965 ;
        RECT -219.215 94.795 -219.045 94.965 ;
        RECT -210.660 94.795 -210.490 94.965 ;
        RECT -209.295 94.795 -209.125 94.965 ;
        RECT -200.740 94.795 -200.570 94.965 ;
        RECT -199.375 94.795 -199.205 94.965 ;
        RECT -190.820 94.795 -190.650 94.965 ;
        RECT -189.455 94.795 -189.285 94.965 ;
        RECT -180.900 94.795 -180.730 94.965 ;
        RECT -179.535 94.795 -179.365 94.965 ;
        RECT -170.980 94.795 -170.810 94.965 ;
        RECT -169.615 94.795 -169.445 94.965 ;
        RECT -161.060 94.795 -160.890 94.965 ;
        RECT -159.695 94.795 -159.525 94.965 ;
        RECT -151.140 94.795 -150.970 94.965 ;
        RECT -149.775 94.795 -149.605 94.965 ;
        RECT -141.220 94.795 -141.050 94.965 ;
        RECT -139.855 94.795 -139.685 94.965 ;
        RECT -131.300 94.795 -131.130 94.965 ;
        RECT -129.935 94.795 -129.765 94.965 ;
        RECT -121.380 94.795 -121.210 94.965 ;
        RECT -120.015 94.795 -119.845 94.965 ;
        RECT -111.460 94.795 -111.290 94.965 ;
        RECT -110.095 94.795 -109.925 94.965 ;
        RECT -101.540 94.795 -101.370 94.965 ;
        RECT -100.175 94.795 -100.005 94.965 ;
        RECT -91.620 94.795 -91.450 94.965 ;
        RECT -90.255 94.795 -90.085 94.965 ;
        RECT -81.700 94.795 -81.530 94.965 ;
        RECT -80.335 94.795 -80.165 94.965 ;
        RECT -71.780 94.795 -71.610 94.965 ;
        RECT -70.415 94.795 -70.245 94.965 ;
        RECT -61.860 94.795 -61.690 94.965 ;
        RECT -60.495 94.795 -60.325 94.965 ;
        RECT -51.940 94.795 -51.770 94.965 ;
        RECT -50.575 94.795 -50.405 94.965 ;
        RECT -42.020 94.795 -41.850 94.965 ;
        RECT -40.655 94.795 -40.485 94.965 ;
        RECT -32.100 94.795 -31.930 94.965 ;
        RECT -30.735 94.795 -30.565 94.965 ;
        RECT -22.180 94.795 -22.010 94.965 ;
        RECT -20.815 94.795 -20.645 94.965 ;
        RECT -12.260 94.795 -12.090 94.965 ;
        RECT -10.895 94.795 -10.725 94.965 ;
        RECT -2.340 94.795 -2.170 94.965 ;
        RECT -0.975 94.795 -0.805 94.965 ;
        RECT 7.580 94.795 7.750 94.965 ;
        RECT 8.945 94.795 9.115 94.965 ;
        RECT 17.500 94.795 17.670 94.965 ;
        RECT 18.865 94.795 19.035 94.965 ;
        RECT -290.845 94.365 -290.675 94.535 ;
        RECT -290.845 93.905 -290.675 94.075 ;
        RECT -289.285 93.945 -289.115 94.115 ;
        RECT -283.425 93.945 -283.255 94.115 ;
        RECT -279.365 93.945 -279.195 94.115 ;
        RECT -273.505 93.945 -273.335 94.115 ;
        RECT -269.445 93.945 -269.275 94.115 ;
        RECT -263.585 93.945 -263.415 94.115 ;
        RECT -259.525 93.945 -259.355 94.115 ;
        RECT -253.665 93.945 -253.495 94.115 ;
        RECT -249.605 93.945 -249.435 94.115 ;
        RECT -243.745 93.945 -243.575 94.115 ;
        RECT -239.685 93.945 -239.515 94.115 ;
        RECT -233.825 93.945 -233.655 94.115 ;
        RECT -229.765 93.945 -229.595 94.115 ;
        RECT -223.905 93.945 -223.735 94.115 ;
        RECT -219.845 93.945 -219.675 94.115 ;
        RECT -213.985 93.945 -213.815 94.115 ;
        RECT -209.925 93.945 -209.755 94.115 ;
        RECT -204.065 93.945 -203.895 94.115 ;
        RECT -200.005 93.945 -199.835 94.115 ;
        RECT -194.145 93.945 -193.975 94.115 ;
        RECT -190.085 93.945 -189.915 94.115 ;
        RECT -184.225 93.945 -184.055 94.115 ;
        RECT -180.165 93.945 -179.995 94.115 ;
        RECT -174.305 93.945 -174.135 94.115 ;
        RECT -170.245 93.945 -170.075 94.115 ;
        RECT -164.385 93.945 -164.215 94.115 ;
        RECT -160.325 93.945 -160.155 94.115 ;
        RECT -154.465 93.945 -154.295 94.115 ;
        RECT -150.405 93.945 -150.235 94.115 ;
        RECT -144.545 93.945 -144.375 94.115 ;
        RECT -140.485 93.945 -140.315 94.115 ;
        RECT -134.625 93.945 -134.455 94.115 ;
        RECT -130.565 93.945 -130.395 94.115 ;
        RECT -124.705 93.945 -124.535 94.115 ;
        RECT -120.645 93.945 -120.475 94.115 ;
        RECT -114.785 93.945 -114.615 94.115 ;
        RECT -110.725 93.945 -110.555 94.115 ;
        RECT -104.865 93.945 -104.695 94.115 ;
        RECT -100.805 93.945 -100.635 94.115 ;
        RECT -94.945 93.945 -94.775 94.115 ;
        RECT -90.885 93.945 -90.715 94.115 ;
        RECT -85.025 93.945 -84.855 94.115 ;
        RECT -80.965 93.945 -80.795 94.115 ;
        RECT -75.105 93.945 -74.935 94.115 ;
        RECT -71.045 93.945 -70.875 94.115 ;
        RECT -65.185 93.945 -65.015 94.115 ;
        RECT -61.125 93.945 -60.955 94.115 ;
        RECT -55.265 93.945 -55.095 94.115 ;
        RECT -51.205 93.945 -51.035 94.115 ;
        RECT -45.345 93.945 -45.175 94.115 ;
        RECT -41.285 93.945 -41.115 94.115 ;
        RECT -35.425 93.945 -35.255 94.115 ;
        RECT -31.365 93.945 -31.195 94.115 ;
        RECT -25.505 93.945 -25.335 94.115 ;
        RECT -21.445 93.945 -21.275 94.115 ;
        RECT -15.585 93.945 -15.415 94.115 ;
        RECT -11.525 93.945 -11.355 94.115 ;
        RECT -5.665 93.945 -5.495 94.115 ;
        RECT -1.605 93.945 -1.435 94.115 ;
        RECT 4.255 93.945 4.425 94.115 ;
        RECT 8.315 93.945 8.485 94.115 ;
        RECT 14.175 93.945 14.345 94.115 ;
        RECT 18.235 93.945 18.405 94.115 ;
        RECT 24.095 93.945 24.265 94.115 ;
        RECT -291.315 93.245 -291.145 93.415 ;
        RECT -290.855 93.245 -290.685 93.415 ;
        RECT -290.395 93.245 -290.225 93.415 ;
        RECT -289.935 93.245 -289.765 93.415 ;
        RECT 24.745 93.245 24.915 93.415 ;
        RECT 25.205 93.245 25.375 93.415 ;
        RECT 25.665 93.245 25.835 93.415 ;
        RECT 26.125 93.245 26.295 93.415 ;
        RECT -289.965 92.525 -289.795 92.695 ;
        RECT -289.980 92.085 -289.810 92.255 ;
        RECT -282.745 92.525 -282.575 92.695 ;
        RECT -287.690 91.685 -287.520 91.855 ;
        RECT -287.705 91.245 -287.535 91.415 ;
        RECT -282.730 92.085 -282.560 92.255 ;
        RECT -285.020 91.685 -284.850 91.855 ;
        RECT -280.045 92.525 -279.875 92.695 ;
        RECT -280.060 92.085 -279.890 92.255 ;
        RECT -272.825 92.525 -272.655 92.695 ;
        RECT -285.005 91.245 -284.835 91.415 ;
        RECT -277.770 91.685 -277.600 91.855 ;
        RECT -277.785 91.245 -277.615 91.415 ;
        RECT -272.810 92.085 -272.640 92.255 ;
        RECT -275.100 91.685 -274.930 91.855 ;
        RECT -270.125 92.525 -269.955 92.695 ;
        RECT -270.140 92.085 -269.970 92.255 ;
        RECT -262.905 92.525 -262.735 92.695 ;
        RECT -275.085 91.245 -274.915 91.415 ;
        RECT -267.850 91.685 -267.680 91.855 ;
        RECT -267.865 91.245 -267.695 91.415 ;
        RECT -262.890 92.085 -262.720 92.255 ;
        RECT -265.180 91.685 -265.010 91.855 ;
        RECT -260.205 92.525 -260.035 92.695 ;
        RECT -260.220 92.085 -260.050 92.255 ;
        RECT -252.985 92.525 -252.815 92.695 ;
        RECT -265.165 91.245 -264.995 91.415 ;
        RECT -257.930 91.685 -257.760 91.855 ;
        RECT -257.945 91.245 -257.775 91.415 ;
        RECT -252.970 92.085 -252.800 92.255 ;
        RECT -255.260 91.685 -255.090 91.855 ;
        RECT -250.285 92.525 -250.115 92.695 ;
        RECT -250.300 92.085 -250.130 92.255 ;
        RECT -243.065 92.525 -242.895 92.695 ;
        RECT -255.245 91.245 -255.075 91.415 ;
        RECT -248.010 91.685 -247.840 91.855 ;
        RECT -248.025 91.245 -247.855 91.415 ;
        RECT -243.050 92.085 -242.880 92.255 ;
        RECT -245.340 91.685 -245.170 91.855 ;
        RECT -240.365 92.525 -240.195 92.695 ;
        RECT -240.380 92.085 -240.210 92.255 ;
        RECT -233.145 92.525 -232.975 92.695 ;
        RECT -245.325 91.245 -245.155 91.415 ;
        RECT -238.090 91.685 -237.920 91.855 ;
        RECT -238.105 91.245 -237.935 91.415 ;
        RECT -233.130 92.085 -232.960 92.255 ;
        RECT -235.420 91.685 -235.250 91.855 ;
        RECT -230.445 92.525 -230.275 92.695 ;
        RECT -230.460 92.085 -230.290 92.255 ;
        RECT -223.225 92.525 -223.055 92.695 ;
        RECT -235.405 91.245 -235.235 91.415 ;
        RECT -228.170 91.685 -228.000 91.855 ;
        RECT -228.185 91.245 -228.015 91.415 ;
        RECT -223.210 92.085 -223.040 92.255 ;
        RECT -225.500 91.685 -225.330 91.855 ;
        RECT -220.525 92.525 -220.355 92.695 ;
        RECT -220.540 92.085 -220.370 92.255 ;
        RECT -213.305 92.525 -213.135 92.695 ;
        RECT -225.485 91.245 -225.315 91.415 ;
        RECT -218.250 91.685 -218.080 91.855 ;
        RECT -218.265 91.245 -218.095 91.415 ;
        RECT -213.290 92.085 -213.120 92.255 ;
        RECT -215.580 91.685 -215.410 91.855 ;
        RECT -210.605 92.525 -210.435 92.695 ;
        RECT -210.620 92.085 -210.450 92.255 ;
        RECT -203.385 92.525 -203.215 92.695 ;
        RECT -215.565 91.245 -215.395 91.415 ;
        RECT -208.330 91.685 -208.160 91.855 ;
        RECT -208.345 91.245 -208.175 91.415 ;
        RECT -203.370 92.085 -203.200 92.255 ;
        RECT -205.660 91.685 -205.490 91.855 ;
        RECT -200.685 92.525 -200.515 92.695 ;
        RECT -200.700 92.085 -200.530 92.255 ;
        RECT -193.465 92.525 -193.295 92.695 ;
        RECT -205.645 91.245 -205.475 91.415 ;
        RECT -198.410 91.685 -198.240 91.855 ;
        RECT -198.425 91.245 -198.255 91.415 ;
        RECT -193.450 92.085 -193.280 92.255 ;
        RECT -195.740 91.685 -195.570 91.855 ;
        RECT -190.765 92.525 -190.595 92.695 ;
        RECT -190.780 92.085 -190.610 92.255 ;
        RECT -183.545 92.525 -183.375 92.695 ;
        RECT -195.725 91.245 -195.555 91.415 ;
        RECT -188.490 91.685 -188.320 91.855 ;
        RECT -188.505 91.245 -188.335 91.415 ;
        RECT -183.530 92.085 -183.360 92.255 ;
        RECT -185.820 91.685 -185.650 91.855 ;
        RECT -180.845 92.525 -180.675 92.695 ;
        RECT -180.860 92.085 -180.690 92.255 ;
        RECT -173.625 92.525 -173.455 92.695 ;
        RECT -185.805 91.245 -185.635 91.415 ;
        RECT -178.570 91.685 -178.400 91.855 ;
        RECT -178.585 91.245 -178.415 91.415 ;
        RECT -173.610 92.085 -173.440 92.255 ;
        RECT -175.900 91.685 -175.730 91.855 ;
        RECT -170.925 92.525 -170.755 92.695 ;
        RECT -170.940 92.085 -170.770 92.255 ;
        RECT -163.705 92.525 -163.535 92.695 ;
        RECT -175.885 91.245 -175.715 91.415 ;
        RECT -168.650 91.685 -168.480 91.855 ;
        RECT -168.665 91.245 -168.495 91.415 ;
        RECT -163.690 92.085 -163.520 92.255 ;
        RECT -165.980 91.685 -165.810 91.855 ;
        RECT -161.005 92.525 -160.835 92.695 ;
        RECT -161.020 92.085 -160.850 92.255 ;
        RECT -153.785 92.525 -153.615 92.695 ;
        RECT -165.965 91.245 -165.795 91.415 ;
        RECT -158.730 91.685 -158.560 91.855 ;
        RECT -158.745 91.245 -158.575 91.415 ;
        RECT -153.770 92.085 -153.600 92.255 ;
        RECT -156.060 91.685 -155.890 91.855 ;
        RECT -151.085 92.525 -150.915 92.695 ;
        RECT -151.100 92.085 -150.930 92.255 ;
        RECT -143.865 92.525 -143.695 92.695 ;
        RECT -156.045 91.245 -155.875 91.415 ;
        RECT -148.810 91.685 -148.640 91.855 ;
        RECT -148.825 91.245 -148.655 91.415 ;
        RECT -143.850 92.085 -143.680 92.255 ;
        RECT -146.140 91.685 -145.970 91.855 ;
        RECT -141.165 92.525 -140.995 92.695 ;
        RECT -141.180 92.085 -141.010 92.255 ;
        RECT -133.945 92.525 -133.775 92.695 ;
        RECT -146.125 91.245 -145.955 91.415 ;
        RECT -138.890 91.685 -138.720 91.855 ;
        RECT -138.905 91.245 -138.735 91.415 ;
        RECT -133.930 92.085 -133.760 92.255 ;
        RECT -136.220 91.685 -136.050 91.855 ;
        RECT -131.245 92.525 -131.075 92.695 ;
        RECT -131.260 92.085 -131.090 92.255 ;
        RECT -124.025 92.525 -123.855 92.695 ;
        RECT -136.205 91.245 -136.035 91.415 ;
        RECT -128.970 91.685 -128.800 91.855 ;
        RECT -128.985 91.245 -128.815 91.415 ;
        RECT -124.010 92.085 -123.840 92.255 ;
        RECT -126.300 91.685 -126.130 91.855 ;
        RECT -121.325 92.525 -121.155 92.695 ;
        RECT -121.340 92.085 -121.170 92.255 ;
        RECT -114.105 92.525 -113.935 92.695 ;
        RECT -126.285 91.245 -126.115 91.415 ;
        RECT -119.050 91.685 -118.880 91.855 ;
        RECT -119.065 91.245 -118.895 91.415 ;
        RECT -114.090 92.085 -113.920 92.255 ;
        RECT -116.380 91.685 -116.210 91.855 ;
        RECT -111.405 92.525 -111.235 92.695 ;
        RECT -111.420 92.085 -111.250 92.255 ;
        RECT -104.185 92.525 -104.015 92.695 ;
        RECT -116.365 91.245 -116.195 91.415 ;
        RECT -109.130 91.685 -108.960 91.855 ;
        RECT -109.145 91.245 -108.975 91.415 ;
        RECT -104.170 92.085 -104.000 92.255 ;
        RECT -106.460 91.685 -106.290 91.855 ;
        RECT -101.485 92.525 -101.315 92.695 ;
        RECT -101.500 92.085 -101.330 92.255 ;
        RECT -94.265 92.525 -94.095 92.695 ;
        RECT -106.445 91.245 -106.275 91.415 ;
        RECT -99.210 91.685 -99.040 91.855 ;
        RECT -99.225 91.245 -99.055 91.415 ;
        RECT -94.250 92.085 -94.080 92.255 ;
        RECT -96.540 91.685 -96.370 91.855 ;
        RECT -91.565 92.525 -91.395 92.695 ;
        RECT -91.580 92.085 -91.410 92.255 ;
        RECT -84.345 92.525 -84.175 92.695 ;
        RECT -96.525 91.245 -96.355 91.415 ;
        RECT -89.290 91.685 -89.120 91.855 ;
        RECT -89.305 91.245 -89.135 91.415 ;
        RECT -84.330 92.085 -84.160 92.255 ;
        RECT -86.620 91.685 -86.450 91.855 ;
        RECT -81.645 92.525 -81.475 92.695 ;
        RECT -81.660 92.085 -81.490 92.255 ;
        RECT -74.425 92.525 -74.255 92.695 ;
        RECT -86.605 91.245 -86.435 91.415 ;
        RECT -79.370 91.685 -79.200 91.855 ;
        RECT -79.385 91.245 -79.215 91.415 ;
        RECT -74.410 92.085 -74.240 92.255 ;
        RECT -76.700 91.685 -76.530 91.855 ;
        RECT -71.725 92.525 -71.555 92.695 ;
        RECT -71.740 92.085 -71.570 92.255 ;
        RECT -64.505 92.525 -64.335 92.695 ;
        RECT -76.685 91.245 -76.515 91.415 ;
        RECT -69.450 91.685 -69.280 91.855 ;
        RECT -69.465 91.245 -69.295 91.415 ;
        RECT -64.490 92.085 -64.320 92.255 ;
        RECT -66.780 91.685 -66.610 91.855 ;
        RECT -61.805 92.525 -61.635 92.695 ;
        RECT -61.820 92.085 -61.650 92.255 ;
        RECT -54.585 92.525 -54.415 92.695 ;
        RECT -66.765 91.245 -66.595 91.415 ;
        RECT -59.530 91.685 -59.360 91.855 ;
        RECT -59.545 91.245 -59.375 91.415 ;
        RECT -54.570 92.085 -54.400 92.255 ;
        RECT -56.860 91.685 -56.690 91.855 ;
        RECT -51.885 92.525 -51.715 92.695 ;
        RECT -51.900 92.085 -51.730 92.255 ;
        RECT -44.665 92.525 -44.495 92.695 ;
        RECT -56.845 91.245 -56.675 91.415 ;
        RECT -49.610 91.685 -49.440 91.855 ;
        RECT -49.625 91.245 -49.455 91.415 ;
        RECT -44.650 92.085 -44.480 92.255 ;
        RECT -46.940 91.685 -46.770 91.855 ;
        RECT -41.965 92.525 -41.795 92.695 ;
        RECT -41.980 92.085 -41.810 92.255 ;
        RECT -34.745 92.525 -34.575 92.695 ;
        RECT -46.925 91.245 -46.755 91.415 ;
        RECT -39.690 91.685 -39.520 91.855 ;
        RECT -39.705 91.245 -39.535 91.415 ;
        RECT -34.730 92.085 -34.560 92.255 ;
        RECT -37.020 91.685 -36.850 91.855 ;
        RECT -32.045 92.525 -31.875 92.695 ;
        RECT -32.060 92.085 -31.890 92.255 ;
        RECT -24.825 92.525 -24.655 92.695 ;
        RECT -37.005 91.245 -36.835 91.415 ;
        RECT -29.770 91.685 -29.600 91.855 ;
        RECT -29.785 91.245 -29.615 91.415 ;
        RECT -24.810 92.085 -24.640 92.255 ;
        RECT -27.100 91.685 -26.930 91.855 ;
        RECT -22.125 92.525 -21.955 92.695 ;
        RECT -22.140 92.085 -21.970 92.255 ;
        RECT -14.905 92.525 -14.735 92.695 ;
        RECT -27.085 91.245 -26.915 91.415 ;
        RECT -19.850 91.685 -19.680 91.855 ;
        RECT -19.865 91.245 -19.695 91.415 ;
        RECT -14.890 92.085 -14.720 92.255 ;
        RECT -17.180 91.685 -17.010 91.855 ;
        RECT -12.205 92.525 -12.035 92.695 ;
        RECT -12.220 92.085 -12.050 92.255 ;
        RECT -4.985 92.525 -4.815 92.695 ;
        RECT -17.165 91.245 -16.995 91.415 ;
        RECT -9.930 91.685 -9.760 91.855 ;
        RECT -9.945 91.245 -9.775 91.415 ;
        RECT -4.970 92.085 -4.800 92.255 ;
        RECT -7.260 91.685 -7.090 91.855 ;
        RECT -2.285 92.525 -2.115 92.695 ;
        RECT -2.300 92.085 -2.130 92.255 ;
        RECT 4.935 92.525 5.105 92.695 ;
        RECT -7.245 91.245 -7.075 91.415 ;
        RECT -0.010 91.685 0.160 91.855 ;
        RECT -0.025 91.245 0.145 91.415 ;
        RECT 4.950 92.085 5.120 92.255 ;
        RECT 2.660 91.685 2.830 91.855 ;
        RECT 7.635 92.525 7.805 92.695 ;
        RECT 7.620 92.085 7.790 92.255 ;
        RECT 14.855 92.525 15.025 92.695 ;
        RECT 2.675 91.245 2.845 91.415 ;
        RECT 9.910 91.685 10.080 91.855 ;
        RECT 9.895 91.245 10.065 91.415 ;
        RECT 14.870 92.085 15.040 92.255 ;
        RECT 12.580 91.685 12.750 91.855 ;
        RECT 17.555 92.525 17.725 92.695 ;
        RECT 17.540 92.085 17.710 92.255 ;
        RECT 24.775 92.525 24.945 92.695 ;
        RECT 12.595 91.245 12.765 91.415 ;
        RECT 19.830 91.685 20.000 91.855 ;
        RECT 19.815 91.245 19.985 91.415 ;
        RECT 24.790 92.085 24.960 92.255 ;
        RECT 22.500 91.685 22.670 91.855 ;
        RECT 22.515 91.245 22.685 91.415 ;
        RECT -291.315 90.525 -291.145 90.695 ;
        RECT -290.855 90.525 -290.685 90.695 ;
        RECT -290.395 90.525 -290.225 90.695 ;
        RECT -289.935 90.525 -289.765 90.695 ;
        RECT -289.545 89.865 -289.375 90.035 ;
        RECT -289.545 89.405 -289.375 89.575 ;
        RECT -288.385 89.825 -288.215 89.995 ;
        RECT -284.325 89.825 -284.155 89.995 ;
        RECT -278.465 89.825 -278.295 89.995 ;
        RECT -274.405 89.825 -274.235 89.995 ;
        RECT -268.545 89.825 -268.375 89.995 ;
        RECT -264.485 89.825 -264.315 89.995 ;
        RECT -258.625 89.825 -258.455 89.995 ;
        RECT -254.565 89.825 -254.395 89.995 ;
        RECT -248.705 89.825 -248.535 89.995 ;
        RECT -244.645 89.825 -244.475 89.995 ;
        RECT -238.785 89.825 -238.615 89.995 ;
        RECT -234.725 89.825 -234.555 89.995 ;
        RECT -228.865 89.825 -228.695 89.995 ;
        RECT -224.805 89.825 -224.635 89.995 ;
        RECT -218.945 89.825 -218.775 89.995 ;
        RECT -214.885 89.825 -214.715 89.995 ;
        RECT -209.025 89.825 -208.855 89.995 ;
        RECT -204.965 89.825 -204.795 89.995 ;
        RECT -199.105 89.825 -198.935 89.995 ;
        RECT -195.045 89.825 -194.875 89.995 ;
        RECT -189.185 89.825 -189.015 89.995 ;
        RECT -185.125 89.825 -184.955 89.995 ;
        RECT -179.265 89.825 -179.095 89.995 ;
        RECT -175.205 89.825 -175.035 89.995 ;
        RECT -169.345 89.825 -169.175 89.995 ;
        RECT -165.285 89.825 -165.115 89.995 ;
        RECT -159.425 89.825 -159.255 89.995 ;
        RECT -155.365 89.825 -155.195 89.995 ;
        RECT -149.505 89.825 -149.335 89.995 ;
        RECT -145.445 89.825 -145.275 89.995 ;
        RECT -139.585 89.825 -139.415 89.995 ;
        RECT -135.525 89.825 -135.355 89.995 ;
        RECT -129.665 89.825 -129.495 89.995 ;
        RECT -125.605 89.825 -125.435 89.995 ;
        RECT -119.745 89.825 -119.575 89.995 ;
        RECT -115.685 89.825 -115.515 89.995 ;
        RECT -109.825 89.825 -109.655 89.995 ;
        RECT -105.765 89.825 -105.595 89.995 ;
        RECT -99.905 89.825 -99.735 89.995 ;
        RECT -95.845 89.825 -95.675 89.995 ;
        RECT -89.985 89.825 -89.815 89.995 ;
        RECT -85.925 89.825 -85.755 89.995 ;
        RECT -80.065 89.825 -79.895 89.995 ;
        RECT -76.005 89.825 -75.835 89.995 ;
        RECT -70.145 89.825 -69.975 89.995 ;
        RECT -66.085 89.825 -65.915 89.995 ;
        RECT -60.225 89.825 -60.055 89.995 ;
        RECT -56.165 89.825 -55.995 89.995 ;
        RECT -50.305 89.825 -50.135 89.995 ;
        RECT -46.245 89.825 -46.075 89.995 ;
        RECT -40.385 89.825 -40.215 89.995 ;
        RECT -36.325 89.825 -36.155 89.995 ;
        RECT -30.465 89.825 -30.295 89.995 ;
        RECT -26.405 89.825 -26.235 89.995 ;
        RECT -20.545 89.825 -20.375 89.995 ;
        RECT -16.485 89.825 -16.315 89.995 ;
        RECT -10.625 89.825 -10.455 89.995 ;
        RECT -6.565 89.825 -6.395 89.995 ;
        RECT -0.705 89.825 -0.535 89.995 ;
        RECT 3.355 89.825 3.525 89.995 ;
        RECT 9.215 89.825 9.385 89.995 ;
        RECT 13.275 89.825 13.445 89.995 ;
        RECT 19.135 89.825 19.305 89.995 ;
        RECT 23.195 89.825 23.365 89.995 ;
        RECT 24.355 89.865 24.525 90.035 ;
        RECT 24.355 89.405 24.525 89.575 ;
        RECT -290.015 88.955 -289.845 89.125 ;
        RECT -289.545 88.945 -289.375 89.115 ;
        RECT -285.060 88.975 -284.890 89.145 ;
        RECT -283.695 88.975 -283.525 89.145 ;
        RECT -275.140 88.975 -274.970 89.145 ;
        RECT -273.775 88.975 -273.605 89.145 ;
        RECT -265.220 88.975 -265.050 89.145 ;
        RECT -263.855 88.975 -263.685 89.145 ;
        RECT -255.300 88.975 -255.130 89.145 ;
        RECT -253.935 88.975 -253.765 89.145 ;
        RECT -245.380 88.975 -245.210 89.145 ;
        RECT -244.015 88.975 -243.845 89.145 ;
        RECT -235.460 88.975 -235.290 89.145 ;
        RECT -234.095 88.975 -233.925 89.145 ;
        RECT -225.540 88.975 -225.370 89.145 ;
        RECT -224.175 88.975 -224.005 89.145 ;
        RECT -215.620 88.975 -215.450 89.145 ;
        RECT -214.255 88.975 -214.085 89.145 ;
        RECT -205.700 88.975 -205.530 89.145 ;
        RECT -204.335 88.975 -204.165 89.145 ;
        RECT -195.780 88.975 -195.610 89.145 ;
        RECT -194.415 88.975 -194.245 89.145 ;
        RECT -185.860 88.975 -185.690 89.145 ;
        RECT -184.495 88.975 -184.325 89.145 ;
        RECT -175.940 88.975 -175.770 89.145 ;
        RECT -174.575 88.975 -174.405 89.145 ;
        RECT -166.020 88.975 -165.850 89.145 ;
        RECT -164.655 88.975 -164.485 89.145 ;
        RECT -156.100 88.975 -155.930 89.145 ;
        RECT -154.735 88.975 -154.565 89.145 ;
        RECT -146.180 88.975 -146.010 89.145 ;
        RECT -144.815 88.975 -144.645 89.145 ;
        RECT -136.260 88.975 -136.090 89.145 ;
        RECT -134.895 88.975 -134.725 89.145 ;
        RECT -126.340 88.975 -126.170 89.145 ;
        RECT -124.975 88.975 -124.805 89.145 ;
        RECT -116.420 88.975 -116.250 89.145 ;
        RECT -115.055 88.975 -114.885 89.145 ;
        RECT -106.500 88.975 -106.330 89.145 ;
        RECT -105.135 88.975 -104.965 89.145 ;
        RECT -96.580 88.975 -96.410 89.145 ;
        RECT -95.215 88.975 -95.045 89.145 ;
        RECT -86.660 88.975 -86.490 89.145 ;
        RECT -85.295 88.975 -85.125 89.145 ;
        RECT -76.740 88.975 -76.570 89.145 ;
        RECT -75.375 88.975 -75.205 89.145 ;
        RECT -66.820 88.975 -66.650 89.145 ;
        RECT -65.455 88.975 -65.285 89.145 ;
        RECT -56.900 88.975 -56.730 89.145 ;
        RECT -55.535 88.975 -55.365 89.145 ;
        RECT -46.980 88.975 -46.810 89.145 ;
        RECT -45.615 88.975 -45.445 89.145 ;
        RECT -37.060 88.975 -36.890 89.145 ;
        RECT -35.695 88.975 -35.525 89.145 ;
        RECT -27.140 88.975 -26.970 89.145 ;
        RECT -25.775 88.975 -25.605 89.145 ;
        RECT -17.220 88.975 -17.050 89.145 ;
        RECT -15.855 88.975 -15.685 89.145 ;
        RECT -7.300 88.975 -7.130 89.145 ;
        RECT -5.935 88.975 -5.765 89.145 ;
        RECT 2.620 88.975 2.790 89.145 ;
        RECT 3.985 88.975 4.155 89.145 ;
        RECT 12.540 88.975 12.710 89.145 ;
        RECT 13.905 88.975 14.075 89.145 ;
        RECT 22.460 88.975 22.630 89.145 ;
        RECT 23.825 88.975 23.995 89.145 ;
        RECT 24.355 88.945 24.525 89.115 ;
        RECT 24.825 88.955 24.995 89.125 ;
        RECT -293.335 10.770 -293.165 10.940 ;
        RECT -292.865 10.775 -292.695 10.945 ;
        RECT -292.040 10.745 -291.870 10.915 ;
        RECT -290.675 10.745 -290.505 10.915 ;
        RECT -282.120 10.745 -281.950 10.915 ;
        RECT -280.755 10.745 -280.585 10.915 ;
        RECT -272.200 10.745 -272.030 10.915 ;
        RECT -270.835 10.745 -270.665 10.915 ;
        RECT -262.280 10.745 -262.110 10.915 ;
        RECT -260.915 10.745 -260.745 10.915 ;
        RECT -252.360 10.745 -252.190 10.915 ;
        RECT -250.995 10.745 -250.825 10.915 ;
        RECT -242.440 10.745 -242.270 10.915 ;
        RECT -241.075 10.745 -240.905 10.915 ;
        RECT -232.520 10.745 -232.350 10.915 ;
        RECT -231.155 10.745 -230.985 10.915 ;
        RECT -222.600 10.745 -222.430 10.915 ;
        RECT -221.235 10.745 -221.065 10.915 ;
        RECT -212.680 10.745 -212.510 10.915 ;
        RECT -211.315 10.745 -211.145 10.915 ;
        RECT -202.760 10.745 -202.590 10.915 ;
        RECT -201.395 10.745 -201.225 10.915 ;
        RECT -192.840 10.745 -192.670 10.915 ;
        RECT -191.475 10.745 -191.305 10.915 ;
        RECT -182.920 10.745 -182.750 10.915 ;
        RECT -181.555 10.745 -181.385 10.915 ;
        RECT -173.000 10.745 -172.830 10.915 ;
        RECT -171.635 10.745 -171.465 10.915 ;
        RECT -163.080 10.745 -162.910 10.915 ;
        RECT -161.715 10.745 -161.545 10.915 ;
        RECT -153.160 10.745 -152.990 10.915 ;
        RECT -151.795 10.745 -151.625 10.915 ;
        RECT -143.240 10.745 -143.070 10.915 ;
        RECT -141.875 10.745 -141.705 10.915 ;
        RECT -133.320 10.745 -133.150 10.915 ;
        RECT -131.955 10.745 -131.785 10.915 ;
        RECT -123.400 10.745 -123.230 10.915 ;
        RECT -122.035 10.745 -121.865 10.915 ;
        RECT -113.480 10.745 -113.310 10.915 ;
        RECT -112.115 10.745 -111.945 10.915 ;
        RECT -103.560 10.745 -103.390 10.915 ;
        RECT -102.195 10.745 -102.025 10.915 ;
        RECT -93.640 10.745 -93.470 10.915 ;
        RECT -92.275 10.745 -92.105 10.915 ;
        RECT -83.720 10.745 -83.550 10.915 ;
        RECT -82.355 10.745 -82.185 10.915 ;
        RECT -73.800 10.745 -73.630 10.915 ;
        RECT -72.435 10.745 -72.265 10.915 ;
        RECT -63.880 10.745 -63.710 10.915 ;
        RECT -62.515 10.745 -62.345 10.915 ;
        RECT -53.960 10.745 -53.790 10.915 ;
        RECT -52.595 10.745 -52.425 10.915 ;
        RECT -44.040 10.745 -43.870 10.915 ;
        RECT -42.675 10.745 -42.505 10.915 ;
        RECT -34.120 10.745 -33.950 10.915 ;
        RECT -32.755 10.745 -32.585 10.915 ;
        RECT -24.200 10.745 -24.030 10.915 ;
        RECT -22.835 10.745 -22.665 10.915 ;
        RECT -14.280 10.745 -14.110 10.915 ;
        RECT -12.915 10.745 -12.745 10.915 ;
        RECT -4.360 10.745 -4.190 10.915 ;
        RECT -2.995 10.745 -2.825 10.915 ;
        RECT 5.560 10.745 5.730 10.915 ;
        RECT 6.925 10.745 7.095 10.915 ;
        RECT 15.480 10.745 15.650 10.915 ;
        RECT 16.845 10.745 17.015 10.915 ;
        RECT -292.865 10.315 -292.695 10.485 ;
        RECT -292.865 9.855 -292.695 10.025 ;
        RECT -291.305 9.895 -291.135 10.065 ;
        RECT -285.445 9.895 -285.275 10.065 ;
        RECT -281.385 9.895 -281.215 10.065 ;
        RECT -275.525 9.895 -275.355 10.065 ;
        RECT -271.465 9.895 -271.295 10.065 ;
        RECT -265.605 9.895 -265.435 10.065 ;
        RECT -261.545 9.895 -261.375 10.065 ;
        RECT -255.685 9.895 -255.515 10.065 ;
        RECT -251.625 9.895 -251.455 10.065 ;
        RECT -245.765 9.895 -245.595 10.065 ;
        RECT -241.705 9.895 -241.535 10.065 ;
        RECT -235.845 9.895 -235.675 10.065 ;
        RECT -231.785 9.895 -231.615 10.065 ;
        RECT -225.925 9.895 -225.755 10.065 ;
        RECT -221.865 9.895 -221.695 10.065 ;
        RECT -216.005 9.895 -215.835 10.065 ;
        RECT -211.945 9.895 -211.775 10.065 ;
        RECT -206.085 9.895 -205.915 10.065 ;
        RECT -202.025 9.895 -201.855 10.065 ;
        RECT -196.165 9.895 -195.995 10.065 ;
        RECT -192.105 9.895 -191.935 10.065 ;
        RECT -186.245 9.895 -186.075 10.065 ;
        RECT -182.185 9.895 -182.015 10.065 ;
        RECT -176.325 9.895 -176.155 10.065 ;
        RECT -172.265 9.895 -172.095 10.065 ;
        RECT -166.405 9.895 -166.235 10.065 ;
        RECT -162.345 9.895 -162.175 10.065 ;
        RECT -156.485 9.895 -156.315 10.065 ;
        RECT -152.425 9.895 -152.255 10.065 ;
        RECT -146.565 9.895 -146.395 10.065 ;
        RECT -142.505 9.895 -142.335 10.065 ;
        RECT -136.645 9.895 -136.475 10.065 ;
        RECT -132.585 9.895 -132.415 10.065 ;
        RECT -126.725 9.895 -126.555 10.065 ;
        RECT -122.665 9.895 -122.495 10.065 ;
        RECT -116.805 9.895 -116.635 10.065 ;
        RECT -112.745 9.895 -112.575 10.065 ;
        RECT -106.885 9.895 -106.715 10.065 ;
        RECT -102.825 9.895 -102.655 10.065 ;
        RECT -96.965 9.895 -96.795 10.065 ;
        RECT -92.905 9.895 -92.735 10.065 ;
        RECT -87.045 9.895 -86.875 10.065 ;
        RECT -82.985 9.895 -82.815 10.065 ;
        RECT -77.125 9.895 -76.955 10.065 ;
        RECT -73.065 9.895 -72.895 10.065 ;
        RECT -67.205 9.895 -67.035 10.065 ;
        RECT -63.145 9.895 -62.975 10.065 ;
        RECT -57.285 9.895 -57.115 10.065 ;
        RECT -53.225 9.895 -53.055 10.065 ;
        RECT -47.365 9.895 -47.195 10.065 ;
        RECT -43.305 9.895 -43.135 10.065 ;
        RECT -37.445 9.895 -37.275 10.065 ;
        RECT -33.385 9.895 -33.215 10.065 ;
        RECT -27.525 9.895 -27.355 10.065 ;
        RECT -23.465 9.895 -23.295 10.065 ;
        RECT -17.605 9.895 -17.435 10.065 ;
        RECT -13.545 9.895 -13.375 10.065 ;
        RECT -7.685 9.895 -7.515 10.065 ;
        RECT -3.625 9.895 -3.455 10.065 ;
        RECT 2.235 9.895 2.405 10.065 ;
        RECT 6.295 9.895 6.465 10.065 ;
        RECT 12.155 9.895 12.325 10.065 ;
        RECT 16.215 9.895 16.385 10.065 ;
        RECT 22.075 9.895 22.245 10.065 ;
        RECT -293.335 9.195 -293.165 9.365 ;
        RECT -292.875 9.195 -292.705 9.365 ;
        RECT -292.415 9.195 -292.245 9.365 ;
        RECT -291.955 9.195 -291.785 9.365 ;
        RECT 22.725 9.195 22.895 9.365 ;
        RECT 23.185 9.195 23.355 9.365 ;
        RECT 23.645 9.195 23.815 9.365 ;
        RECT 24.105 9.195 24.275 9.365 ;
        RECT -291.985 8.475 -291.815 8.645 ;
        RECT -292.000 8.035 -291.830 8.205 ;
        RECT -284.765 8.475 -284.595 8.645 ;
        RECT -289.710 7.635 -289.540 7.805 ;
        RECT -289.725 7.195 -289.555 7.365 ;
        RECT -284.750 8.035 -284.580 8.205 ;
        RECT -287.040 7.635 -286.870 7.805 ;
        RECT -282.065 8.475 -281.895 8.645 ;
        RECT -282.080 8.035 -281.910 8.205 ;
        RECT -274.845 8.475 -274.675 8.645 ;
        RECT -287.025 7.195 -286.855 7.365 ;
        RECT -279.790 7.635 -279.620 7.805 ;
        RECT -279.805 7.195 -279.635 7.365 ;
        RECT -274.830 8.035 -274.660 8.205 ;
        RECT -277.120 7.635 -276.950 7.805 ;
        RECT -272.145 8.475 -271.975 8.645 ;
        RECT -272.160 8.035 -271.990 8.205 ;
        RECT -264.925 8.475 -264.755 8.645 ;
        RECT -277.105 7.195 -276.935 7.365 ;
        RECT -269.870 7.635 -269.700 7.805 ;
        RECT -269.885 7.195 -269.715 7.365 ;
        RECT -264.910 8.035 -264.740 8.205 ;
        RECT -267.200 7.635 -267.030 7.805 ;
        RECT -262.225 8.475 -262.055 8.645 ;
        RECT -262.240 8.035 -262.070 8.205 ;
        RECT -255.005 8.475 -254.835 8.645 ;
        RECT -267.185 7.195 -267.015 7.365 ;
        RECT -259.950 7.635 -259.780 7.805 ;
        RECT -259.965 7.195 -259.795 7.365 ;
        RECT -254.990 8.035 -254.820 8.205 ;
        RECT -257.280 7.635 -257.110 7.805 ;
        RECT -252.305 8.475 -252.135 8.645 ;
        RECT -252.320 8.035 -252.150 8.205 ;
        RECT -245.085 8.475 -244.915 8.645 ;
        RECT -257.265 7.195 -257.095 7.365 ;
        RECT -250.030 7.635 -249.860 7.805 ;
        RECT -250.045 7.195 -249.875 7.365 ;
        RECT -245.070 8.035 -244.900 8.205 ;
        RECT -247.360 7.635 -247.190 7.805 ;
        RECT -242.385 8.475 -242.215 8.645 ;
        RECT -242.400 8.035 -242.230 8.205 ;
        RECT -235.165 8.475 -234.995 8.645 ;
        RECT -247.345 7.195 -247.175 7.365 ;
        RECT -240.110 7.635 -239.940 7.805 ;
        RECT -240.125 7.195 -239.955 7.365 ;
        RECT -235.150 8.035 -234.980 8.205 ;
        RECT -237.440 7.635 -237.270 7.805 ;
        RECT -232.465 8.475 -232.295 8.645 ;
        RECT -232.480 8.035 -232.310 8.205 ;
        RECT -225.245 8.475 -225.075 8.645 ;
        RECT -237.425 7.195 -237.255 7.365 ;
        RECT -230.190 7.635 -230.020 7.805 ;
        RECT -230.205 7.195 -230.035 7.365 ;
        RECT -225.230 8.035 -225.060 8.205 ;
        RECT -227.520 7.635 -227.350 7.805 ;
        RECT -222.545 8.475 -222.375 8.645 ;
        RECT -222.560 8.035 -222.390 8.205 ;
        RECT -215.325 8.475 -215.155 8.645 ;
        RECT -227.505 7.195 -227.335 7.365 ;
        RECT -220.270 7.635 -220.100 7.805 ;
        RECT -220.285 7.195 -220.115 7.365 ;
        RECT -215.310 8.035 -215.140 8.205 ;
        RECT -217.600 7.635 -217.430 7.805 ;
        RECT -212.625 8.475 -212.455 8.645 ;
        RECT -212.640 8.035 -212.470 8.205 ;
        RECT -205.405 8.475 -205.235 8.645 ;
        RECT -217.585 7.195 -217.415 7.365 ;
        RECT -210.350 7.635 -210.180 7.805 ;
        RECT -210.365 7.195 -210.195 7.365 ;
        RECT -205.390 8.035 -205.220 8.205 ;
        RECT -207.680 7.635 -207.510 7.805 ;
        RECT -202.705 8.475 -202.535 8.645 ;
        RECT -202.720 8.035 -202.550 8.205 ;
        RECT -195.485 8.475 -195.315 8.645 ;
        RECT -207.665 7.195 -207.495 7.365 ;
        RECT -200.430 7.635 -200.260 7.805 ;
        RECT -200.445 7.195 -200.275 7.365 ;
        RECT -195.470 8.035 -195.300 8.205 ;
        RECT -197.760 7.635 -197.590 7.805 ;
        RECT -192.785 8.475 -192.615 8.645 ;
        RECT -192.800 8.035 -192.630 8.205 ;
        RECT -185.565 8.475 -185.395 8.645 ;
        RECT -197.745 7.195 -197.575 7.365 ;
        RECT -190.510 7.635 -190.340 7.805 ;
        RECT -190.525 7.195 -190.355 7.365 ;
        RECT -185.550 8.035 -185.380 8.205 ;
        RECT -187.840 7.635 -187.670 7.805 ;
        RECT -182.865 8.475 -182.695 8.645 ;
        RECT -182.880 8.035 -182.710 8.205 ;
        RECT -175.645 8.475 -175.475 8.645 ;
        RECT -187.825 7.195 -187.655 7.365 ;
        RECT -180.590 7.635 -180.420 7.805 ;
        RECT -180.605 7.195 -180.435 7.365 ;
        RECT -175.630 8.035 -175.460 8.205 ;
        RECT -177.920 7.635 -177.750 7.805 ;
        RECT -172.945 8.475 -172.775 8.645 ;
        RECT -172.960 8.035 -172.790 8.205 ;
        RECT -165.725 8.475 -165.555 8.645 ;
        RECT -177.905 7.195 -177.735 7.365 ;
        RECT -170.670 7.635 -170.500 7.805 ;
        RECT -170.685 7.195 -170.515 7.365 ;
        RECT -165.710 8.035 -165.540 8.205 ;
        RECT -168.000 7.635 -167.830 7.805 ;
        RECT -163.025 8.475 -162.855 8.645 ;
        RECT -163.040 8.035 -162.870 8.205 ;
        RECT -155.805 8.475 -155.635 8.645 ;
        RECT -167.985 7.195 -167.815 7.365 ;
        RECT -160.750 7.635 -160.580 7.805 ;
        RECT -160.765 7.195 -160.595 7.365 ;
        RECT -155.790 8.035 -155.620 8.205 ;
        RECT -158.080 7.635 -157.910 7.805 ;
        RECT -153.105 8.475 -152.935 8.645 ;
        RECT -153.120 8.035 -152.950 8.205 ;
        RECT -145.885 8.475 -145.715 8.645 ;
        RECT -158.065 7.195 -157.895 7.365 ;
        RECT -150.830 7.635 -150.660 7.805 ;
        RECT -150.845 7.195 -150.675 7.365 ;
        RECT -145.870 8.035 -145.700 8.205 ;
        RECT -148.160 7.635 -147.990 7.805 ;
        RECT -143.185 8.475 -143.015 8.645 ;
        RECT -143.200 8.035 -143.030 8.205 ;
        RECT -135.965 8.475 -135.795 8.645 ;
        RECT -148.145 7.195 -147.975 7.365 ;
        RECT -140.910 7.635 -140.740 7.805 ;
        RECT -140.925 7.195 -140.755 7.365 ;
        RECT -135.950 8.035 -135.780 8.205 ;
        RECT -138.240 7.635 -138.070 7.805 ;
        RECT -133.265 8.475 -133.095 8.645 ;
        RECT -133.280 8.035 -133.110 8.205 ;
        RECT -126.045 8.475 -125.875 8.645 ;
        RECT -138.225 7.195 -138.055 7.365 ;
        RECT -130.990 7.635 -130.820 7.805 ;
        RECT -131.005 7.195 -130.835 7.365 ;
        RECT -126.030 8.035 -125.860 8.205 ;
        RECT -128.320 7.635 -128.150 7.805 ;
        RECT -123.345 8.475 -123.175 8.645 ;
        RECT -123.360 8.035 -123.190 8.205 ;
        RECT -116.125 8.475 -115.955 8.645 ;
        RECT -128.305 7.195 -128.135 7.365 ;
        RECT -121.070 7.635 -120.900 7.805 ;
        RECT -121.085 7.195 -120.915 7.365 ;
        RECT -116.110 8.035 -115.940 8.205 ;
        RECT -118.400 7.635 -118.230 7.805 ;
        RECT -113.425 8.475 -113.255 8.645 ;
        RECT -113.440 8.035 -113.270 8.205 ;
        RECT -106.205 8.475 -106.035 8.645 ;
        RECT -118.385 7.195 -118.215 7.365 ;
        RECT -111.150 7.635 -110.980 7.805 ;
        RECT -111.165 7.195 -110.995 7.365 ;
        RECT -106.190 8.035 -106.020 8.205 ;
        RECT -108.480 7.635 -108.310 7.805 ;
        RECT -103.505 8.475 -103.335 8.645 ;
        RECT -103.520 8.035 -103.350 8.205 ;
        RECT -96.285 8.475 -96.115 8.645 ;
        RECT -108.465 7.195 -108.295 7.365 ;
        RECT -101.230 7.635 -101.060 7.805 ;
        RECT -101.245 7.195 -101.075 7.365 ;
        RECT -96.270 8.035 -96.100 8.205 ;
        RECT -98.560 7.635 -98.390 7.805 ;
        RECT -93.585 8.475 -93.415 8.645 ;
        RECT -93.600 8.035 -93.430 8.205 ;
        RECT -86.365 8.475 -86.195 8.645 ;
        RECT -98.545 7.195 -98.375 7.365 ;
        RECT -91.310 7.635 -91.140 7.805 ;
        RECT -91.325 7.195 -91.155 7.365 ;
        RECT -86.350 8.035 -86.180 8.205 ;
        RECT -88.640 7.635 -88.470 7.805 ;
        RECT -83.665 8.475 -83.495 8.645 ;
        RECT -83.680 8.035 -83.510 8.205 ;
        RECT -76.445 8.475 -76.275 8.645 ;
        RECT -88.625 7.195 -88.455 7.365 ;
        RECT -81.390 7.635 -81.220 7.805 ;
        RECT -81.405 7.195 -81.235 7.365 ;
        RECT -76.430 8.035 -76.260 8.205 ;
        RECT -78.720 7.635 -78.550 7.805 ;
        RECT -73.745 8.475 -73.575 8.645 ;
        RECT -73.760 8.035 -73.590 8.205 ;
        RECT -66.525 8.475 -66.355 8.645 ;
        RECT -78.705 7.195 -78.535 7.365 ;
        RECT -71.470 7.635 -71.300 7.805 ;
        RECT -71.485 7.195 -71.315 7.365 ;
        RECT -66.510 8.035 -66.340 8.205 ;
        RECT -68.800 7.635 -68.630 7.805 ;
        RECT -63.825 8.475 -63.655 8.645 ;
        RECT -63.840 8.035 -63.670 8.205 ;
        RECT -56.605 8.475 -56.435 8.645 ;
        RECT -68.785 7.195 -68.615 7.365 ;
        RECT -61.550 7.635 -61.380 7.805 ;
        RECT -61.565 7.195 -61.395 7.365 ;
        RECT -56.590 8.035 -56.420 8.205 ;
        RECT -58.880 7.635 -58.710 7.805 ;
        RECT -53.905 8.475 -53.735 8.645 ;
        RECT -53.920 8.035 -53.750 8.205 ;
        RECT -46.685 8.475 -46.515 8.645 ;
        RECT -58.865 7.195 -58.695 7.365 ;
        RECT -51.630 7.635 -51.460 7.805 ;
        RECT -51.645 7.195 -51.475 7.365 ;
        RECT -46.670 8.035 -46.500 8.205 ;
        RECT -48.960 7.635 -48.790 7.805 ;
        RECT -43.985 8.475 -43.815 8.645 ;
        RECT -44.000 8.035 -43.830 8.205 ;
        RECT -36.765 8.475 -36.595 8.645 ;
        RECT -48.945 7.195 -48.775 7.365 ;
        RECT -41.710 7.635 -41.540 7.805 ;
        RECT -41.725 7.195 -41.555 7.365 ;
        RECT -36.750 8.035 -36.580 8.205 ;
        RECT -39.040 7.635 -38.870 7.805 ;
        RECT -34.065 8.475 -33.895 8.645 ;
        RECT -34.080 8.035 -33.910 8.205 ;
        RECT -26.845 8.475 -26.675 8.645 ;
        RECT -39.025 7.195 -38.855 7.365 ;
        RECT -31.790 7.635 -31.620 7.805 ;
        RECT -31.805 7.195 -31.635 7.365 ;
        RECT -26.830 8.035 -26.660 8.205 ;
        RECT -29.120 7.635 -28.950 7.805 ;
        RECT -24.145 8.475 -23.975 8.645 ;
        RECT -24.160 8.035 -23.990 8.205 ;
        RECT -16.925 8.475 -16.755 8.645 ;
        RECT -29.105 7.195 -28.935 7.365 ;
        RECT -21.870 7.635 -21.700 7.805 ;
        RECT -21.885 7.195 -21.715 7.365 ;
        RECT -16.910 8.035 -16.740 8.205 ;
        RECT -19.200 7.635 -19.030 7.805 ;
        RECT -14.225 8.475 -14.055 8.645 ;
        RECT -14.240 8.035 -14.070 8.205 ;
        RECT -7.005 8.475 -6.835 8.645 ;
        RECT -19.185 7.195 -19.015 7.365 ;
        RECT -11.950 7.635 -11.780 7.805 ;
        RECT -11.965 7.195 -11.795 7.365 ;
        RECT -6.990 8.035 -6.820 8.205 ;
        RECT -9.280 7.635 -9.110 7.805 ;
        RECT -4.305 8.475 -4.135 8.645 ;
        RECT -4.320 8.035 -4.150 8.205 ;
        RECT 2.915 8.475 3.085 8.645 ;
        RECT -9.265 7.195 -9.095 7.365 ;
        RECT -2.030 7.635 -1.860 7.805 ;
        RECT -2.045 7.195 -1.875 7.365 ;
        RECT 2.930 8.035 3.100 8.205 ;
        RECT 0.640 7.635 0.810 7.805 ;
        RECT 5.615 8.475 5.785 8.645 ;
        RECT 5.600 8.035 5.770 8.205 ;
        RECT 12.835 8.475 13.005 8.645 ;
        RECT 0.655 7.195 0.825 7.365 ;
        RECT 7.890 7.635 8.060 7.805 ;
        RECT 7.875 7.195 8.045 7.365 ;
        RECT 12.850 8.035 13.020 8.205 ;
        RECT 10.560 7.635 10.730 7.805 ;
        RECT 15.535 8.475 15.705 8.645 ;
        RECT 15.520 8.035 15.690 8.205 ;
        RECT 22.755 8.475 22.925 8.645 ;
        RECT 10.575 7.195 10.745 7.365 ;
        RECT 17.810 7.635 17.980 7.805 ;
        RECT 17.795 7.195 17.965 7.365 ;
        RECT 22.770 8.035 22.940 8.205 ;
        RECT 20.480 7.635 20.650 7.805 ;
        RECT 20.495 7.195 20.665 7.365 ;
        RECT -293.335 6.475 -293.165 6.645 ;
        RECT -292.875 6.475 -292.705 6.645 ;
        RECT -292.415 6.475 -292.245 6.645 ;
        RECT -291.955 6.475 -291.785 6.645 ;
        RECT -291.565 5.815 -291.395 5.985 ;
        RECT -291.565 5.355 -291.395 5.525 ;
        RECT -290.405 5.775 -290.235 5.945 ;
        RECT -286.345 5.775 -286.175 5.945 ;
        RECT -280.485 5.775 -280.315 5.945 ;
        RECT -276.425 5.775 -276.255 5.945 ;
        RECT -270.565 5.775 -270.395 5.945 ;
        RECT -266.505 5.775 -266.335 5.945 ;
        RECT -260.645 5.775 -260.475 5.945 ;
        RECT -256.585 5.775 -256.415 5.945 ;
        RECT -250.725 5.775 -250.555 5.945 ;
        RECT -246.665 5.775 -246.495 5.945 ;
        RECT -240.805 5.775 -240.635 5.945 ;
        RECT -236.745 5.775 -236.575 5.945 ;
        RECT -230.885 5.775 -230.715 5.945 ;
        RECT -226.825 5.775 -226.655 5.945 ;
        RECT -220.965 5.775 -220.795 5.945 ;
        RECT -216.905 5.775 -216.735 5.945 ;
        RECT -211.045 5.775 -210.875 5.945 ;
        RECT -206.985 5.775 -206.815 5.945 ;
        RECT -201.125 5.775 -200.955 5.945 ;
        RECT -197.065 5.775 -196.895 5.945 ;
        RECT -191.205 5.775 -191.035 5.945 ;
        RECT -187.145 5.775 -186.975 5.945 ;
        RECT -181.285 5.775 -181.115 5.945 ;
        RECT -177.225 5.775 -177.055 5.945 ;
        RECT -171.365 5.775 -171.195 5.945 ;
        RECT -167.305 5.775 -167.135 5.945 ;
        RECT -161.445 5.775 -161.275 5.945 ;
        RECT -157.385 5.775 -157.215 5.945 ;
        RECT -151.525 5.775 -151.355 5.945 ;
        RECT -147.465 5.775 -147.295 5.945 ;
        RECT -141.605 5.775 -141.435 5.945 ;
        RECT -137.545 5.775 -137.375 5.945 ;
        RECT -131.685 5.775 -131.515 5.945 ;
        RECT -127.625 5.775 -127.455 5.945 ;
        RECT -121.765 5.775 -121.595 5.945 ;
        RECT -117.705 5.775 -117.535 5.945 ;
        RECT -111.845 5.775 -111.675 5.945 ;
        RECT -107.785 5.775 -107.615 5.945 ;
        RECT -101.925 5.775 -101.755 5.945 ;
        RECT -97.865 5.775 -97.695 5.945 ;
        RECT -92.005 5.775 -91.835 5.945 ;
        RECT -87.945 5.775 -87.775 5.945 ;
        RECT -82.085 5.775 -81.915 5.945 ;
        RECT -78.025 5.775 -77.855 5.945 ;
        RECT -72.165 5.775 -71.995 5.945 ;
        RECT -68.105 5.775 -67.935 5.945 ;
        RECT -62.245 5.775 -62.075 5.945 ;
        RECT -58.185 5.775 -58.015 5.945 ;
        RECT -52.325 5.775 -52.155 5.945 ;
        RECT -48.265 5.775 -48.095 5.945 ;
        RECT -42.405 5.775 -42.235 5.945 ;
        RECT -38.345 5.775 -38.175 5.945 ;
        RECT -32.485 5.775 -32.315 5.945 ;
        RECT -28.425 5.775 -28.255 5.945 ;
        RECT -22.565 5.775 -22.395 5.945 ;
        RECT -18.505 5.775 -18.335 5.945 ;
        RECT -12.645 5.775 -12.475 5.945 ;
        RECT -8.585 5.775 -8.415 5.945 ;
        RECT -2.725 5.775 -2.555 5.945 ;
        RECT 1.335 5.775 1.505 5.945 ;
        RECT 7.195 5.775 7.365 5.945 ;
        RECT 11.255 5.775 11.425 5.945 ;
        RECT 17.115 5.775 17.285 5.945 ;
        RECT 21.175 5.775 21.345 5.945 ;
        RECT 22.335 5.815 22.505 5.985 ;
        RECT 22.335 5.355 22.505 5.525 ;
        RECT -292.035 4.905 -291.865 5.075 ;
        RECT -291.565 4.895 -291.395 5.065 ;
        RECT -287.080 4.925 -286.910 5.095 ;
        RECT -285.715 4.925 -285.545 5.095 ;
        RECT -277.160 4.925 -276.990 5.095 ;
        RECT -275.795 4.925 -275.625 5.095 ;
        RECT -267.240 4.925 -267.070 5.095 ;
        RECT -265.875 4.925 -265.705 5.095 ;
        RECT -257.320 4.925 -257.150 5.095 ;
        RECT -255.955 4.925 -255.785 5.095 ;
        RECT -247.400 4.925 -247.230 5.095 ;
        RECT -246.035 4.925 -245.865 5.095 ;
        RECT -237.480 4.925 -237.310 5.095 ;
        RECT -236.115 4.925 -235.945 5.095 ;
        RECT -227.560 4.925 -227.390 5.095 ;
        RECT -226.195 4.925 -226.025 5.095 ;
        RECT -217.640 4.925 -217.470 5.095 ;
        RECT -216.275 4.925 -216.105 5.095 ;
        RECT -207.720 4.925 -207.550 5.095 ;
        RECT -206.355 4.925 -206.185 5.095 ;
        RECT -197.800 4.925 -197.630 5.095 ;
        RECT -196.435 4.925 -196.265 5.095 ;
        RECT -187.880 4.925 -187.710 5.095 ;
        RECT -186.515 4.925 -186.345 5.095 ;
        RECT -177.960 4.925 -177.790 5.095 ;
        RECT -176.595 4.925 -176.425 5.095 ;
        RECT -168.040 4.925 -167.870 5.095 ;
        RECT -166.675 4.925 -166.505 5.095 ;
        RECT -158.120 4.925 -157.950 5.095 ;
        RECT -156.755 4.925 -156.585 5.095 ;
        RECT -148.200 4.925 -148.030 5.095 ;
        RECT -146.835 4.925 -146.665 5.095 ;
        RECT -138.280 4.925 -138.110 5.095 ;
        RECT -136.915 4.925 -136.745 5.095 ;
        RECT -128.360 4.925 -128.190 5.095 ;
        RECT -126.995 4.925 -126.825 5.095 ;
        RECT -118.440 4.925 -118.270 5.095 ;
        RECT -117.075 4.925 -116.905 5.095 ;
        RECT -108.520 4.925 -108.350 5.095 ;
        RECT -107.155 4.925 -106.985 5.095 ;
        RECT -98.600 4.925 -98.430 5.095 ;
        RECT -97.235 4.925 -97.065 5.095 ;
        RECT -88.680 4.925 -88.510 5.095 ;
        RECT -87.315 4.925 -87.145 5.095 ;
        RECT -78.760 4.925 -78.590 5.095 ;
        RECT -77.395 4.925 -77.225 5.095 ;
        RECT -68.840 4.925 -68.670 5.095 ;
        RECT -67.475 4.925 -67.305 5.095 ;
        RECT -58.920 4.925 -58.750 5.095 ;
        RECT -57.555 4.925 -57.385 5.095 ;
        RECT -49.000 4.925 -48.830 5.095 ;
        RECT -47.635 4.925 -47.465 5.095 ;
        RECT -39.080 4.925 -38.910 5.095 ;
        RECT -37.715 4.925 -37.545 5.095 ;
        RECT -29.160 4.925 -28.990 5.095 ;
        RECT -27.795 4.925 -27.625 5.095 ;
        RECT -19.240 4.925 -19.070 5.095 ;
        RECT -17.875 4.925 -17.705 5.095 ;
        RECT -9.320 4.925 -9.150 5.095 ;
        RECT -7.955 4.925 -7.785 5.095 ;
        RECT 0.600 4.925 0.770 5.095 ;
        RECT 1.965 4.925 2.135 5.095 ;
        RECT 10.520 4.925 10.690 5.095 ;
        RECT 11.885 4.925 12.055 5.095 ;
        RECT 20.440 4.925 20.610 5.095 ;
        RECT 21.805 4.925 21.975 5.095 ;
        RECT 22.335 4.895 22.505 5.065 ;
        RECT 22.805 4.905 22.975 5.075 ;
        RECT -292.975 -78.180 -292.805 -78.010 ;
        RECT -292.505 -78.175 -292.335 -78.005 ;
        RECT -291.680 -78.205 -291.510 -78.035 ;
        RECT -290.315 -78.205 -290.145 -78.035 ;
        RECT -281.760 -78.205 -281.590 -78.035 ;
        RECT -280.395 -78.205 -280.225 -78.035 ;
        RECT -271.840 -78.205 -271.670 -78.035 ;
        RECT -270.475 -78.205 -270.305 -78.035 ;
        RECT -261.920 -78.205 -261.750 -78.035 ;
        RECT -260.555 -78.205 -260.385 -78.035 ;
        RECT -252.000 -78.205 -251.830 -78.035 ;
        RECT -250.635 -78.205 -250.465 -78.035 ;
        RECT -242.080 -78.205 -241.910 -78.035 ;
        RECT -240.715 -78.205 -240.545 -78.035 ;
        RECT -232.160 -78.205 -231.990 -78.035 ;
        RECT -230.795 -78.205 -230.625 -78.035 ;
        RECT -222.240 -78.205 -222.070 -78.035 ;
        RECT -220.875 -78.205 -220.705 -78.035 ;
        RECT -212.320 -78.205 -212.150 -78.035 ;
        RECT -210.955 -78.205 -210.785 -78.035 ;
        RECT -202.400 -78.205 -202.230 -78.035 ;
        RECT -201.035 -78.205 -200.865 -78.035 ;
        RECT -192.480 -78.205 -192.310 -78.035 ;
        RECT -191.115 -78.205 -190.945 -78.035 ;
        RECT -182.560 -78.205 -182.390 -78.035 ;
        RECT -181.195 -78.205 -181.025 -78.035 ;
        RECT -172.640 -78.205 -172.470 -78.035 ;
        RECT -171.275 -78.205 -171.105 -78.035 ;
        RECT -162.720 -78.205 -162.550 -78.035 ;
        RECT -161.355 -78.205 -161.185 -78.035 ;
        RECT -152.800 -78.205 -152.630 -78.035 ;
        RECT -151.435 -78.205 -151.265 -78.035 ;
        RECT -142.880 -78.205 -142.710 -78.035 ;
        RECT -141.515 -78.205 -141.345 -78.035 ;
        RECT -132.960 -78.205 -132.790 -78.035 ;
        RECT -131.595 -78.205 -131.425 -78.035 ;
        RECT -123.040 -78.205 -122.870 -78.035 ;
        RECT -121.675 -78.205 -121.505 -78.035 ;
        RECT -113.120 -78.205 -112.950 -78.035 ;
        RECT -111.755 -78.205 -111.585 -78.035 ;
        RECT -103.200 -78.205 -103.030 -78.035 ;
        RECT -101.835 -78.205 -101.665 -78.035 ;
        RECT -93.280 -78.205 -93.110 -78.035 ;
        RECT -91.915 -78.205 -91.745 -78.035 ;
        RECT -83.360 -78.205 -83.190 -78.035 ;
        RECT -81.995 -78.205 -81.825 -78.035 ;
        RECT -73.440 -78.205 -73.270 -78.035 ;
        RECT -72.075 -78.205 -71.905 -78.035 ;
        RECT -63.520 -78.205 -63.350 -78.035 ;
        RECT -62.155 -78.205 -61.985 -78.035 ;
        RECT -53.600 -78.205 -53.430 -78.035 ;
        RECT -52.235 -78.205 -52.065 -78.035 ;
        RECT -43.680 -78.205 -43.510 -78.035 ;
        RECT -42.315 -78.205 -42.145 -78.035 ;
        RECT -33.760 -78.205 -33.590 -78.035 ;
        RECT -32.395 -78.205 -32.225 -78.035 ;
        RECT -23.840 -78.205 -23.670 -78.035 ;
        RECT -22.475 -78.205 -22.305 -78.035 ;
        RECT -13.920 -78.205 -13.750 -78.035 ;
        RECT -12.555 -78.205 -12.385 -78.035 ;
        RECT -4.000 -78.205 -3.830 -78.035 ;
        RECT -2.635 -78.205 -2.465 -78.035 ;
        RECT 5.920 -78.205 6.090 -78.035 ;
        RECT 7.285 -78.205 7.455 -78.035 ;
        RECT 15.840 -78.205 16.010 -78.035 ;
        RECT 17.205 -78.205 17.375 -78.035 ;
        RECT -292.505 -78.635 -292.335 -78.465 ;
        RECT -292.505 -79.095 -292.335 -78.925 ;
        RECT -290.945 -79.055 -290.775 -78.885 ;
        RECT -285.085 -79.055 -284.915 -78.885 ;
        RECT -281.025 -79.055 -280.855 -78.885 ;
        RECT -275.165 -79.055 -274.995 -78.885 ;
        RECT -271.105 -79.055 -270.935 -78.885 ;
        RECT -265.245 -79.055 -265.075 -78.885 ;
        RECT -261.185 -79.055 -261.015 -78.885 ;
        RECT -255.325 -79.055 -255.155 -78.885 ;
        RECT -251.265 -79.055 -251.095 -78.885 ;
        RECT -245.405 -79.055 -245.235 -78.885 ;
        RECT -241.345 -79.055 -241.175 -78.885 ;
        RECT -235.485 -79.055 -235.315 -78.885 ;
        RECT -231.425 -79.055 -231.255 -78.885 ;
        RECT -225.565 -79.055 -225.395 -78.885 ;
        RECT -221.505 -79.055 -221.335 -78.885 ;
        RECT -215.645 -79.055 -215.475 -78.885 ;
        RECT -211.585 -79.055 -211.415 -78.885 ;
        RECT -205.725 -79.055 -205.555 -78.885 ;
        RECT -201.665 -79.055 -201.495 -78.885 ;
        RECT -195.805 -79.055 -195.635 -78.885 ;
        RECT -191.745 -79.055 -191.575 -78.885 ;
        RECT -185.885 -79.055 -185.715 -78.885 ;
        RECT -181.825 -79.055 -181.655 -78.885 ;
        RECT -175.965 -79.055 -175.795 -78.885 ;
        RECT -171.905 -79.055 -171.735 -78.885 ;
        RECT -166.045 -79.055 -165.875 -78.885 ;
        RECT -161.985 -79.055 -161.815 -78.885 ;
        RECT -156.125 -79.055 -155.955 -78.885 ;
        RECT -152.065 -79.055 -151.895 -78.885 ;
        RECT -146.205 -79.055 -146.035 -78.885 ;
        RECT -142.145 -79.055 -141.975 -78.885 ;
        RECT -136.285 -79.055 -136.115 -78.885 ;
        RECT -132.225 -79.055 -132.055 -78.885 ;
        RECT -126.365 -79.055 -126.195 -78.885 ;
        RECT -122.305 -79.055 -122.135 -78.885 ;
        RECT -116.445 -79.055 -116.275 -78.885 ;
        RECT -112.385 -79.055 -112.215 -78.885 ;
        RECT -106.525 -79.055 -106.355 -78.885 ;
        RECT -102.465 -79.055 -102.295 -78.885 ;
        RECT -96.605 -79.055 -96.435 -78.885 ;
        RECT -92.545 -79.055 -92.375 -78.885 ;
        RECT -86.685 -79.055 -86.515 -78.885 ;
        RECT -82.625 -79.055 -82.455 -78.885 ;
        RECT -76.765 -79.055 -76.595 -78.885 ;
        RECT -72.705 -79.055 -72.535 -78.885 ;
        RECT -66.845 -79.055 -66.675 -78.885 ;
        RECT -62.785 -79.055 -62.615 -78.885 ;
        RECT -56.925 -79.055 -56.755 -78.885 ;
        RECT -52.865 -79.055 -52.695 -78.885 ;
        RECT -47.005 -79.055 -46.835 -78.885 ;
        RECT -42.945 -79.055 -42.775 -78.885 ;
        RECT -37.085 -79.055 -36.915 -78.885 ;
        RECT -33.025 -79.055 -32.855 -78.885 ;
        RECT -27.165 -79.055 -26.995 -78.885 ;
        RECT -23.105 -79.055 -22.935 -78.885 ;
        RECT -17.245 -79.055 -17.075 -78.885 ;
        RECT -13.185 -79.055 -13.015 -78.885 ;
        RECT -7.325 -79.055 -7.155 -78.885 ;
        RECT -3.265 -79.055 -3.095 -78.885 ;
        RECT 2.595 -79.055 2.765 -78.885 ;
        RECT 6.655 -79.055 6.825 -78.885 ;
        RECT 12.515 -79.055 12.685 -78.885 ;
        RECT 16.575 -79.055 16.745 -78.885 ;
        RECT 22.435 -79.055 22.605 -78.885 ;
        RECT -292.975 -79.755 -292.805 -79.585 ;
        RECT -292.515 -79.755 -292.345 -79.585 ;
        RECT -292.055 -79.755 -291.885 -79.585 ;
        RECT -291.595 -79.755 -291.425 -79.585 ;
        RECT 23.085 -79.755 23.255 -79.585 ;
        RECT 23.545 -79.755 23.715 -79.585 ;
        RECT 24.005 -79.755 24.175 -79.585 ;
        RECT 24.465 -79.755 24.635 -79.585 ;
        RECT -291.625 -80.475 -291.455 -80.305 ;
        RECT -291.640 -80.915 -291.470 -80.745 ;
        RECT -284.405 -80.475 -284.235 -80.305 ;
        RECT -289.350 -81.315 -289.180 -81.145 ;
        RECT -289.365 -81.755 -289.195 -81.585 ;
        RECT -284.390 -80.915 -284.220 -80.745 ;
        RECT -286.680 -81.315 -286.510 -81.145 ;
        RECT -281.705 -80.475 -281.535 -80.305 ;
        RECT -281.720 -80.915 -281.550 -80.745 ;
        RECT -274.485 -80.475 -274.315 -80.305 ;
        RECT -286.665 -81.755 -286.495 -81.585 ;
        RECT -279.430 -81.315 -279.260 -81.145 ;
        RECT -279.445 -81.755 -279.275 -81.585 ;
        RECT -274.470 -80.915 -274.300 -80.745 ;
        RECT -276.760 -81.315 -276.590 -81.145 ;
        RECT -271.785 -80.475 -271.615 -80.305 ;
        RECT -271.800 -80.915 -271.630 -80.745 ;
        RECT -264.565 -80.475 -264.395 -80.305 ;
        RECT -276.745 -81.755 -276.575 -81.585 ;
        RECT -269.510 -81.315 -269.340 -81.145 ;
        RECT -269.525 -81.755 -269.355 -81.585 ;
        RECT -264.550 -80.915 -264.380 -80.745 ;
        RECT -266.840 -81.315 -266.670 -81.145 ;
        RECT -261.865 -80.475 -261.695 -80.305 ;
        RECT -261.880 -80.915 -261.710 -80.745 ;
        RECT -254.645 -80.475 -254.475 -80.305 ;
        RECT -266.825 -81.755 -266.655 -81.585 ;
        RECT -259.590 -81.315 -259.420 -81.145 ;
        RECT -259.605 -81.755 -259.435 -81.585 ;
        RECT -254.630 -80.915 -254.460 -80.745 ;
        RECT -256.920 -81.315 -256.750 -81.145 ;
        RECT -251.945 -80.475 -251.775 -80.305 ;
        RECT -251.960 -80.915 -251.790 -80.745 ;
        RECT -244.725 -80.475 -244.555 -80.305 ;
        RECT -256.905 -81.755 -256.735 -81.585 ;
        RECT -249.670 -81.315 -249.500 -81.145 ;
        RECT -249.685 -81.755 -249.515 -81.585 ;
        RECT -244.710 -80.915 -244.540 -80.745 ;
        RECT -247.000 -81.315 -246.830 -81.145 ;
        RECT -242.025 -80.475 -241.855 -80.305 ;
        RECT -242.040 -80.915 -241.870 -80.745 ;
        RECT -234.805 -80.475 -234.635 -80.305 ;
        RECT -246.985 -81.755 -246.815 -81.585 ;
        RECT -239.750 -81.315 -239.580 -81.145 ;
        RECT -239.765 -81.755 -239.595 -81.585 ;
        RECT -234.790 -80.915 -234.620 -80.745 ;
        RECT -237.080 -81.315 -236.910 -81.145 ;
        RECT -232.105 -80.475 -231.935 -80.305 ;
        RECT -232.120 -80.915 -231.950 -80.745 ;
        RECT -224.885 -80.475 -224.715 -80.305 ;
        RECT -237.065 -81.755 -236.895 -81.585 ;
        RECT -229.830 -81.315 -229.660 -81.145 ;
        RECT -229.845 -81.755 -229.675 -81.585 ;
        RECT -224.870 -80.915 -224.700 -80.745 ;
        RECT -227.160 -81.315 -226.990 -81.145 ;
        RECT -222.185 -80.475 -222.015 -80.305 ;
        RECT -222.200 -80.915 -222.030 -80.745 ;
        RECT -214.965 -80.475 -214.795 -80.305 ;
        RECT -227.145 -81.755 -226.975 -81.585 ;
        RECT -219.910 -81.315 -219.740 -81.145 ;
        RECT -219.925 -81.755 -219.755 -81.585 ;
        RECT -214.950 -80.915 -214.780 -80.745 ;
        RECT -217.240 -81.315 -217.070 -81.145 ;
        RECT -212.265 -80.475 -212.095 -80.305 ;
        RECT -212.280 -80.915 -212.110 -80.745 ;
        RECT -205.045 -80.475 -204.875 -80.305 ;
        RECT -217.225 -81.755 -217.055 -81.585 ;
        RECT -209.990 -81.315 -209.820 -81.145 ;
        RECT -210.005 -81.755 -209.835 -81.585 ;
        RECT -205.030 -80.915 -204.860 -80.745 ;
        RECT -207.320 -81.315 -207.150 -81.145 ;
        RECT -202.345 -80.475 -202.175 -80.305 ;
        RECT -202.360 -80.915 -202.190 -80.745 ;
        RECT -195.125 -80.475 -194.955 -80.305 ;
        RECT -207.305 -81.755 -207.135 -81.585 ;
        RECT -200.070 -81.315 -199.900 -81.145 ;
        RECT -200.085 -81.755 -199.915 -81.585 ;
        RECT -195.110 -80.915 -194.940 -80.745 ;
        RECT -197.400 -81.315 -197.230 -81.145 ;
        RECT -192.425 -80.475 -192.255 -80.305 ;
        RECT -192.440 -80.915 -192.270 -80.745 ;
        RECT -185.205 -80.475 -185.035 -80.305 ;
        RECT -197.385 -81.755 -197.215 -81.585 ;
        RECT -190.150 -81.315 -189.980 -81.145 ;
        RECT -190.165 -81.755 -189.995 -81.585 ;
        RECT -185.190 -80.915 -185.020 -80.745 ;
        RECT -187.480 -81.315 -187.310 -81.145 ;
        RECT -182.505 -80.475 -182.335 -80.305 ;
        RECT -182.520 -80.915 -182.350 -80.745 ;
        RECT -175.285 -80.475 -175.115 -80.305 ;
        RECT -187.465 -81.755 -187.295 -81.585 ;
        RECT -180.230 -81.315 -180.060 -81.145 ;
        RECT -180.245 -81.755 -180.075 -81.585 ;
        RECT -175.270 -80.915 -175.100 -80.745 ;
        RECT -177.560 -81.315 -177.390 -81.145 ;
        RECT -172.585 -80.475 -172.415 -80.305 ;
        RECT -172.600 -80.915 -172.430 -80.745 ;
        RECT -165.365 -80.475 -165.195 -80.305 ;
        RECT -177.545 -81.755 -177.375 -81.585 ;
        RECT -170.310 -81.315 -170.140 -81.145 ;
        RECT -170.325 -81.755 -170.155 -81.585 ;
        RECT -165.350 -80.915 -165.180 -80.745 ;
        RECT -167.640 -81.315 -167.470 -81.145 ;
        RECT -162.665 -80.475 -162.495 -80.305 ;
        RECT -162.680 -80.915 -162.510 -80.745 ;
        RECT -155.445 -80.475 -155.275 -80.305 ;
        RECT -167.625 -81.755 -167.455 -81.585 ;
        RECT -160.390 -81.315 -160.220 -81.145 ;
        RECT -160.405 -81.755 -160.235 -81.585 ;
        RECT -155.430 -80.915 -155.260 -80.745 ;
        RECT -157.720 -81.315 -157.550 -81.145 ;
        RECT -152.745 -80.475 -152.575 -80.305 ;
        RECT -152.760 -80.915 -152.590 -80.745 ;
        RECT -145.525 -80.475 -145.355 -80.305 ;
        RECT -157.705 -81.755 -157.535 -81.585 ;
        RECT -150.470 -81.315 -150.300 -81.145 ;
        RECT -150.485 -81.755 -150.315 -81.585 ;
        RECT -145.510 -80.915 -145.340 -80.745 ;
        RECT -147.800 -81.315 -147.630 -81.145 ;
        RECT -142.825 -80.475 -142.655 -80.305 ;
        RECT -142.840 -80.915 -142.670 -80.745 ;
        RECT -135.605 -80.475 -135.435 -80.305 ;
        RECT -147.785 -81.755 -147.615 -81.585 ;
        RECT -140.550 -81.315 -140.380 -81.145 ;
        RECT -140.565 -81.755 -140.395 -81.585 ;
        RECT -135.590 -80.915 -135.420 -80.745 ;
        RECT -137.880 -81.315 -137.710 -81.145 ;
        RECT -132.905 -80.475 -132.735 -80.305 ;
        RECT -132.920 -80.915 -132.750 -80.745 ;
        RECT -125.685 -80.475 -125.515 -80.305 ;
        RECT -137.865 -81.755 -137.695 -81.585 ;
        RECT -130.630 -81.315 -130.460 -81.145 ;
        RECT -130.645 -81.755 -130.475 -81.585 ;
        RECT -125.670 -80.915 -125.500 -80.745 ;
        RECT -127.960 -81.315 -127.790 -81.145 ;
        RECT -122.985 -80.475 -122.815 -80.305 ;
        RECT -123.000 -80.915 -122.830 -80.745 ;
        RECT -115.765 -80.475 -115.595 -80.305 ;
        RECT -127.945 -81.755 -127.775 -81.585 ;
        RECT -120.710 -81.315 -120.540 -81.145 ;
        RECT -120.725 -81.755 -120.555 -81.585 ;
        RECT -115.750 -80.915 -115.580 -80.745 ;
        RECT -118.040 -81.315 -117.870 -81.145 ;
        RECT -113.065 -80.475 -112.895 -80.305 ;
        RECT -113.080 -80.915 -112.910 -80.745 ;
        RECT -105.845 -80.475 -105.675 -80.305 ;
        RECT -118.025 -81.755 -117.855 -81.585 ;
        RECT -110.790 -81.315 -110.620 -81.145 ;
        RECT -110.805 -81.755 -110.635 -81.585 ;
        RECT -105.830 -80.915 -105.660 -80.745 ;
        RECT -108.120 -81.315 -107.950 -81.145 ;
        RECT -103.145 -80.475 -102.975 -80.305 ;
        RECT -103.160 -80.915 -102.990 -80.745 ;
        RECT -95.925 -80.475 -95.755 -80.305 ;
        RECT -108.105 -81.755 -107.935 -81.585 ;
        RECT -100.870 -81.315 -100.700 -81.145 ;
        RECT -100.885 -81.755 -100.715 -81.585 ;
        RECT -95.910 -80.915 -95.740 -80.745 ;
        RECT -98.200 -81.315 -98.030 -81.145 ;
        RECT -93.225 -80.475 -93.055 -80.305 ;
        RECT -93.240 -80.915 -93.070 -80.745 ;
        RECT -86.005 -80.475 -85.835 -80.305 ;
        RECT -98.185 -81.755 -98.015 -81.585 ;
        RECT -90.950 -81.315 -90.780 -81.145 ;
        RECT -90.965 -81.755 -90.795 -81.585 ;
        RECT -85.990 -80.915 -85.820 -80.745 ;
        RECT -88.280 -81.315 -88.110 -81.145 ;
        RECT -83.305 -80.475 -83.135 -80.305 ;
        RECT -83.320 -80.915 -83.150 -80.745 ;
        RECT -76.085 -80.475 -75.915 -80.305 ;
        RECT -88.265 -81.755 -88.095 -81.585 ;
        RECT -81.030 -81.315 -80.860 -81.145 ;
        RECT -81.045 -81.755 -80.875 -81.585 ;
        RECT -76.070 -80.915 -75.900 -80.745 ;
        RECT -78.360 -81.315 -78.190 -81.145 ;
        RECT -73.385 -80.475 -73.215 -80.305 ;
        RECT -73.400 -80.915 -73.230 -80.745 ;
        RECT -66.165 -80.475 -65.995 -80.305 ;
        RECT -78.345 -81.755 -78.175 -81.585 ;
        RECT -71.110 -81.315 -70.940 -81.145 ;
        RECT -71.125 -81.755 -70.955 -81.585 ;
        RECT -66.150 -80.915 -65.980 -80.745 ;
        RECT -68.440 -81.315 -68.270 -81.145 ;
        RECT -63.465 -80.475 -63.295 -80.305 ;
        RECT -63.480 -80.915 -63.310 -80.745 ;
        RECT -56.245 -80.475 -56.075 -80.305 ;
        RECT -68.425 -81.755 -68.255 -81.585 ;
        RECT -61.190 -81.315 -61.020 -81.145 ;
        RECT -61.205 -81.755 -61.035 -81.585 ;
        RECT -56.230 -80.915 -56.060 -80.745 ;
        RECT -58.520 -81.315 -58.350 -81.145 ;
        RECT -53.545 -80.475 -53.375 -80.305 ;
        RECT -53.560 -80.915 -53.390 -80.745 ;
        RECT -46.325 -80.475 -46.155 -80.305 ;
        RECT -58.505 -81.755 -58.335 -81.585 ;
        RECT -51.270 -81.315 -51.100 -81.145 ;
        RECT -51.285 -81.755 -51.115 -81.585 ;
        RECT -46.310 -80.915 -46.140 -80.745 ;
        RECT -48.600 -81.315 -48.430 -81.145 ;
        RECT -43.625 -80.475 -43.455 -80.305 ;
        RECT -43.640 -80.915 -43.470 -80.745 ;
        RECT -36.405 -80.475 -36.235 -80.305 ;
        RECT -48.585 -81.755 -48.415 -81.585 ;
        RECT -41.350 -81.315 -41.180 -81.145 ;
        RECT -41.365 -81.755 -41.195 -81.585 ;
        RECT -36.390 -80.915 -36.220 -80.745 ;
        RECT -38.680 -81.315 -38.510 -81.145 ;
        RECT -33.705 -80.475 -33.535 -80.305 ;
        RECT -33.720 -80.915 -33.550 -80.745 ;
        RECT -26.485 -80.475 -26.315 -80.305 ;
        RECT -38.665 -81.755 -38.495 -81.585 ;
        RECT -31.430 -81.315 -31.260 -81.145 ;
        RECT -31.445 -81.755 -31.275 -81.585 ;
        RECT -26.470 -80.915 -26.300 -80.745 ;
        RECT -28.760 -81.315 -28.590 -81.145 ;
        RECT -23.785 -80.475 -23.615 -80.305 ;
        RECT -23.800 -80.915 -23.630 -80.745 ;
        RECT -16.565 -80.475 -16.395 -80.305 ;
        RECT -28.745 -81.755 -28.575 -81.585 ;
        RECT -21.510 -81.315 -21.340 -81.145 ;
        RECT -21.525 -81.755 -21.355 -81.585 ;
        RECT -16.550 -80.915 -16.380 -80.745 ;
        RECT -18.840 -81.315 -18.670 -81.145 ;
        RECT -13.865 -80.475 -13.695 -80.305 ;
        RECT -13.880 -80.915 -13.710 -80.745 ;
        RECT -6.645 -80.475 -6.475 -80.305 ;
        RECT -18.825 -81.755 -18.655 -81.585 ;
        RECT -11.590 -81.315 -11.420 -81.145 ;
        RECT -11.605 -81.755 -11.435 -81.585 ;
        RECT -6.630 -80.915 -6.460 -80.745 ;
        RECT -8.920 -81.315 -8.750 -81.145 ;
        RECT -3.945 -80.475 -3.775 -80.305 ;
        RECT -3.960 -80.915 -3.790 -80.745 ;
        RECT 3.275 -80.475 3.445 -80.305 ;
        RECT -8.905 -81.755 -8.735 -81.585 ;
        RECT -1.670 -81.315 -1.500 -81.145 ;
        RECT -1.685 -81.755 -1.515 -81.585 ;
        RECT 3.290 -80.915 3.460 -80.745 ;
        RECT 1.000 -81.315 1.170 -81.145 ;
        RECT 5.975 -80.475 6.145 -80.305 ;
        RECT 5.960 -80.915 6.130 -80.745 ;
        RECT 13.195 -80.475 13.365 -80.305 ;
        RECT 1.015 -81.755 1.185 -81.585 ;
        RECT 8.250 -81.315 8.420 -81.145 ;
        RECT 8.235 -81.755 8.405 -81.585 ;
        RECT 13.210 -80.915 13.380 -80.745 ;
        RECT 10.920 -81.315 11.090 -81.145 ;
        RECT 15.895 -80.475 16.065 -80.305 ;
        RECT 15.880 -80.915 16.050 -80.745 ;
        RECT 23.115 -80.475 23.285 -80.305 ;
        RECT 10.935 -81.755 11.105 -81.585 ;
        RECT 18.170 -81.315 18.340 -81.145 ;
        RECT 18.155 -81.755 18.325 -81.585 ;
        RECT 23.130 -80.915 23.300 -80.745 ;
        RECT 20.840 -81.315 21.010 -81.145 ;
        RECT 20.855 -81.755 21.025 -81.585 ;
        RECT -292.975 -82.475 -292.805 -82.305 ;
        RECT -292.515 -82.475 -292.345 -82.305 ;
        RECT -292.055 -82.475 -291.885 -82.305 ;
        RECT -291.595 -82.475 -291.425 -82.305 ;
        RECT -291.205 -83.135 -291.035 -82.965 ;
        RECT -291.205 -83.595 -291.035 -83.425 ;
        RECT -290.045 -83.175 -289.875 -83.005 ;
        RECT -285.985 -83.175 -285.815 -83.005 ;
        RECT -280.125 -83.175 -279.955 -83.005 ;
        RECT -276.065 -83.175 -275.895 -83.005 ;
        RECT -270.205 -83.175 -270.035 -83.005 ;
        RECT -266.145 -83.175 -265.975 -83.005 ;
        RECT -260.285 -83.175 -260.115 -83.005 ;
        RECT -256.225 -83.175 -256.055 -83.005 ;
        RECT -250.365 -83.175 -250.195 -83.005 ;
        RECT -246.305 -83.175 -246.135 -83.005 ;
        RECT -240.445 -83.175 -240.275 -83.005 ;
        RECT -236.385 -83.175 -236.215 -83.005 ;
        RECT -230.525 -83.175 -230.355 -83.005 ;
        RECT -226.465 -83.175 -226.295 -83.005 ;
        RECT -220.605 -83.175 -220.435 -83.005 ;
        RECT -216.545 -83.175 -216.375 -83.005 ;
        RECT -210.685 -83.175 -210.515 -83.005 ;
        RECT -206.625 -83.175 -206.455 -83.005 ;
        RECT -200.765 -83.175 -200.595 -83.005 ;
        RECT -196.705 -83.175 -196.535 -83.005 ;
        RECT -190.845 -83.175 -190.675 -83.005 ;
        RECT -186.785 -83.175 -186.615 -83.005 ;
        RECT -180.925 -83.175 -180.755 -83.005 ;
        RECT -176.865 -83.175 -176.695 -83.005 ;
        RECT -171.005 -83.175 -170.835 -83.005 ;
        RECT -166.945 -83.175 -166.775 -83.005 ;
        RECT -161.085 -83.175 -160.915 -83.005 ;
        RECT -157.025 -83.175 -156.855 -83.005 ;
        RECT -151.165 -83.175 -150.995 -83.005 ;
        RECT -147.105 -83.175 -146.935 -83.005 ;
        RECT -141.245 -83.175 -141.075 -83.005 ;
        RECT -137.185 -83.175 -137.015 -83.005 ;
        RECT -131.325 -83.175 -131.155 -83.005 ;
        RECT -127.265 -83.175 -127.095 -83.005 ;
        RECT -121.405 -83.175 -121.235 -83.005 ;
        RECT -117.345 -83.175 -117.175 -83.005 ;
        RECT -111.485 -83.175 -111.315 -83.005 ;
        RECT -107.425 -83.175 -107.255 -83.005 ;
        RECT -101.565 -83.175 -101.395 -83.005 ;
        RECT -97.505 -83.175 -97.335 -83.005 ;
        RECT -91.645 -83.175 -91.475 -83.005 ;
        RECT -87.585 -83.175 -87.415 -83.005 ;
        RECT -81.725 -83.175 -81.555 -83.005 ;
        RECT -77.665 -83.175 -77.495 -83.005 ;
        RECT -71.805 -83.175 -71.635 -83.005 ;
        RECT -67.745 -83.175 -67.575 -83.005 ;
        RECT -61.885 -83.175 -61.715 -83.005 ;
        RECT -57.825 -83.175 -57.655 -83.005 ;
        RECT -51.965 -83.175 -51.795 -83.005 ;
        RECT -47.905 -83.175 -47.735 -83.005 ;
        RECT -42.045 -83.175 -41.875 -83.005 ;
        RECT -37.985 -83.175 -37.815 -83.005 ;
        RECT -32.125 -83.175 -31.955 -83.005 ;
        RECT -28.065 -83.175 -27.895 -83.005 ;
        RECT -22.205 -83.175 -22.035 -83.005 ;
        RECT -18.145 -83.175 -17.975 -83.005 ;
        RECT -12.285 -83.175 -12.115 -83.005 ;
        RECT -8.225 -83.175 -8.055 -83.005 ;
        RECT -2.365 -83.175 -2.195 -83.005 ;
        RECT 1.695 -83.175 1.865 -83.005 ;
        RECT 7.555 -83.175 7.725 -83.005 ;
        RECT 11.615 -83.175 11.785 -83.005 ;
        RECT 17.475 -83.175 17.645 -83.005 ;
        RECT 21.535 -83.175 21.705 -83.005 ;
        RECT 22.695 -83.135 22.865 -82.965 ;
        RECT 22.695 -83.595 22.865 -83.425 ;
        RECT -291.675 -84.045 -291.505 -83.875 ;
        RECT -291.205 -84.055 -291.035 -83.885 ;
        RECT -286.720 -84.025 -286.550 -83.855 ;
        RECT -285.355 -84.025 -285.185 -83.855 ;
        RECT -276.800 -84.025 -276.630 -83.855 ;
        RECT -275.435 -84.025 -275.265 -83.855 ;
        RECT -266.880 -84.025 -266.710 -83.855 ;
        RECT -265.515 -84.025 -265.345 -83.855 ;
        RECT -256.960 -84.025 -256.790 -83.855 ;
        RECT -255.595 -84.025 -255.425 -83.855 ;
        RECT -247.040 -84.025 -246.870 -83.855 ;
        RECT -245.675 -84.025 -245.505 -83.855 ;
        RECT -237.120 -84.025 -236.950 -83.855 ;
        RECT -235.755 -84.025 -235.585 -83.855 ;
        RECT -227.200 -84.025 -227.030 -83.855 ;
        RECT -225.835 -84.025 -225.665 -83.855 ;
        RECT -217.280 -84.025 -217.110 -83.855 ;
        RECT -215.915 -84.025 -215.745 -83.855 ;
        RECT -207.360 -84.025 -207.190 -83.855 ;
        RECT -205.995 -84.025 -205.825 -83.855 ;
        RECT -197.440 -84.025 -197.270 -83.855 ;
        RECT -196.075 -84.025 -195.905 -83.855 ;
        RECT -187.520 -84.025 -187.350 -83.855 ;
        RECT -186.155 -84.025 -185.985 -83.855 ;
        RECT -177.600 -84.025 -177.430 -83.855 ;
        RECT -176.235 -84.025 -176.065 -83.855 ;
        RECT -167.680 -84.025 -167.510 -83.855 ;
        RECT -166.315 -84.025 -166.145 -83.855 ;
        RECT -157.760 -84.025 -157.590 -83.855 ;
        RECT -156.395 -84.025 -156.225 -83.855 ;
        RECT -147.840 -84.025 -147.670 -83.855 ;
        RECT -146.475 -84.025 -146.305 -83.855 ;
        RECT -137.920 -84.025 -137.750 -83.855 ;
        RECT -136.555 -84.025 -136.385 -83.855 ;
        RECT -128.000 -84.025 -127.830 -83.855 ;
        RECT -126.635 -84.025 -126.465 -83.855 ;
        RECT -118.080 -84.025 -117.910 -83.855 ;
        RECT -116.715 -84.025 -116.545 -83.855 ;
        RECT -108.160 -84.025 -107.990 -83.855 ;
        RECT -106.795 -84.025 -106.625 -83.855 ;
        RECT -98.240 -84.025 -98.070 -83.855 ;
        RECT -96.875 -84.025 -96.705 -83.855 ;
        RECT -88.320 -84.025 -88.150 -83.855 ;
        RECT -86.955 -84.025 -86.785 -83.855 ;
        RECT -78.400 -84.025 -78.230 -83.855 ;
        RECT -77.035 -84.025 -76.865 -83.855 ;
        RECT -68.480 -84.025 -68.310 -83.855 ;
        RECT -67.115 -84.025 -66.945 -83.855 ;
        RECT -58.560 -84.025 -58.390 -83.855 ;
        RECT -57.195 -84.025 -57.025 -83.855 ;
        RECT -48.640 -84.025 -48.470 -83.855 ;
        RECT -47.275 -84.025 -47.105 -83.855 ;
        RECT -38.720 -84.025 -38.550 -83.855 ;
        RECT -37.355 -84.025 -37.185 -83.855 ;
        RECT -28.800 -84.025 -28.630 -83.855 ;
        RECT -27.435 -84.025 -27.265 -83.855 ;
        RECT -18.880 -84.025 -18.710 -83.855 ;
        RECT -17.515 -84.025 -17.345 -83.855 ;
        RECT -8.960 -84.025 -8.790 -83.855 ;
        RECT -7.595 -84.025 -7.425 -83.855 ;
        RECT 0.960 -84.025 1.130 -83.855 ;
        RECT 2.325 -84.025 2.495 -83.855 ;
        RECT 10.880 -84.025 11.050 -83.855 ;
        RECT 12.245 -84.025 12.415 -83.855 ;
        RECT 20.800 -84.025 20.970 -83.855 ;
        RECT 22.165 -84.025 22.335 -83.855 ;
        RECT 22.695 -84.055 22.865 -83.885 ;
        RECT 23.165 -84.045 23.335 -83.875 ;
        RECT -294.735 -172.760 -294.565 -172.590 ;
        RECT -294.265 -172.755 -294.095 -172.585 ;
        RECT -293.440 -172.785 -293.270 -172.615 ;
        RECT -292.075 -172.785 -291.905 -172.615 ;
        RECT -283.520 -172.785 -283.350 -172.615 ;
        RECT -282.155 -172.785 -281.985 -172.615 ;
        RECT -273.600 -172.785 -273.430 -172.615 ;
        RECT -272.235 -172.785 -272.065 -172.615 ;
        RECT -263.680 -172.785 -263.510 -172.615 ;
        RECT -262.315 -172.785 -262.145 -172.615 ;
        RECT -253.760 -172.785 -253.590 -172.615 ;
        RECT -252.395 -172.785 -252.225 -172.615 ;
        RECT -243.840 -172.785 -243.670 -172.615 ;
        RECT -242.475 -172.785 -242.305 -172.615 ;
        RECT -233.920 -172.785 -233.750 -172.615 ;
        RECT -232.555 -172.785 -232.385 -172.615 ;
        RECT -224.000 -172.785 -223.830 -172.615 ;
        RECT -222.635 -172.785 -222.465 -172.615 ;
        RECT -214.080 -172.785 -213.910 -172.615 ;
        RECT -212.715 -172.785 -212.545 -172.615 ;
        RECT -204.160 -172.785 -203.990 -172.615 ;
        RECT -202.795 -172.785 -202.625 -172.615 ;
        RECT -194.240 -172.785 -194.070 -172.615 ;
        RECT -192.875 -172.785 -192.705 -172.615 ;
        RECT -184.320 -172.785 -184.150 -172.615 ;
        RECT -182.955 -172.785 -182.785 -172.615 ;
        RECT -174.400 -172.785 -174.230 -172.615 ;
        RECT -173.035 -172.785 -172.865 -172.615 ;
        RECT -164.480 -172.785 -164.310 -172.615 ;
        RECT -163.115 -172.785 -162.945 -172.615 ;
        RECT -154.560 -172.785 -154.390 -172.615 ;
        RECT -153.195 -172.785 -153.025 -172.615 ;
        RECT -144.640 -172.785 -144.470 -172.615 ;
        RECT -143.275 -172.785 -143.105 -172.615 ;
        RECT -134.720 -172.785 -134.550 -172.615 ;
        RECT -133.355 -172.785 -133.185 -172.615 ;
        RECT -124.800 -172.785 -124.630 -172.615 ;
        RECT -123.435 -172.785 -123.265 -172.615 ;
        RECT -114.880 -172.785 -114.710 -172.615 ;
        RECT -113.515 -172.785 -113.345 -172.615 ;
        RECT -104.960 -172.785 -104.790 -172.615 ;
        RECT -103.595 -172.785 -103.425 -172.615 ;
        RECT -95.040 -172.785 -94.870 -172.615 ;
        RECT -93.675 -172.785 -93.505 -172.615 ;
        RECT -85.120 -172.785 -84.950 -172.615 ;
        RECT -83.755 -172.785 -83.585 -172.615 ;
        RECT -75.200 -172.785 -75.030 -172.615 ;
        RECT -73.835 -172.785 -73.665 -172.615 ;
        RECT -65.280 -172.785 -65.110 -172.615 ;
        RECT -63.915 -172.785 -63.745 -172.615 ;
        RECT -55.360 -172.785 -55.190 -172.615 ;
        RECT -53.995 -172.785 -53.825 -172.615 ;
        RECT -45.440 -172.785 -45.270 -172.615 ;
        RECT -44.075 -172.785 -43.905 -172.615 ;
        RECT -35.520 -172.785 -35.350 -172.615 ;
        RECT -34.155 -172.785 -33.985 -172.615 ;
        RECT -25.600 -172.785 -25.430 -172.615 ;
        RECT -24.235 -172.785 -24.065 -172.615 ;
        RECT -15.680 -172.785 -15.510 -172.615 ;
        RECT -14.315 -172.785 -14.145 -172.615 ;
        RECT -5.760 -172.785 -5.590 -172.615 ;
        RECT -4.395 -172.785 -4.225 -172.615 ;
        RECT 4.160 -172.785 4.330 -172.615 ;
        RECT 5.525 -172.785 5.695 -172.615 ;
        RECT 14.080 -172.785 14.250 -172.615 ;
        RECT 15.445 -172.785 15.615 -172.615 ;
        RECT -294.265 -173.215 -294.095 -173.045 ;
        RECT -294.265 -173.675 -294.095 -173.505 ;
        RECT -292.705 -173.635 -292.535 -173.465 ;
        RECT -286.845 -173.635 -286.675 -173.465 ;
        RECT -282.785 -173.635 -282.615 -173.465 ;
        RECT -276.925 -173.635 -276.755 -173.465 ;
        RECT -272.865 -173.635 -272.695 -173.465 ;
        RECT -267.005 -173.635 -266.835 -173.465 ;
        RECT -262.945 -173.635 -262.775 -173.465 ;
        RECT -257.085 -173.635 -256.915 -173.465 ;
        RECT -253.025 -173.635 -252.855 -173.465 ;
        RECT -247.165 -173.635 -246.995 -173.465 ;
        RECT -243.105 -173.635 -242.935 -173.465 ;
        RECT -237.245 -173.635 -237.075 -173.465 ;
        RECT -233.185 -173.635 -233.015 -173.465 ;
        RECT -227.325 -173.635 -227.155 -173.465 ;
        RECT -223.265 -173.635 -223.095 -173.465 ;
        RECT -217.405 -173.635 -217.235 -173.465 ;
        RECT -213.345 -173.635 -213.175 -173.465 ;
        RECT -207.485 -173.635 -207.315 -173.465 ;
        RECT -203.425 -173.635 -203.255 -173.465 ;
        RECT -197.565 -173.635 -197.395 -173.465 ;
        RECT -193.505 -173.635 -193.335 -173.465 ;
        RECT -187.645 -173.635 -187.475 -173.465 ;
        RECT -183.585 -173.635 -183.415 -173.465 ;
        RECT -177.725 -173.635 -177.555 -173.465 ;
        RECT -173.665 -173.635 -173.495 -173.465 ;
        RECT -167.805 -173.635 -167.635 -173.465 ;
        RECT -163.745 -173.635 -163.575 -173.465 ;
        RECT -157.885 -173.635 -157.715 -173.465 ;
        RECT -153.825 -173.635 -153.655 -173.465 ;
        RECT -147.965 -173.635 -147.795 -173.465 ;
        RECT -143.905 -173.635 -143.735 -173.465 ;
        RECT -138.045 -173.635 -137.875 -173.465 ;
        RECT -133.985 -173.635 -133.815 -173.465 ;
        RECT -128.125 -173.635 -127.955 -173.465 ;
        RECT -124.065 -173.635 -123.895 -173.465 ;
        RECT -118.205 -173.635 -118.035 -173.465 ;
        RECT -114.145 -173.635 -113.975 -173.465 ;
        RECT -108.285 -173.635 -108.115 -173.465 ;
        RECT -104.225 -173.635 -104.055 -173.465 ;
        RECT -98.365 -173.635 -98.195 -173.465 ;
        RECT -94.305 -173.635 -94.135 -173.465 ;
        RECT -88.445 -173.635 -88.275 -173.465 ;
        RECT -84.385 -173.635 -84.215 -173.465 ;
        RECT -78.525 -173.635 -78.355 -173.465 ;
        RECT -74.465 -173.635 -74.295 -173.465 ;
        RECT -68.605 -173.635 -68.435 -173.465 ;
        RECT -64.545 -173.635 -64.375 -173.465 ;
        RECT -58.685 -173.635 -58.515 -173.465 ;
        RECT -54.625 -173.635 -54.455 -173.465 ;
        RECT -48.765 -173.635 -48.595 -173.465 ;
        RECT -44.705 -173.635 -44.535 -173.465 ;
        RECT -38.845 -173.635 -38.675 -173.465 ;
        RECT -34.785 -173.635 -34.615 -173.465 ;
        RECT -28.925 -173.635 -28.755 -173.465 ;
        RECT -24.865 -173.635 -24.695 -173.465 ;
        RECT -19.005 -173.635 -18.835 -173.465 ;
        RECT -14.945 -173.635 -14.775 -173.465 ;
        RECT -9.085 -173.635 -8.915 -173.465 ;
        RECT -5.025 -173.635 -4.855 -173.465 ;
        RECT 0.835 -173.635 1.005 -173.465 ;
        RECT 4.895 -173.635 5.065 -173.465 ;
        RECT 10.755 -173.635 10.925 -173.465 ;
        RECT 14.815 -173.635 14.985 -173.465 ;
        RECT 20.675 -173.635 20.845 -173.465 ;
        RECT -294.735 -174.335 -294.565 -174.165 ;
        RECT -294.275 -174.335 -294.105 -174.165 ;
        RECT -293.815 -174.335 -293.645 -174.165 ;
        RECT -293.355 -174.335 -293.185 -174.165 ;
        RECT 21.325 -174.335 21.495 -174.165 ;
        RECT 21.785 -174.335 21.955 -174.165 ;
        RECT 22.245 -174.335 22.415 -174.165 ;
        RECT 22.705 -174.335 22.875 -174.165 ;
        RECT -293.385 -175.055 -293.215 -174.885 ;
        RECT -293.400 -175.495 -293.230 -175.325 ;
        RECT -286.165 -175.055 -285.995 -174.885 ;
        RECT -291.110 -175.895 -290.940 -175.725 ;
        RECT -291.125 -176.335 -290.955 -176.165 ;
        RECT -286.150 -175.495 -285.980 -175.325 ;
        RECT -288.440 -175.895 -288.270 -175.725 ;
        RECT -283.465 -175.055 -283.295 -174.885 ;
        RECT -283.480 -175.495 -283.310 -175.325 ;
        RECT -276.245 -175.055 -276.075 -174.885 ;
        RECT -288.425 -176.335 -288.255 -176.165 ;
        RECT -281.190 -175.895 -281.020 -175.725 ;
        RECT -281.205 -176.335 -281.035 -176.165 ;
        RECT -276.230 -175.495 -276.060 -175.325 ;
        RECT -278.520 -175.895 -278.350 -175.725 ;
        RECT -273.545 -175.055 -273.375 -174.885 ;
        RECT -273.560 -175.495 -273.390 -175.325 ;
        RECT -266.325 -175.055 -266.155 -174.885 ;
        RECT -278.505 -176.335 -278.335 -176.165 ;
        RECT -271.270 -175.895 -271.100 -175.725 ;
        RECT -271.285 -176.335 -271.115 -176.165 ;
        RECT -266.310 -175.495 -266.140 -175.325 ;
        RECT -268.600 -175.895 -268.430 -175.725 ;
        RECT -263.625 -175.055 -263.455 -174.885 ;
        RECT -263.640 -175.495 -263.470 -175.325 ;
        RECT -256.405 -175.055 -256.235 -174.885 ;
        RECT -268.585 -176.335 -268.415 -176.165 ;
        RECT -261.350 -175.895 -261.180 -175.725 ;
        RECT -261.365 -176.335 -261.195 -176.165 ;
        RECT -256.390 -175.495 -256.220 -175.325 ;
        RECT -258.680 -175.895 -258.510 -175.725 ;
        RECT -253.705 -175.055 -253.535 -174.885 ;
        RECT -253.720 -175.495 -253.550 -175.325 ;
        RECT -246.485 -175.055 -246.315 -174.885 ;
        RECT -258.665 -176.335 -258.495 -176.165 ;
        RECT -251.430 -175.895 -251.260 -175.725 ;
        RECT -251.445 -176.335 -251.275 -176.165 ;
        RECT -246.470 -175.495 -246.300 -175.325 ;
        RECT -248.760 -175.895 -248.590 -175.725 ;
        RECT -243.785 -175.055 -243.615 -174.885 ;
        RECT -243.800 -175.495 -243.630 -175.325 ;
        RECT -236.565 -175.055 -236.395 -174.885 ;
        RECT -248.745 -176.335 -248.575 -176.165 ;
        RECT -241.510 -175.895 -241.340 -175.725 ;
        RECT -241.525 -176.335 -241.355 -176.165 ;
        RECT -236.550 -175.495 -236.380 -175.325 ;
        RECT -238.840 -175.895 -238.670 -175.725 ;
        RECT -233.865 -175.055 -233.695 -174.885 ;
        RECT -233.880 -175.495 -233.710 -175.325 ;
        RECT -226.645 -175.055 -226.475 -174.885 ;
        RECT -238.825 -176.335 -238.655 -176.165 ;
        RECT -231.590 -175.895 -231.420 -175.725 ;
        RECT -231.605 -176.335 -231.435 -176.165 ;
        RECT -226.630 -175.495 -226.460 -175.325 ;
        RECT -228.920 -175.895 -228.750 -175.725 ;
        RECT -223.945 -175.055 -223.775 -174.885 ;
        RECT -223.960 -175.495 -223.790 -175.325 ;
        RECT -216.725 -175.055 -216.555 -174.885 ;
        RECT -228.905 -176.335 -228.735 -176.165 ;
        RECT -221.670 -175.895 -221.500 -175.725 ;
        RECT -221.685 -176.335 -221.515 -176.165 ;
        RECT -216.710 -175.495 -216.540 -175.325 ;
        RECT -219.000 -175.895 -218.830 -175.725 ;
        RECT -214.025 -175.055 -213.855 -174.885 ;
        RECT -214.040 -175.495 -213.870 -175.325 ;
        RECT -206.805 -175.055 -206.635 -174.885 ;
        RECT -218.985 -176.335 -218.815 -176.165 ;
        RECT -211.750 -175.895 -211.580 -175.725 ;
        RECT -211.765 -176.335 -211.595 -176.165 ;
        RECT -206.790 -175.495 -206.620 -175.325 ;
        RECT -209.080 -175.895 -208.910 -175.725 ;
        RECT -204.105 -175.055 -203.935 -174.885 ;
        RECT -204.120 -175.495 -203.950 -175.325 ;
        RECT -196.885 -175.055 -196.715 -174.885 ;
        RECT -209.065 -176.335 -208.895 -176.165 ;
        RECT -201.830 -175.895 -201.660 -175.725 ;
        RECT -201.845 -176.335 -201.675 -176.165 ;
        RECT -196.870 -175.495 -196.700 -175.325 ;
        RECT -199.160 -175.895 -198.990 -175.725 ;
        RECT -194.185 -175.055 -194.015 -174.885 ;
        RECT -194.200 -175.495 -194.030 -175.325 ;
        RECT -186.965 -175.055 -186.795 -174.885 ;
        RECT -199.145 -176.335 -198.975 -176.165 ;
        RECT -191.910 -175.895 -191.740 -175.725 ;
        RECT -191.925 -176.335 -191.755 -176.165 ;
        RECT -186.950 -175.495 -186.780 -175.325 ;
        RECT -189.240 -175.895 -189.070 -175.725 ;
        RECT -184.265 -175.055 -184.095 -174.885 ;
        RECT -184.280 -175.495 -184.110 -175.325 ;
        RECT -177.045 -175.055 -176.875 -174.885 ;
        RECT -189.225 -176.335 -189.055 -176.165 ;
        RECT -181.990 -175.895 -181.820 -175.725 ;
        RECT -182.005 -176.335 -181.835 -176.165 ;
        RECT -177.030 -175.495 -176.860 -175.325 ;
        RECT -179.320 -175.895 -179.150 -175.725 ;
        RECT -174.345 -175.055 -174.175 -174.885 ;
        RECT -174.360 -175.495 -174.190 -175.325 ;
        RECT -167.125 -175.055 -166.955 -174.885 ;
        RECT -179.305 -176.335 -179.135 -176.165 ;
        RECT -172.070 -175.895 -171.900 -175.725 ;
        RECT -172.085 -176.335 -171.915 -176.165 ;
        RECT -167.110 -175.495 -166.940 -175.325 ;
        RECT -169.400 -175.895 -169.230 -175.725 ;
        RECT -164.425 -175.055 -164.255 -174.885 ;
        RECT -164.440 -175.495 -164.270 -175.325 ;
        RECT -157.205 -175.055 -157.035 -174.885 ;
        RECT -169.385 -176.335 -169.215 -176.165 ;
        RECT -162.150 -175.895 -161.980 -175.725 ;
        RECT -162.165 -176.335 -161.995 -176.165 ;
        RECT -157.190 -175.495 -157.020 -175.325 ;
        RECT -159.480 -175.895 -159.310 -175.725 ;
        RECT -154.505 -175.055 -154.335 -174.885 ;
        RECT -154.520 -175.495 -154.350 -175.325 ;
        RECT -147.285 -175.055 -147.115 -174.885 ;
        RECT -159.465 -176.335 -159.295 -176.165 ;
        RECT -152.230 -175.895 -152.060 -175.725 ;
        RECT -152.245 -176.335 -152.075 -176.165 ;
        RECT -147.270 -175.495 -147.100 -175.325 ;
        RECT -149.560 -175.895 -149.390 -175.725 ;
        RECT -144.585 -175.055 -144.415 -174.885 ;
        RECT -144.600 -175.495 -144.430 -175.325 ;
        RECT -137.365 -175.055 -137.195 -174.885 ;
        RECT -149.545 -176.335 -149.375 -176.165 ;
        RECT -142.310 -175.895 -142.140 -175.725 ;
        RECT -142.325 -176.335 -142.155 -176.165 ;
        RECT -137.350 -175.495 -137.180 -175.325 ;
        RECT -139.640 -175.895 -139.470 -175.725 ;
        RECT -134.665 -175.055 -134.495 -174.885 ;
        RECT -134.680 -175.495 -134.510 -175.325 ;
        RECT -127.445 -175.055 -127.275 -174.885 ;
        RECT -139.625 -176.335 -139.455 -176.165 ;
        RECT -132.390 -175.895 -132.220 -175.725 ;
        RECT -132.405 -176.335 -132.235 -176.165 ;
        RECT -127.430 -175.495 -127.260 -175.325 ;
        RECT -129.720 -175.895 -129.550 -175.725 ;
        RECT -124.745 -175.055 -124.575 -174.885 ;
        RECT -124.760 -175.495 -124.590 -175.325 ;
        RECT -117.525 -175.055 -117.355 -174.885 ;
        RECT -129.705 -176.335 -129.535 -176.165 ;
        RECT -122.470 -175.895 -122.300 -175.725 ;
        RECT -122.485 -176.335 -122.315 -176.165 ;
        RECT -117.510 -175.495 -117.340 -175.325 ;
        RECT -119.800 -175.895 -119.630 -175.725 ;
        RECT -114.825 -175.055 -114.655 -174.885 ;
        RECT -114.840 -175.495 -114.670 -175.325 ;
        RECT -107.605 -175.055 -107.435 -174.885 ;
        RECT -119.785 -176.335 -119.615 -176.165 ;
        RECT -112.550 -175.895 -112.380 -175.725 ;
        RECT -112.565 -176.335 -112.395 -176.165 ;
        RECT -107.590 -175.495 -107.420 -175.325 ;
        RECT -109.880 -175.895 -109.710 -175.725 ;
        RECT -104.905 -175.055 -104.735 -174.885 ;
        RECT -104.920 -175.495 -104.750 -175.325 ;
        RECT -97.685 -175.055 -97.515 -174.885 ;
        RECT -109.865 -176.335 -109.695 -176.165 ;
        RECT -102.630 -175.895 -102.460 -175.725 ;
        RECT -102.645 -176.335 -102.475 -176.165 ;
        RECT -97.670 -175.495 -97.500 -175.325 ;
        RECT -99.960 -175.895 -99.790 -175.725 ;
        RECT -94.985 -175.055 -94.815 -174.885 ;
        RECT -95.000 -175.495 -94.830 -175.325 ;
        RECT -87.765 -175.055 -87.595 -174.885 ;
        RECT -99.945 -176.335 -99.775 -176.165 ;
        RECT -92.710 -175.895 -92.540 -175.725 ;
        RECT -92.725 -176.335 -92.555 -176.165 ;
        RECT -87.750 -175.495 -87.580 -175.325 ;
        RECT -90.040 -175.895 -89.870 -175.725 ;
        RECT -85.065 -175.055 -84.895 -174.885 ;
        RECT -85.080 -175.495 -84.910 -175.325 ;
        RECT -77.845 -175.055 -77.675 -174.885 ;
        RECT -90.025 -176.335 -89.855 -176.165 ;
        RECT -82.790 -175.895 -82.620 -175.725 ;
        RECT -82.805 -176.335 -82.635 -176.165 ;
        RECT -77.830 -175.495 -77.660 -175.325 ;
        RECT -80.120 -175.895 -79.950 -175.725 ;
        RECT -75.145 -175.055 -74.975 -174.885 ;
        RECT -75.160 -175.495 -74.990 -175.325 ;
        RECT -67.925 -175.055 -67.755 -174.885 ;
        RECT -80.105 -176.335 -79.935 -176.165 ;
        RECT -72.870 -175.895 -72.700 -175.725 ;
        RECT -72.885 -176.335 -72.715 -176.165 ;
        RECT -67.910 -175.495 -67.740 -175.325 ;
        RECT -70.200 -175.895 -70.030 -175.725 ;
        RECT -65.225 -175.055 -65.055 -174.885 ;
        RECT -65.240 -175.495 -65.070 -175.325 ;
        RECT -58.005 -175.055 -57.835 -174.885 ;
        RECT -70.185 -176.335 -70.015 -176.165 ;
        RECT -62.950 -175.895 -62.780 -175.725 ;
        RECT -62.965 -176.335 -62.795 -176.165 ;
        RECT -57.990 -175.495 -57.820 -175.325 ;
        RECT -60.280 -175.895 -60.110 -175.725 ;
        RECT -55.305 -175.055 -55.135 -174.885 ;
        RECT -55.320 -175.495 -55.150 -175.325 ;
        RECT -48.085 -175.055 -47.915 -174.885 ;
        RECT -60.265 -176.335 -60.095 -176.165 ;
        RECT -53.030 -175.895 -52.860 -175.725 ;
        RECT -53.045 -176.335 -52.875 -176.165 ;
        RECT -48.070 -175.495 -47.900 -175.325 ;
        RECT -50.360 -175.895 -50.190 -175.725 ;
        RECT -45.385 -175.055 -45.215 -174.885 ;
        RECT -45.400 -175.495 -45.230 -175.325 ;
        RECT -38.165 -175.055 -37.995 -174.885 ;
        RECT -50.345 -176.335 -50.175 -176.165 ;
        RECT -43.110 -175.895 -42.940 -175.725 ;
        RECT -43.125 -176.335 -42.955 -176.165 ;
        RECT -38.150 -175.495 -37.980 -175.325 ;
        RECT -40.440 -175.895 -40.270 -175.725 ;
        RECT -35.465 -175.055 -35.295 -174.885 ;
        RECT -35.480 -175.495 -35.310 -175.325 ;
        RECT -28.245 -175.055 -28.075 -174.885 ;
        RECT -40.425 -176.335 -40.255 -176.165 ;
        RECT -33.190 -175.895 -33.020 -175.725 ;
        RECT -33.205 -176.335 -33.035 -176.165 ;
        RECT -28.230 -175.495 -28.060 -175.325 ;
        RECT -30.520 -175.895 -30.350 -175.725 ;
        RECT -25.545 -175.055 -25.375 -174.885 ;
        RECT -25.560 -175.495 -25.390 -175.325 ;
        RECT -18.325 -175.055 -18.155 -174.885 ;
        RECT -30.505 -176.335 -30.335 -176.165 ;
        RECT -23.270 -175.895 -23.100 -175.725 ;
        RECT -23.285 -176.335 -23.115 -176.165 ;
        RECT -18.310 -175.495 -18.140 -175.325 ;
        RECT -20.600 -175.895 -20.430 -175.725 ;
        RECT -15.625 -175.055 -15.455 -174.885 ;
        RECT -15.640 -175.495 -15.470 -175.325 ;
        RECT -8.405 -175.055 -8.235 -174.885 ;
        RECT -20.585 -176.335 -20.415 -176.165 ;
        RECT -13.350 -175.895 -13.180 -175.725 ;
        RECT -13.365 -176.335 -13.195 -176.165 ;
        RECT -8.390 -175.495 -8.220 -175.325 ;
        RECT -10.680 -175.895 -10.510 -175.725 ;
        RECT -5.705 -175.055 -5.535 -174.885 ;
        RECT -5.720 -175.495 -5.550 -175.325 ;
        RECT 1.515 -175.055 1.685 -174.885 ;
        RECT -10.665 -176.335 -10.495 -176.165 ;
        RECT -3.430 -175.895 -3.260 -175.725 ;
        RECT -3.445 -176.335 -3.275 -176.165 ;
        RECT 1.530 -175.495 1.700 -175.325 ;
        RECT -0.760 -175.895 -0.590 -175.725 ;
        RECT 4.215 -175.055 4.385 -174.885 ;
        RECT 4.200 -175.495 4.370 -175.325 ;
        RECT 11.435 -175.055 11.605 -174.885 ;
        RECT -0.745 -176.335 -0.575 -176.165 ;
        RECT 6.490 -175.895 6.660 -175.725 ;
        RECT 6.475 -176.335 6.645 -176.165 ;
        RECT 11.450 -175.495 11.620 -175.325 ;
        RECT 9.160 -175.895 9.330 -175.725 ;
        RECT 14.135 -175.055 14.305 -174.885 ;
        RECT 14.120 -175.495 14.290 -175.325 ;
        RECT 21.355 -175.055 21.525 -174.885 ;
        RECT 9.175 -176.335 9.345 -176.165 ;
        RECT 16.410 -175.895 16.580 -175.725 ;
        RECT 16.395 -176.335 16.565 -176.165 ;
        RECT 21.370 -175.495 21.540 -175.325 ;
        RECT 19.080 -175.895 19.250 -175.725 ;
        RECT 19.095 -176.335 19.265 -176.165 ;
        RECT -294.735 -177.055 -294.565 -176.885 ;
        RECT -294.275 -177.055 -294.105 -176.885 ;
        RECT -293.815 -177.055 -293.645 -176.885 ;
        RECT -293.355 -177.055 -293.185 -176.885 ;
        RECT -292.965 -177.715 -292.795 -177.545 ;
        RECT -292.965 -178.175 -292.795 -178.005 ;
        RECT -291.805 -177.755 -291.635 -177.585 ;
        RECT -287.745 -177.755 -287.575 -177.585 ;
        RECT -281.885 -177.755 -281.715 -177.585 ;
        RECT -277.825 -177.755 -277.655 -177.585 ;
        RECT -271.965 -177.755 -271.795 -177.585 ;
        RECT -267.905 -177.755 -267.735 -177.585 ;
        RECT -262.045 -177.755 -261.875 -177.585 ;
        RECT -257.985 -177.755 -257.815 -177.585 ;
        RECT -252.125 -177.755 -251.955 -177.585 ;
        RECT -248.065 -177.755 -247.895 -177.585 ;
        RECT -242.205 -177.755 -242.035 -177.585 ;
        RECT -238.145 -177.755 -237.975 -177.585 ;
        RECT -232.285 -177.755 -232.115 -177.585 ;
        RECT -228.225 -177.755 -228.055 -177.585 ;
        RECT -222.365 -177.755 -222.195 -177.585 ;
        RECT -218.305 -177.755 -218.135 -177.585 ;
        RECT -212.445 -177.755 -212.275 -177.585 ;
        RECT -208.385 -177.755 -208.215 -177.585 ;
        RECT -202.525 -177.755 -202.355 -177.585 ;
        RECT -198.465 -177.755 -198.295 -177.585 ;
        RECT -192.605 -177.755 -192.435 -177.585 ;
        RECT -188.545 -177.755 -188.375 -177.585 ;
        RECT -182.685 -177.755 -182.515 -177.585 ;
        RECT -178.625 -177.755 -178.455 -177.585 ;
        RECT -172.765 -177.755 -172.595 -177.585 ;
        RECT -168.705 -177.755 -168.535 -177.585 ;
        RECT -162.845 -177.755 -162.675 -177.585 ;
        RECT -158.785 -177.755 -158.615 -177.585 ;
        RECT -152.925 -177.755 -152.755 -177.585 ;
        RECT -148.865 -177.755 -148.695 -177.585 ;
        RECT -143.005 -177.755 -142.835 -177.585 ;
        RECT -138.945 -177.755 -138.775 -177.585 ;
        RECT -133.085 -177.755 -132.915 -177.585 ;
        RECT -129.025 -177.755 -128.855 -177.585 ;
        RECT -123.165 -177.755 -122.995 -177.585 ;
        RECT -119.105 -177.755 -118.935 -177.585 ;
        RECT -113.245 -177.755 -113.075 -177.585 ;
        RECT -109.185 -177.755 -109.015 -177.585 ;
        RECT -103.325 -177.755 -103.155 -177.585 ;
        RECT -99.265 -177.755 -99.095 -177.585 ;
        RECT -93.405 -177.755 -93.235 -177.585 ;
        RECT -89.345 -177.755 -89.175 -177.585 ;
        RECT -83.485 -177.755 -83.315 -177.585 ;
        RECT -79.425 -177.755 -79.255 -177.585 ;
        RECT -73.565 -177.755 -73.395 -177.585 ;
        RECT -69.505 -177.755 -69.335 -177.585 ;
        RECT -63.645 -177.755 -63.475 -177.585 ;
        RECT -59.585 -177.755 -59.415 -177.585 ;
        RECT -53.725 -177.755 -53.555 -177.585 ;
        RECT -49.665 -177.755 -49.495 -177.585 ;
        RECT -43.805 -177.755 -43.635 -177.585 ;
        RECT -39.745 -177.755 -39.575 -177.585 ;
        RECT -33.885 -177.755 -33.715 -177.585 ;
        RECT -29.825 -177.755 -29.655 -177.585 ;
        RECT -23.965 -177.755 -23.795 -177.585 ;
        RECT -19.905 -177.755 -19.735 -177.585 ;
        RECT -14.045 -177.755 -13.875 -177.585 ;
        RECT -9.985 -177.755 -9.815 -177.585 ;
        RECT -4.125 -177.755 -3.955 -177.585 ;
        RECT -0.065 -177.755 0.105 -177.585 ;
        RECT 5.795 -177.755 5.965 -177.585 ;
        RECT 9.855 -177.755 10.025 -177.585 ;
        RECT 15.715 -177.755 15.885 -177.585 ;
        RECT 19.775 -177.755 19.945 -177.585 ;
        RECT 20.935 -177.715 21.105 -177.545 ;
        RECT 20.935 -178.175 21.105 -178.005 ;
        RECT -293.435 -178.625 -293.265 -178.455 ;
        RECT -292.965 -178.635 -292.795 -178.465 ;
        RECT -288.480 -178.605 -288.310 -178.435 ;
        RECT -287.115 -178.605 -286.945 -178.435 ;
        RECT -278.560 -178.605 -278.390 -178.435 ;
        RECT -277.195 -178.605 -277.025 -178.435 ;
        RECT -268.640 -178.605 -268.470 -178.435 ;
        RECT -267.275 -178.605 -267.105 -178.435 ;
        RECT -258.720 -178.605 -258.550 -178.435 ;
        RECT -257.355 -178.605 -257.185 -178.435 ;
        RECT -248.800 -178.605 -248.630 -178.435 ;
        RECT -247.435 -178.605 -247.265 -178.435 ;
        RECT -238.880 -178.605 -238.710 -178.435 ;
        RECT -237.515 -178.605 -237.345 -178.435 ;
        RECT -228.960 -178.605 -228.790 -178.435 ;
        RECT -227.595 -178.605 -227.425 -178.435 ;
        RECT -219.040 -178.605 -218.870 -178.435 ;
        RECT -217.675 -178.605 -217.505 -178.435 ;
        RECT -209.120 -178.605 -208.950 -178.435 ;
        RECT -207.755 -178.605 -207.585 -178.435 ;
        RECT -199.200 -178.605 -199.030 -178.435 ;
        RECT -197.835 -178.605 -197.665 -178.435 ;
        RECT -189.280 -178.605 -189.110 -178.435 ;
        RECT -187.915 -178.605 -187.745 -178.435 ;
        RECT -179.360 -178.605 -179.190 -178.435 ;
        RECT -177.995 -178.605 -177.825 -178.435 ;
        RECT -169.440 -178.605 -169.270 -178.435 ;
        RECT -168.075 -178.605 -167.905 -178.435 ;
        RECT -159.520 -178.605 -159.350 -178.435 ;
        RECT -158.155 -178.605 -157.985 -178.435 ;
        RECT -149.600 -178.605 -149.430 -178.435 ;
        RECT -148.235 -178.605 -148.065 -178.435 ;
        RECT -139.680 -178.605 -139.510 -178.435 ;
        RECT -138.315 -178.605 -138.145 -178.435 ;
        RECT -129.760 -178.605 -129.590 -178.435 ;
        RECT -128.395 -178.605 -128.225 -178.435 ;
        RECT -119.840 -178.605 -119.670 -178.435 ;
        RECT -118.475 -178.605 -118.305 -178.435 ;
        RECT -109.920 -178.605 -109.750 -178.435 ;
        RECT -108.555 -178.605 -108.385 -178.435 ;
        RECT -100.000 -178.605 -99.830 -178.435 ;
        RECT -98.635 -178.605 -98.465 -178.435 ;
        RECT -90.080 -178.605 -89.910 -178.435 ;
        RECT -88.715 -178.605 -88.545 -178.435 ;
        RECT -80.160 -178.605 -79.990 -178.435 ;
        RECT -78.795 -178.605 -78.625 -178.435 ;
        RECT -70.240 -178.605 -70.070 -178.435 ;
        RECT -68.875 -178.605 -68.705 -178.435 ;
        RECT -60.320 -178.605 -60.150 -178.435 ;
        RECT -58.955 -178.605 -58.785 -178.435 ;
        RECT -50.400 -178.605 -50.230 -178.435 ;
        RECT -49.035 -178.605 -48.865 -178.435 ;
        RECT -40.480 -178.605 -40.310 -178.435 ;
        RECT -39.115 -178.605 -38.945 -178.435 ;
        RECT -30.560 -178.605 -30.390 -178.435 ;
        RECT -29.195 -178.605 -29.025 -178.435 ;
        RECT -20.640 -178.605 -20.470 -178.435 ;
        RECT -19.275 -178.605 -19.105 -178.435 ;
        RECT -10.720 -178.605 -10.550 -178.435 ;
        RECT -9.355 -178.605 -9.185 -178.435 ;
        RECT -0.800 -178.605 -0.630 -178.435 ;
        RECT 0.565 -178.605 0.735 -178.435 ;
        RECT 9.120 -178.605 9.290 -178.435 ;
        RECT 10.485 -178.605 10.655 -178.435 ;
        RECT 19.040 -178.605 19.210 -178.435 ;
        RECT 20.405 -178.605 20.575 -178.435 ;
        RECT 20.935 -178.635 21.105 -178.465 ;
        RECT 21.405 -178.625 21.575 -178.455 ;
      LAYER met1 ;
        RECT -291.460 95.140 -291.000 95.145 ;
        RECT -291.460 94.665 -290.520 95.140 ;
        RECT -289.600 95.060 -288.600 95.760 ;
        RECT -279.680 95.060 -278.680 95.760 ;
        RECT -269.760 95.060 -268.760 95.760 ;
        RECT -259.840 95.060 -258.840 95.760 ;
        RECT -249.920 95.060 -248.920 95.760 ;
        RECT -240.000 95.060 -239.000 95.760 ;
        RECT -230.080 95.060 -229.080 95.760 ;
        RECT -220.160 95.060 -219.160 95.760 ;
        RECT -210.240 95.060 -209.240 95.760 ;
        RECT -200.320 95.060 -199.320 95.760 ;
        RECT -190.400 95.060 -189.400 95.760 ;
        RECT -180.480 95.060 -179.480 95.760 ;
        RECT -170.560 95.060 -169.560 95.760 ;
        RECT -160.640 95.060 -159.640 95.760 ;
        RECT -150.720 95.060 -149.720 95.760 ;
        RECT -140.800 95.060 -139.800 95.760 ;
        RECT -130.880 95.060 -129.880 95.760 ;
        RECT -120.960 95.060 -119.960 95.760 ;
        RECT -111.040 95.060 -110.040 95.760 ;
        RECT -101.120 95.060 -100.120 95.760 ;
        RECT -91.200 95.060 -90.200 95.760 ;
        RECT -81.280 95.060 -80.280 95.760 ;
        RECT -71.360 95.060 -70.360 95.760 ;
        RECT -61.440 95.060 -60.440 95.760 ;
        RECT -51.520 95.060 -50.520 95.760 ;
        RECT -41.600 95.060 -40.600 95.760 ;
        RECT -31.680 95.060 -30.680 95.760 ;
        RECT -21.760 95.060 -20.760 95.760 ;
        RECT -11.840 95.060 -10.840 95.760 ;
        RECT -1.920 95.060 -0.920 95.760 ;
        RECT 8.000 95.060 9.000 95.760 ;
        RECT 17.920 95.060 18.920 95.760 ;
        RECT -290.110 94.760 -288.420 95.060 ;
        RECT -280.190 94.760 -278.500 95.060 ;
        RECT -270.270 94.760 -268.580 95.060 ;
        RECT -260.350 94.760 -258.660 95.060 ;
        RECT -250.430 94.760 -248.740 95.060 ;
        RECT -240.510 94.760 -238.820 95.060 ;
        RECT -230.590 94.760 -228.900 95.060 ;
        RECT -220.670 94.760 -218.980 95.060 ;
        RECT -210.750 94.760 -209.060 95.060 ;
        RECT -200.830 94.760 -199.140 95.060 ;
        RECT -190.910 94.760 -189.220 95.060 ;
        RECT -180.990 94.760 -179.300 95.060 ;
        RECT -171.070 94.760 -169.380 95.060 ;
        RECT -161.150 94.760 -159.460 95.060 ;
        RECT -151.230 94.760 -149.540 95.060 ;
        RECT -141.310 94.760 -139.620 95.060 ;
        RECT -131.390 94.760 -129.700 95.060 ;
        RECT -121.470 94.760 -119.780 95.060 ;
        RECT -111.550 94.760 -109.860 95.060 ;
        RECT -101.630 94.760 -99.940 95.060 ;
        RECT -91.710 94.760 -90.020 95.060 ;
        RECT -81.790 94.760 -80.100 95.060 ;
        RECT -71.870 94.760 -70.180 95.060 ;
        RECT -61.950 94.760 -60.260 95.060 ;
        RECT -52.030 94.760 -50.340 95.060 ;
        RECT -42.110 94.760 -40.420 95.060 ;
        RECT -32.190 94.760 -30.500 95.060 ;
        RECT -22.270 94.760 -20.580 95.060 ;
        RECT -12.350 94.760 -10.660 95.060 ;
        RECT -2.430 94.760 -0.740 95.060 ;
        RECT 7.490 94.760 9.180 95.060 ;
        RECT 17.410 94.760 19.100 95.060 ;
        RECT -291.000 93.760 -290.520 94.665 ;
        RECT -289.370 93.890 -289.050 94.180 ;
        RECT -283.490 93.890 -283.170 94.180 ;
        RECT -279.450 93.890 -279.130 94.180 ;
        RECT -273.570 93.890 -273.250 94.180 ;
        RECT -269.530 93.890 -269.210 94.180 ;
        RECT -263.650 93.890 -263.330 94.180 ;
        RECT -259.610 93.890 -259.290 94.180 ;
        RECT -253.730 93.890 -253.410 94.180 ;
        RECT -249.690 93.890 -249.370 94.180 ;
        RECT -243.810 93.890 -243.490 94.180 ;
        RECT -239.770 93.890 -239.450 94.180 ;
        RECT -233.890 93.890 -233.570 94.180 ;
        RECT -229.850 93.890 -229.530 94.180 ;
        RECT -223.970 93.890 -223.650 94.180 ;
        RECT -219.930 93.890 -219.610 94.180 ;
        RECT -214.050 93.890 -213.730 94.180 ;
        RECT -210.010 93.890 -209.690 94.180 ;
        RECT -204.130 93.890 -203.810 94.180 ;
        RECT -200.090 93.890 -199.770 94.180 ;
        RECT -194.210 93.890 -193.890 94.180 ;
        RECT -190.170 93.890 -189.850 94.180 ;
        RECT -184.290 93.890 -183.970 94.180 ;
        RECT -180.250 93.890 -179.930 94.180 ;
        RECT -174.370 93.890 -174.050 94.180 ;
        RECT -170.330 93.890 -170.010 94.180 ;
        RECT -164.450 93.890 -164.130 94.180 ;
        RECT -160.410 93.890 -160.090 94.180 ;
        RECT -154.530 93.890 -154.210 94.180 ;
        RECT -150.490 93.890 -150.170 94.180 ;
        RECT -144.610 93.890 -144.290 94.180 ;
        RECT -140.570 93.890 -140.250 94.180 ;
        RECT -134.690 93.890 -134.370 94.180 ;
        RECT -130.650 93.890 -130.330 94.180 ;
        RECT -124.770 93.890 -124.450 94.180 ;
        RECT -120.730 93.890 -120.410 94.180 ;
        RECT -114.850 93.890 -114.530 94.180 ;
        RECT -110.810 93.890 -110.490 94.180 ;
        RECT -104.930 93.890 -104.610 94.180 ;
        RECT -100.890 93.890 -100.570 94.180 ;
        RECT -95.010 93.890 -94.690 94.180 ;
        RECT -90.970 93.890 -90.650 94.180 ;
        RECT -85.090 93.890 -84.770 94.180 ;
        RECT -81.050 93.890 -80.730 94.180 ;
        RECT -75.170 93.890 -74.850 94.180 ;
        RECT -71.130 93.890 -70.810 94.180 ;
        RECT -65.250 93.890 -64.930 94.180 ;
        RECT -61.210 93.890 -60.890 94.180 ;
        RECT -55.330 93.890 -55.010 94.180 ;
        RECT -51.290 93.890 -50.970 94.180 ;
        RECT -45.410 93.890 -45.090 94.180 ;
        RECT -41.370 93.890 -41.050 94.180 ;
        RECT -35.490 93.890 -35.170 94.180 ;
        RECT -31.450 93.890 -31.130 94.180 ;
        RECT -25.570 93.890 -25.250 94.180 ;
        RECT -21.530 93.890 -21.210 94.180 ;
        RECT -15.650 93.890 -15.330 94.180 ;
        RECT -11.610 93.890 -11.290 94.180 ;
        RECT -5.730 93.890 -5.410 94.180 ;
        RECT -1.690 93.890 -1.370 94.180 ;
        RECT 4.190 93.890 4.510 94.180 ;
        RECT 8.230 93.890 8.550 94.180 ;
        RECT 14.110 93.890 14.430 94.180 ;
        RECT 18.150 93.890 18.470 94.180 ;
        RECT 24.030 93.890 24.350 94.180 ;
        RECT -291.460 93.090 -289.620 93.570 ;
        RECT -289.290 92.760 -289.100 93.890 ;
        RECT -283.440 92.760 -283.250 93.890 ;
        RECT -279.370 92.760 -279.180 93.890 ;
        RECT -273.520 92.760 -273.330 93.890 ;
        RECT -269.450 92.760 -269.260 93.890 ;
        RECT -263.600 92.760 -263.410 93.890 ;
        RECT -259.530 92.760 -259.340 93.890 ;
        RECT -253.680 92.760 -253.490 93.890 ;
        RECT -249.610 92.760 -249.420 93.890 ;
        RECT -243.760 92.760 -243.570 93.890 ;
        RECT -239.690 92.760 -239.500 93.890 ;
        RECT -233.840 92.760 -233.650 93.890 ;
        RECT -229.770 92.760 -229.580 93.890 ;
        RECT -223.920 92.760 -223.730 93.890 ;
        RECT -219.850 92.760 -219.660 93.890 ;
        RECT -214.000 92.760 -213.810 93.890 ;
        RECT -209.930 92.760 -209.740 93.890 ;
        RECT -204.080 92.760 -203.890 93.890 ;
        RECT -200.010 92.760 -199.820 93.890 ;
        RECT -194.160 92.760 -193.970 93.890 ;
        RECT -190.090 92.760 -189.900 93.890 ;
        RECT -184.240 92.760 -184.050 93.890 ;
        RECT -180.170 92.760 -179.980 93.890 ;
        RECT -174.320 92.760 -174.130 93.890 ;
        RECT -170.250 92.760 -170.060 93.890 ;
        RECT -164.400 92.760 -164.210 93.890 ;
        RECT -160.330 92.760 -160.140 93.890 ;
        RECT -154.480 92.760 -154.290 93.890 ;
        RECT -150.410 92.760 -150.220 93.890 ;
        RECT -144.560 92.760 -144.370 93.890 ;
        RECT -140.490 92.760 -140.300 93.890 ;
        RECT -134.640 92.760 -134.450 93.890 ;
        RECT -130.570 92.760 -130.380 93.890 ;
        RECT -124.720 92.760 -124.530 93.890 ;
        RECT -120.650 92.760 -120.460 93.890 ;
        RECT -114.800 92.760 -114.610 93.890 ;
        RECT -110.730 92.760 -110.540 93.890 ;
        RECT -104.880 92.760 -104.690 93.890 ;
        RECT -100.810 92.760 -100.620 93.890 ;
        RECT -94.960 92.760 -94.770 93.890 ;
        RECT -90.890 92.760 -90.700 93.890 ;
        RECT -85.040 92.760 -84.850 93.890 ;
        RECT -80.970 92.760 -80.780 93.890 ;
        RECT -75.120 92.760 -74.930 93.890 ;
        RECT -71.050 92.760 -70.860 93.890 ;
        RECT -65.200 92.760 -65.010 93.890 ;
        RECT -61.130 92.760 -60.940 93.890 ;
        RECT -55.280 92.760 -55.090 93.890 ;
        RECT -51.210 92.760 -51.020 93.890 ;
        RECT -45.360 92.760 -45.170 93.890 ;
        RECT -41.290 92.760 -41.100 93.890 ;
        RECT -35.440 92.760 -35.250 93.890 ;
        RECT -31.370 92.760 -31.180 93.890 ;
        RECT -25.520 92.760 -25.330 93.890 ;
        RECT -21.450 92.760 -21.260 93.890 ;
        RECT -15.600 92.760 -15.410 93.890 ;
        RECT -11.530 92.760 -11.340 93.890 ;
        RECT -5.680 92.760 -5.490 93.890 ;
        RECT -1.610 92.760 -1.420 93.890 ;
        RECT 4.240 92.760 4.430 93.890 ;
        RECT 8.310 92.760 8.500 93.890 ;
        RECT 14.160 92.760 14.350 93.890 ;
        RECT 18.230 92.760 18.420 93.890 ;
        RECT 24.080 92.760 24.270 93.890 ;
        RECT 24.600 93.090 26.440 93.570 ;
        RECT -290.050 92.610 -288.110 92.760 ;
        RECT -290.050 92.460 -289.710 92.610 ;
        RECT -290.050 92.260 -289.730 92.290 ;
        RECT -290.050 92.120 -289.230 92.260 ;
        RECT -290.050 92.010 -289.730 92.120 ;
        RECT -289.390 91.330 -289.230 92.120 ;
        RECT -288.270 91.820 -288.110 92.610 ;
        RECT -284.430 92.610 -282.490 92.760 ;
        RECT -287.770 91.820 -287.450 91.930 ;
        RECT -288.270 91.680 -287.450 91.820 ;
        RECT -287.770 91.650 -287.450 91.680 ;
        RECT -285.090 91.820 -284.770 91.930 ;
        RECT -284.430 91.820 -284.270 92.610 ;
        RECT -282.830 92.460 -282.490 92.610 ;
        RECT -280.130 92.610 -278.190 92.760 ;
        RECT -280.130 92.460 -279.790 92.610 ;
        RECT -282.810 92.260 -282.490 92.290 ;
        RECT -285.090 91.680 -284.270 91.820 ;
        RECT -283.310 92.120 -282.490 92.260 ;
        RECT -285.090 91.650 -284.770 91.680 ;
        RECT -287.790 91.330 -287.450 91.480 ;
        RECT -289.390 91.180 -287.450 91.330 ;
        RECT -285.090 91.330 -284.750 91.480 ;
        RECT -283.310 91.330 -283.150 92.120 ;
        RECT -282.810 92.010 -282.490 92.120 ;
        RECT -280.130 92.260 -279.810 92.290 ;
        RECT -280.130 92.120 -279.310 92.260 ;
        RECT -280.130 92.010 -279.810 92.120 ;
        RECT -285.090 91.180 -283.150 91.330 ;
        RECT -279.470 91.330 -279.310 92.120 ;
        RECT -278.350 91.820 -278.190 92.610 ;
        RECT -274.510 92.610 -272.570 92.760 ;
        RECT -277.850 91.820 -277.530 91.930 ;
        RECT -278.350 91.680 -277.530 91.820 ;
        RECT -277.850 91.650 -277.530 91.680 ;
        RECT -275.170 91.820 -274.850 91.930 ;
        RECT -274.510 91.820 -274.350 92.610 ;
        RECT -272.910 92.460 -272.570 92.610 ;
        RECT -270.210 92.610 -268.270 92.760 ;
        RECT -270.210 92.460 -269.870 92.610 ;
        RECT -272.890 92.260 -272.570 92.290 ;
        RECT -275.170 91.680 -274.350 91.820 ;
        RECT -273.390 92.120 -272.570 92.260 ;
        RECT -275.170 91.650 -274.850 91.680 ;
        RECT -277.870 91.330 -277.530 91.480 ;
        RECT -279.470 91.180 -277.530 91.330 ;
        RECT -275.170 91.330 -274.830 91.480 ;
        RECT -273.390 91.330 -273.230 92.120 ;
        RECT -272.890 92.010 -272.570 92.120 ;
        RECT -270.210 92.260 -269.890 92.290 ;
        RECT -270.210 92.120 -269.390 92.260 ;
        RECT -270.210 92.010 -269.890 92.120 ;
        RECT -275.170 91.180 -273.230 91.330 ;
        RECT -269.550 91.330 -269.390 92.120 ;
        RECT -268.430 91.820 -268.270 92.610 ;
        RECT -264.590 92.610 -262.650 92.760 ;
        RECT -267.930 91.820 -267.610 91.930 ;
        RECT -268.430 91.680 -267.610 91.820 ;
        RECT -267.930 91.650 -267.610 91.680 ;
        RECT -265.250 91.820 -264.930 91.930 ;
        RECT -264.590 91.820 -264.430 92.610 ;
        RECT -262.990 92.460 -262.650 92.610 ;
        RECT -260.290 92.610 -258.350 92.760 ;
        RECT -260.290 92.460 -259.950 92.610 ;
        RECT -262.970 92.260 -262.650 92.290 ;
        RECT -265.250 91.680 -264.430 91.820 ;
        RECT -263.470 92.120 -262.650 92.260 ;
        RECT -265.250 91.650 -264.930 91.680 ;
        RECT -267.950 91.330 -267.610 91.480 ;
        RECT -269.550 91.180 -267.610 91.330 ;
        RECT -265.250 91.330 -264.910 91.480 ;
        RECT -263.470 91.330 -263.310 92.120 ;
        RECT -262.970 92.010 -262.650 92.120 ;
        RECT -260.290 92.260 -259.970 92.290 ;
        RECT -260.290 92.120 -259.470 92.260 ;
        RECT -260.290 92.010 -259.970 92.120 ;
        RECT -265.250 91.180 -263.310 91.330 ;
        RECT -259.630 91.330 -259.470 92.120 ;
        RECT -258.510 91.820 -258.350 92.610 ;
        RECT -254.670 92.610 -252.730 92.760 ;
        RECT -258.010 91.820 -257.690 91.930 ;
        RECT -258.510 91.680 -257.690 91.820 ;
        RECT -258.010 91.650 -257.690 91.680 ;
        RECT -255.330 91.820 -255.010 91.930 ;
        RECT -254.670 91.820 -254.510 92.610 ;
        RECT -253.070 92.460 -252.730 92.610 ;
        RECT -250.370 92.610 -248.430 92.760 ;
        RECT -250.370 92.460 -250.030 92.610 ;
        RECT -253.050 92.260 -252.730 92.290 ;
        RECT -255.330 91.680 -254.510 91.820 ;
        RECT -253.550 92.120 -252.730 92.260 ;
        RECT -255.330 91.650 -255.010 91.680 ;
        RECT -258.030 91.330 -257.690 91.480 ;
        RECT -259.630 91.180 -257.690 91.330 ;
        RECT -255.330 91.330 -254.990 91.480 ;
        RECT -253.550 91.330 -253.390 92.120 ;
        RECT -253.050 92.010 -252.730 92.120 ;
        RECT -250.370 92.260 -250.050 92.290 ;
        RECT -250.370 92.120 -249.550 92.260 ;
        RECT -250.370 92.010 -250.050 92.120 ;
        RECT -255.330 91.180 -253.390 91.330 ;
        RECT -249.710 91.330 -249.550 92.120 ;
        RECT -248.590 91.820 -248.430 92.610 ;
        RECT -244.750 92.610 -242.810 92.760 ;
        RECT -248.090 91.820 -247.770 91.930 ;
        RECT -248.590 91.680 -247.770 91.820 ;
        RECT -248.090 91.650 -247.770 91.680 ;
        RECT -245.410 91.820 -245.090 91.930 ;
        RECT -244.750 91.820 -244.590 92.610 ;
        RECT -243.150 92.460 -242.810 92.610 ;
        RECT -240.450 92.610 -238.510 92.760 ;
        RECT -240.450 92.460 -240.110 92.610 ;
        RECT -243.130 92.260 -242.810 92.290 ;
        RECT -245.410 91.680 -244.590 91.820 ;
        RECT -243.630 92.120 -242.810 92.260 ;
        RECT -245.410 91.650 -245.090 91.680 ;
        RECT -248.110 91.330 -247.770 91.480 ;
        RECT -249.710 91.180 -247.770 91.330 ;
        RECT -245.410 91.330 -245.070 91.480 ;
        RECT -243.630 91.330 -243.470 92.120 ;
        RECT -243.130 92.010 -242.810 92.120 ;
        RECT -240.450 92.260 -240.130 92.290 ;
        RECT -240.450 92.120 -239.630 92.260 ;
        RECT -240.450 92.010 -240.130 92.120 ;
        RECT -245.410 91.180 -243.470 91.330 ;
        RECT -239.790 91.330 -239.630 92.120 ;
        RECT -238.670 91.820 -238.510 92.610 ;
        RECT -234.830 92.610 -232.890 92.760 ;
        RECT -238.170 91.820 -237.850 91.930 ;
        RECT -238.670 91.680 -237.850 91.820 ;
        RECT -238.170 91.650 -237.850 91.680 ;
        RECT -235.490 91.820 -235.170 91.930 ;
        RECT -234.830 91.820 -234.670 92.610 ;
        RECT -233.230 92.460 -232.890 92.610 ;
        RECT -230.530 92.610 -228.590 92.760 ;
        RECT -230.530 92.460 -230.190 92.610 ;
        RECT -233.210 92.260 -232.890 92.290 ;
        RECT -235.490 91.680 -234.670 91.820 ;
        RECT -233.710 92.120 -232.890 92.260 ;
        RECT -235.490 91.650 -235.170 91.680 ;
        RECT -238.190 91.330 -237.850 91.480 ;
        RECT -239.790 91.180 -237.850 91.330 ;
        RECT -235.490 91.330 -235.150 91.480 ;
        RECT -233.710 91.330 -233.550 92.120 ;
        RECT -233.210 92.010 -232.890 92.120 ;
        RECT -230.530 92.260 -230.210 92.290 ;
        RECT -230.530 92.120 -229.710 92.260 ;
        RECT -230.530 92.010 -230.210 92.120 ;
        RECT -235.490 91.180 -233.550 91.330 ;
        RECT -229.870 91.330 -229.710 92.120 ;
        RECT -228.750 91.820 -228.590 92.610 ;
        RECT -224.910 92.610 -222.970 92.760 ;
        RECT -228.250 91.820 -227.930 91.930 ;
        RECT -228.750 91.680 -227.930 91.820 ;
        RECT -228.250 91.650 -227.930 91.680 ;
        RECT -225.570 91.820 -225.250 91.930 ;
        RECT -224.910 91.820 -224.750 92.610 ;
        RECT -223.310 92.460 -222.970 92.610 ;
        RECT -220.610 92.610 -218.670 92.760 ;
        RECT -220.610 92.460 -220.270 92.610 ;
        RECT -223.290 92.260 -222.970 92.290 ;
        RECT -225.570 91.680 -224.750 91.820 ;
        RECT -223.790 92.120 -222.970 92.260 ;
        RECT -225.570 91.650 -225.250 91.680 ;
        RECT -228.270 91.330 -227.930 91.480 ;
        RECT -229.870 91.180 -227.930 91.330 ;
        RECT -225.570 91.330 -225.230 91.480 ;
        RECT -223.790 91.330 -223.630 92.120 ;
        RECT -223.290 92.010 -222.970 92.120 ;
        RECT -220.610 92.260 -220.290 92.290 ;
        RECT -220.610 92.120 -219.790 92.260 ;
        RECT -220.610 92.010 -220.290 92.120 ;
        RECT -225.570 91.180 -223.630 91.330 ;
        RECT -219.950 91.330 -219.790 92.120 ;
        RECT -218.830 91.820 -218.670 92.610 ;
        RECT -214.990 92.610 -213.050 92.760 ;
        RECT -218.330 91.820 -218.010 91.930 ;
        RECT -218.830 91.680 -218.010 91.820 ;
        RECT -218.330 91.650 -218.010 91.680 ;
        RECT -215.650 91.820 -215.330 91.930 ;
        RECT -214.990 91.820 -214.830 92.610 ;
        RECT -213.390 92.460 -213.050 92.610 ;
        RECT -210.690 92.610 -208.750 92.760 ;
        RECT -210.690 92.460 -210.350 92.610 ;
        RECT -213.370 92.260 -213.050 92.290 ;
        RECT -215.650 91.680 -214.830 91.820 ;
        RECT -213.870 92.120 -213.050 92.260 ;
        RECT -215.650 91.650 -215.330 91.680 ;
        RECT -218.350 91.330 -218.010 91.480 ;
        RECT -219.950 91.180 -218.010 91.330 ;
        RECT -215.650 91.330 -215.310 91.480 ;
        RECT -213.870 91.330 -213.710 92.120 ;
        RECT -213.370 92.010 -213.050 92.120 ;
        RECT -210.690 92.260 -210.370 92.290 ;
        RECT -210.690 92.120 -209.870 92.260 ;
        RECT -210.690 92.010 -210.370 92.120 ;
        RECT -215.650 91.180 -213.710 91.330 ;
        RECT -210.030 91.330 -209.870 92.120 ;
        RECT -208.910 91.820 -208.750 92.610 ;
        RECT -205.070 92.610 -203.130 92.760 ;
        RECT -208.410 91.820 -208.090 91.930 ;
        RECT -208.910 91.680 -208.090 91.820 ;
        RECT -208.410 91.650 -208.090 91.680 ;
        RECT -205.730 91.820 -205.410 91.930 ;
        RECT -205.070 91.820 -204.910 92.610 ;
        RECT -203.470 92.460 -203.130 92.610 ;
        RECT -200.770 92.610 -198.830 92.760 ;
        RECT -200.770 92.460 -200.430 92.610 ;
        RECT -203.450 92.260 -203.130 92.290 ;
        RECT -205.730 91.680 -204.910 91.820 ;
        RECT -203.950 92.120 -203.130 92.260 ;
        RECT -205.730 91.650 -205.410 91.680 ;
        RECT -208.430 91.330 -208.090 91.480 ;
        RECT -210.030 91.180 -208.090 91.330 ;
        RECT -205.730 91.330 -205.390 91.480 ;
        RECT -203.950 91.330 -203.790 92.120 ;
        RECT -203.450 92.010 -203.130 92.120 ;
        RECT -200.770 92.260 -200.450 92.290 ;
        RECT -200.770 92.120 -199.950 92.260 ;
        RECT -200.770 92.010 -200.450 92.120 ;
        RECT -205.730 91.180 -203.790 91.330 ;
        RECT -200.110 91.330 -199.950 92.120 ;
        RECT -198.990 91.820 -198.830 92.610 ;
        RECT -195.150 92.610 -193.210 92.760 ;
        RECT -198.490 91.820 -198.170 91.930 ;
        RECT -198.990 91.680 -198.170 91.820 ;
        RECT -198.490 91.650 -198.170 91.680 ;
        RECT -195.810 91.820 -195.490 91.930 ;
        RECT -195.150 91.820 -194.990 92.610 ;
        RECT -193.550 92.460 -193.210 92.610 ;
        RECT -190.850 92.610 -188.910 92.760 ;
        RECT -190.850 92.460 -190.510 92.610 ;
        RECT -193.530 92.260 -193.210 92.290 ;
        RECT -195.810 91.680 -194.990 91.820 ;
        RECT -194.030 92.120 -193.210 92.260 ;
        RECT -195.810 91.650 -195.490 91.680 ;
        RECT -198.510 91.330 -198.170 91.480 ;
        RECT -200.110 91.180 -198.170 91.330 ;
        RECT -195.810 91.330 -195.470 91.480 ;
        RECT -194.030 91.330 -193.870 92.120 ;
        RECT -193.530 92.010 -193.210 92.120 ;
        RECT -190.850 92.260 -190.530 92.290 ;
        RECT -190.850 92.120 -190.030 92.260 ;
        RECT -190.850 92.010 -190.530 92.120 ;
        RECT -195.810 91.180 -193.870 91.330 ;
        RECT -190.190 91.330 -190.030 92.120 ;
        RECT -189.070 91.820 -188.910 92.610 ;
        RECT -185.230 92.610 -183.290 92.760 ;
        RECT -188.570 91.820 -188.250 91.930 ;
        RECT -189.070 91.680 -188.250 91.820 ;
        RECT -188.570 91.650 -188.250 91.680 ;
        RECT -185.890 91.820 -185.570 91.930 ;
        RECT -185.230 91.820 -185.070 92.610 ;
        RECT -183.630 92.460 -183.290 92.610 ;
        RECT -180.930 92.610 -178.990 92.760 ;
        RECT -180.930 92.460 -180.590 92.610 ;
        RECT -183.610 92.260 -183.290 92.290 ;
        RECT -185.890 91.680 -185.070 91.820 ;
        RECT -184.110 92.120 -183.290 92.260 ;
        RECT -185.890 91.650 -185.570 91.680 ;
        RECT -188.590 91.330 -188.250 91.480 ;
        RECT -190.190 91.180 -188.250 91.330 ;
        RECT -185.890 91.330 -185.550 91.480 ;
        RECT -184.110 91.330 -183.950 92.120 ;
        RECT -183.610 92.010 -183.290 92.120 ;
        RECT -180.930 92.260 -180.610 92.290 ;
        RECT -180.930 92.120 -180.110 92.260 ;
        RECT -180.930 92.010 -180.610 92.120 ;
        RECT -185.890 91.180 -183.950 91.330 ;
        RECT -180.270 91.330 -180.110 92.120 ;
        RECT -179.150 91.820 -178.990 92.610 ;
        RECT -175.310 92.610 -173.370 92.760 ;
        RECT -178.650 91.820 -178.330 91.930 ;
        RECT -179.150 91.680 -178.330 91.820 ;
        RECT -178.650 91.650 -178.330 91.680 ;
        RECT -175.970 91.820 -175.650 91.930 ;
        RECT -175.310 91.820 -175.150 92.610 ;
        RECT -173.710 92.460 -173.370 92.610 ;
        RECT -171.010 92.610 -169.070 92.760 ;
        RECT -171.010 92.460 -170.670 92.610 ;
        RECT -173.690 92.260 -173.370 92.290 ;
        RECT -175.970 91.680 -175.150 91.820 ;
        RECT -174.190 92.120 -173.370 92.260 ;
        RECT -175.970 91.650 -175.650 91.680 ;
        RECT -178.670 91.330 -178.330 91.480 ;
        RECT -180.270 91.180 -178.330 91.330 ;
        RECT -175.970 91.330 -175.630 91.480 ;
        RECT -174.190 91.330 -174.030 92.120 ;
        RECT -173.690 92.010 -173.370 92.120 ;
        RECT -171.010 92.260 -170.690 92.290 ;
        RECT -171.010 92.120 -170.190 92.260 ;
        RECT -171.010 92.010 -170.690 92.120 ;
        RECT -175.970 91.180 -174.030 91.330 ;
        RECT -170.350 91.330 -170.190 92.120 ;
        RECT -169.230 91.820 -169.070 92.610 ;
        RECT -165.390 92.610 -163.450 92.760 ;
        RECT -168.730 91.820 -168.410 91.930 ;
        RECT -169.230 91.680 -168.410 91.820 ;
        RECT -168.730 91.650 -168.410 91.680 ;
        RECT -166.050 91.820 -165.730 91.930 ;
        RECT -165.390 91.820 -165.230 92.610 ;
        RECT -163.790 92.460 -163.450 92.610 ;
        RECT -161.090 92.610 -159.150 92.760 ;
        RECT -161.090 92.460 -160.750 92.610 ;
        RECT -163.770 92.260 -163.450 92.290 ;
        RECT -166.050 91.680 -165.230 91.820 ;
        RECT -164.270 92.120 -163.450 92.260 ;
        RECT -166.050 91.650 -165.730 91.680 ;
        RECT -168.750 91.330 -168.410 91.480 ;
        RECT -170.350 91.180 -168.410 91.330 ;
        RECT -166.050 91.330 -165.710 91.480 ;
        RECT -164.270 91.330 -164.110 92.120 ;
        RECT -163.770 92.010 -163.450 92.120 ;
        RECT -161.090 92.260 -160.770 92.290 ;
        RECT -161.090 92.120 -160.270 92.260 ;
        RECT -161.090 92.010 -160.770 92.120 ;
        RECT -166.050 91.180 -164.110 91.330 ;
        RECT -160.430 91.330 -160.270 92.120 ;
        RECT -159.310 91.820 -159.150 92.610 ;
        RECT -155.470 92.610 -153.530 92.760 ;
        RECT -158.810 91.820 -158.490 91.930 ;
        RECT -159.310 91.680 -158.490 91.820 ;
        RECT -158.810 91.650 -158.490 91.680 ;
        RECT -156.130 91.820 -155.810 91.930 ;
        RECT -155.470 91.820 -155.310 92.610 ;
        RECT -153.870 92.460 -153.530 92.610 ;
        RECT -151.170 92.610 -149.230 92.760 ;
        RECT -151.170 92.460 -150.830 92.610 ;
        RECT -153.850 92.260 -153.530 92.290 ;
        RECT -156.130 91.680 -155.310 91.820 ;
        RECT -154.350 92.120 -153.530 92.260 ;
        RECT -156.130 91.650 -155.810 91.680 ;
        RECT -158.830 91.330 -158.490 91.480 ;
        RECT -160.430 91.180 -158.490 91.330 ;
        RECT -156.130 91.330 -155.790 91.480 ;
        RECT -154.350 91.330 -154.190 92.120 ;
        RECT -153.850 92.010 -153.530 92.120 ;
        RECT -151.170 92.260 -150.850 92.290 ;
        RECT -151.170 92.120 -150.350 92.260 ;
        RECT -151.170 92.010 -150.850 92.120 ;
        RECT -156.130 91.180 -154.190 91.330 ;
        RECT -150.510 91.330 -150.350 92.120 ;
        RECT -149.390 91.820 -149.230 92.610 ;
        RECT -145.550 92.610 -143.610 92.760 ;
        RECT -148.890 91.820 -148.570 91.930 ;
        RECT -149.390 91.680 -148.570 91.820 ;
        RECT -148.890 91.650 -148.570 91.680 ;
        RECT -146.210 91.820 -145.890 91.930 ;
        RECT -145.550 91.820 -145.390 92.610 ;
        RECT -143.950 92.460 -143.610 92.610 ;
        RECT -141.250 92.610 -139.310 92.760 ;
        RECT -141.250 92.460 -140.910 92.610 ;
        RECT -143.930 92.260 -143.610 92.290 ;
        RECT -146.210 91.680 -145.390 91.820 ;
        RECT -144.430 92.120 -143.610 92.260 ;
        RECT -146.210 91.650 -145.890 91.680 ;
        RECT -148.910 91.330 -148.570 91.480 ;
        RECT -150.510 91.180 -148.570 91.330 ;
        RECT -146.210 91.330 -145.870 91.480 ;
        RECT -144.430 91.330 -144.270 92.120 ;
        RECT -143.930 92.010 -143.610 92.120 ;
        RECT -141.250 92.260 -140.930 92.290 ;
        RECT -141.250 92.120 -140.430 92.260 ;
        RECT -141.250 92.010 -140.930 92.120 ;
        RECT -146.210 91.180 -144.270 91.330 ;
        RECT -140.590 91.330 -140.430 92.120 ;
        RECT -139.470 91.820 -139.310 92.610 ;
        RECT -135.630 92.610 -133.690 92.760 ;
        RECT -138.970 91.820 -138.650 91.930 ;
        RECT -139.470 91.680 -138.650 91.820 ;
        RECT -138.970 91.650 -138.650 91.680 ;
        RECT -136.290 91.820 -135.970 91.930 ;
        RECT -135.630 91.820 -135.470 92.610 ;
        RECT -134.030 92.460 -133.690 92.610 ;
        RECT -131.330 92.610 -129.390 92.760 ;
        RECT -131.330 92.460 -130.990 92.610 ;
        RECT -134.010 92.260 -133.690 92.290 ;
        RECT -136.290 91.680 -135.470 91.820 ;
        RECT -134.510 92.120 -133.690 92.260 ;
        RECT -136.290 91.650 -135.970 91.680 ;
        RECT -138.990 91.330 -138.650 91.480 ;
        RECT -140.590 91.180 -138.650 91.330 ;
        RECT -136.290 91.330 -135.950 91.480 ;
        RECT -134.510 91.330 -134.350 92.120 ;
        RECT -134.010 92.010 -133.690 92.120 ;
        RECT -131.330 92.260 -131.010 92.290 ;
        RECT -131.330 92.120 -130.510 92.260 ;
        RECT -131.330 92.010 -131.010 92.120 ;
        RECT -136.290 91.180 -134.350 91.330 ;
        RECT -130.670 91.330 -130.510 92.120 ;
        RECT -129.550 91.820 -129.390 92.610 ;
        RECT -125.710 92.610 -123.770 92.760 ;
        RECT -129.050 91.820 -128.730 91.930 ;
        RECT -129.550 91.680 -128.730 91.820 ;
        RECT -129.050 91.650 -128.730 91.680 ;
        RECT -126.370 91.820 -126.050 91.930 ;
        RECT -125.710 91.820 -125.550 92.610 ;
        RECT -124.110 92.460 -123.770 92.610 ;
        RECT -121.410 92.610 -119.470 92.760 ;
        RECT -121.410 92.460 -121.070 92.610 ;
        RECT -124.090 92.260 -123.770 92.290 ;
        RECT -126.370 91.680 -125.550 91.820 ;
        RECT -124.590 92.120 -123.770 92.260 ;
        RECT -126.370 91.650 -126.050 91.680 ;
        RECT -129.070 91.330 -128.730 91.480 ;
        RECT -130.670 91.180 -128.730 91.330 ;
        RECT -126.370 91.330 -126.030 91.480 ;
        RECT -124.590 91.330 -124.430 92.120 ;
        RECT -124.090 92.010 -123.770 92.120 ;
        RECT -121.410 92.260 -121.090 92.290 ;
        RECT -121.410 92.120 -120.590 92.260 ;
        RECT -121.410 92.010 -121.090 92.120 ;
        RECT -126.370 91.180 -124.430 91.330 ;
        RECT -120.750 91.330 -120.590 92.120 ;
        RECT -119.630 91.820 -119.470 92.610 ;
        RECT -115.790 92.610 -113.850 92.760 ;
        RECT -119.130 91.820 -118.810 91.930 ;
        RECT -119.630 91.680 -118.810 91.820 ;
        RECT -119.130 91.650 -118.810 91.680 ;
        RECT -116.450 91.820 -116.130 91.930 ;
        RECT -115.790 91.820 -115.630 92.610 ;
        RECT -114.190 92.460 -113.850 92.610 ;
        RECT -111.490 92.610 -109.550 92.760 ;
        RECT -111.490 92.460 -111.150 92.610 ;
        RECT -114.170 92.260 -113.850 92.290 ;
        RECT -116.450 91.680 -115.630 91.820 ;
        RECT -114.670 92.120 -113.850 92.260 ;
        RECT -116.450 91.650 -116.130 91.680 ;
        RECT -119.150 91.330 -118.810 91.480 ;
        RECT -120.750 91.180 -118.810 91.330 ;
        RECT -116.450 91.330 -116.110 91.480 ;
        RECT -114.670 91.330 -114.510 92.120 ;
        RECT -114.170 92.010 -113.850 92.120 ;
        RECT -111.490 92.260 -111.170 92.290 ;
        RECT -111.490 92.120 -110.670 92.260 ;
        RECT -111.490 92.010 -111.170 92.120 ;
        RECT -116.450 91.180 -114.510 91.330 ;
        RECT -110.830 91.330 -110.670 92.120 ;
        RECT -109.710 91.820 -109.550 92.610 ;
        RECT -105.870 92.610 -103.930 92.760 ;
        RECT -109.210 91.820 -108.890 91.930 ;
        RECT -109.710 91.680 -108.890 91.820 ;
        RECT -109.210 91.650 -108.890 91.680 ;
        RECT -106.530 91.820 -106.210 91.930 ;
        RECT -105.870 91.820 -105.710 92.610 ;
        RECT -104.270 92.460 -103.930 92.610 ;
        RECT -101.570 92.610 -99.630 92.760 ;
        RECT -101.570 92.460 -101.230 92.610 ;
        RECT -104.250 92.260 -103.930 92.290 ;
        RECT -106.530 91.680 -105.710 91.820 ;
        RECT -104.750 92.120 -103.930 92.260 ;
        RECT -106.530 91.650 -106.210 91.680 ;
        RECT -109.230 91.330 -108.890 91.480 ;
        RECT -110.830 91.180 -108.890 91.330 ;
        RECT -106.530 91.330 -106.190 91.480 ;
        RECT -104.750 91.330 -104.590 92.120 ;
        RECT -104.250 92.010 -103.930 92.120 ;
        RECT -101.570 92.260 -101.250 92.290 ;
        RECT -101.570 92.120 -100.750 92.260 ;
        RECT -101.570 92.010 -101.250 92.120 ;
        RECT -106.530 91.180 -104.590 91.330 ;
        RECT -100.910 91.330 -100.750 92.120 ;
        RECT -99.790 91.820 -99.630 92.610 ;
        RECT -95.950 92.610 -94.010 92.760 ;
        RECT -99.290 91.820 -98.970 91.930 ;
        RECT -99.790 91.680 -98.970 91.820 ;
        RECT -99.290 91.650 -98.970 91.680 ;
        RECT -96.610 91.820 -96.290 91.930 ;
        RECT -95.950 91.820 -95.790 92.610 ;
        RECT -94.350 92.460 -94.010 92.610 ;
        RECT -91.650 92.610 -89.710 92.760 ;
        RECT -91.650 92.460 -91.310 92.610 ;
        RECT -94.330 92.260 -94.010 92.290 ;
        RECT -96.610 91.680 -95.790 91.820 ;
        RECT -94.830 92.120 -94.010 92.260 ;
        RECT -96.610 91.650 -96.290 91.680 ;
        RECT -99.310 91.330 -98.970 91.480 ;
        RECT -100.910 91.180 -98.970 91.330 ;
        RECT -96.610 91.330 -96.270 91.480 ;
        RECT -94.830 91.330 -94.670 92.120 ;
        RECT -94.330 92.010 -94.010 92.120 ;
        RECT -91.650 92.260 -91.330 92.290 ;
        RECT -91.650 92.120 -90.830 92.260 ;
        RECT -91.650 92.010 -91.330 92.120 ;
        RECT -96.610 91.180 -94.670 91.330 ;
        RECT -90.990 91.330 -90.830 92.120 ;
        RECT -89.870 91.820 -89.710 92.610 ;
        RECT -86.030 92.610 -84.090 92.760 ;
        RECT -89.370 91.820 -89.050 91.930 ;
        RECT -89.870 91.680 -89.050 91.820 ;
        RECT -89.370 91.650 -89.050 91.680 ;
        RECT -86.690 91.820 -86.370 91.930 ;
        RECT -86.030 91.820 -85.870 92.610 ;
        RECT -84.430 92.460 -84.090 92.610 ;
        RECT -81.730 92.610 -79.790 92.760 ;
        RECT -81.730 92.460 -81.390 92.610 ;
        RECT -84.410 92.260 -84.090 92.290 ;
        RECT -86.690 91.680 -85.870 91.820 ;
        RECT -84.910 92.120 -84.090 92.260 ;
        RECT -86.690 91.650 -86.370 91.680 ;
        RECT -89.390 91.330 -89.050 91.480 ;
        RECT -90.990 91.180 -89.050 91.330 ;
        RECT -86.690 91.330 -86.350 91.480 ;
        RECT -84.910 91.330 -84.750 92.120 ;
        RECT -84.410 92.010 -84.090 92.120 ;
        RECT -81.730 92.260 -81.410 92.290 ;
        RECT -81.730 92.120 -80.910 92.260 ;
        RECT -81.730 92.010 -81.410 92.120 ;
        RECT -86.690 91.180 -84.750 91.330 ;
        RECT -81.070 91.330 -80.910 92.120 ;
        RECT -79.950 91.820 -79.790 92.610 ;
        RECT -76.110 92.610 -74.170 92.760 ;
        RECT -79.450 91.820 -79.130 91.930 ;
        RECT -79.950 91.680 -79.130 91.820 ;
        RECT -79.450 91.650 -79.130 91.680 ;
        RECT -76.770 91.820 -76.450 91.930 ;
        RECT -76.110 91.820 -75.950 92.610 ;
        RECT -74.510 92.460 -74.170 92.610 ;
        RECT -71.810 92.610 -69.870 92.760 ;
        RECT -71.810 92.460 -71.470 92.610 ;
        RECT -74.490 92.260 -74.170 92.290 ;
        RECT -76.770 91.680 -75.950 91.820 ;
        RECT -74.990 92.120 -74.170 92.260 ;
        RECT -76.770 91.650 -76.450 91.680 ;
        RECT -79.470 91.330 -79.130 91.480 ;
        RECT -81.070 91.180 -79.130 91.330 ;
        RECT -76.770 91.330 -76.430 91.480 ;
        RECT -74.990 91.330 -74.830 92.120 ;
        RECT -74.490 92.010 -74.170 92.120 ;
        RECT -71.810 92.260 -71.490 92.290 ;
        RECT -71.810 92.120 -70.990 92.260 ;
        RECT -71.810 92.010 -71.490 92.120 ;
        RECT -76.770 91.180 -74.830 91.330 ;
        RECT -71.150 91.330 -70.990 92.120 ;
        RECT -70.030 91.820 -69.870 92.610 ;
        RECT -66.190 92.610 -64.250 92.760 ;
        RECT -69.530 91.820 -69.210 91.930 ;
        RECT -70.030 91.680 -69.210 91.820 ;
        RECT -69.530 91.650 -69.210 91.680 ;
        RECT -66.850 91.820 -66.530 91.930 ;
        RECT -66.190 91.820 -66.030 92.610 ;
        RECT -64.590 92.460 -64.250 92.610 ;
        RECT -61.890 92.610 -59.950 92.760 ;
        RECT -61.890 92.460 -61.550 92.610 ;
        RECT -64.570 92.260 -64.250 92.290 ;
        RECT -66.850 91.680 -66.030 91.820 ;
        RECT -65.070 92.120 -64.250 92.260 ;
        RECT -66.850 91.650 -66.530 91.680 ;
        RECT -69.550 91.330 -69.210 91.480 ;
        RECT -71.150 91.180 -69.210 91.330 ;
        RECT -66.850 91.330 -66.510 91.480 ;
        RECT -65.070 91.330 -64.910 92.120 ;
        RECT -64.570 92.010 -64.250 92.120 ;
        RECT -61.890 92.260 -61.570 92.290 ;
        RECT -61.890 92.120 -61.070 92.260 ;
        RECT -61.890 92.010 -61.570 92.120 ;
        RECT -66.850 91.180 -64.910 91.330 ;
        RECT -61.230 91.330 -61.070 92.120 ;
        RECT -60.110 91.820 -59.950 92.610 ;
        RECT -56.270 92.610 -54.330 92.760 ;
        RECT -59.610 91.820 -59.290 91.930 ;
        RECT -60.110 91.680 -59.290 91.820 ;
        RECT -59.610 91.650 -59.290 91.680 ;
        RECT -56.930 91.820 -56.610 91.930 ;
        RECT -56.270 91.820 -56.110 92.610 ;
        RECT -54.670 92.460 -54.330 92.610 ;
        RECT -51.970 92.610 -50.030 92.760 ;
        RECT -51.970 92.460 -51.630 92.610 ;
        RECT -54.650 92.260 -54.330 92.290 ;
        RECT -56.930 91.680 -56.110 91.820 ;
        RECT -55.150 92.120 -54.330 92.260 ;
        RECT -56.930 91.650 -56.610 91.680 ;
        RECT -59.630 91.330 -59.290 91.480 ;
        RECT -61.230 91.180 -59.290 91.330 ;
        RECT -56.930 91.330 -56.590 91.480 ;
        RECT -55.150 91.330 -54.990 92.120 ;
        RECT -54.650 92.010 -54.330 92.120 ;
        RECT -51.970 92.260 -51.650 92.290 ;
        RECT -51.970 92.120 -51.150 92.260 ;
        RECT -51.970 92.010 -51.650 92.120 ;
        RECT -56.930 91.180 -54.990 91.330 ;
        RECT -51.310 91.330 -51.150 92.120 ;
        RECT -50.190 91.820 -50.030 92.610 ;
        RECT -46.350 92.610 -44.410 92.760 ;
        RECT -49.690 91.820 -49.370 91.930 ;
        RECT -50.190 91.680 -49.370 91.820 ;
        RECT -49.690 91.650 -49.370 91.680 ;
        RECT -47.010 91.820 -46.690 91.930 ;
        RECT -46.350 91.820 -46.190 92.610 ;
        RECT -44.750 92.460 -44.410 92.610 ;
        RECT -42.050 92.610 -40.110 92.760 ;
        RECT -42.050 92.460 -41.710 92.610 ;
        RECT -44.730 92.260 -44.410 92.290 ;
        RECT -47.010 91.680 -46.190 91.820 ;
        RECT -45.230 92.120 -44.410 92.260 ;
        RECT -47.010 91.650 -46.690 91.680 ;
        RECT -49.710 91.330 -49.370 91.480 ;
        RECT -51.310 91.180 -49.370 91.330 ;
        RECT -47.010 91.330 -46.670 91.480 ;
        RECT -45.230 91.330 -45.070 92.120 ;
        RECT -44.730 92.010 -44.410 92.120 ;
        RECT -42.050 92.260 -41.730 92.290 ;
        RECT -42.050 92.120 -41.230 92.260 ;
        RECT -42.050 92.010 -41.730 92.120 ;
        RECT -47.010 91.180 -45.070 91.330 ;
        RECT -41.390 91.330 -41.230 92.120 ;
        RECT -40.270 91.820 -40.110 92.610 ;
        RECT -36.430 92.610 -34.490 92.760 ;
        RECT -39.770 91.820 -39.450 91.930 ;
        RECT -40.270 91.680 -39.450 91.820 ;
        RECT -39.770 91.650 -39.450 91.680 ;
        RECT -37.090 91.820 -36.770 91.930 ;
        RECT -36.430 91.820 -36.270 92.610 ;
        RECT -34.830 92.460 -34.490 92.610 ;
        RECT -32.130 92.610 -30.190 92.760 ;
        RECT -32.130 92.460 -31.790 92.610 ;
        RECT -34.810 92.260 -34.490 92.290 ;
        RECT -37.090 91.680 -36.270 91.820 ;
        RECT -35.310 92.120 -34.490 92.260 ;
        RECT -37.090 91.650 -36.770 91.680 ;
        RECT -39.790 91.330 -39.450 91.480 ;
        RECT -41.390 91.180 -39.450 91.330 ;
        RECT -37.090 91.330 -36.750 91.480 ;
        RECT -35.310 91.330 -35.150 92.120 ;
        RECT -34.810 92.010 -34.490 92.120 ;
        RECT -32.130 92.260 -31.810 92.290 ;
        RECT -32.130 92.120 -31.310 92.260 ;
        RECT -32.130 92.010 -31.810 92.120 ;
        RECT -37.090 91.180 -35.150 91.330 ;
        RECT -31.470 91.330 -31.310 92.120 ;
        RECT -30.350 91.820 -30.190 92.610 ;
        RECT -26.510 92.610 -24.570 92.760 ;
        RECT -29.850 91.820 -29.530 91.930 ;
        RECT -30.350 91.680 -29.530 91.820 ;
        RECT -29.850 91.650 -29.530 91.680 ;
        RECT -27.170 91.820 -26.850 91.930 ;
        RECT -26.510 91.820 -26.350 92.610 ;
        RECT -24.910 92.460 -24.570 92.610 ;
        RECT -22.210 92.610 -20.270 92.760 ;
        RECT -22.210 92.460 -21.870 92.610 ;
        RECT -24.890 92.260 -24.570 92.290 ;
        RECT -27.170 91.680 -26.350 91.820 ;
        RECT -25.390 92.120 -24.570 92.260 ;
        RECT -27.170 91.650 -26.850 91.680 ;
        RECT -29.870 91.330 -29.530 91.480 ;
        RECT -31.470 91.180 -29.530 91.330 ;
        RECT -27.170 91.330 -26.830 91.480 ;
        RECT -25.390 91.330 -25.230 92.120 ;
        RECT -24.890 92.010 -24.570 92.120 ;
        RECT -22.210 92.260 -21.890 92.290 ;
        RECT -22.210 92.120 -21.390 92.260 ;
        RECT -22.210 92.010 -21.890 92.120 ;
        RECT -27.170 91.180 -25.230 91.330 ;
        RECT -21.550 91.330 -21.390 92.120 ;
        RECT -20.430 91.820 -20.270 92.610 ;
        RECT -16.590 92.610 -14.650 92.760 ;
        RECT -19.930 91.820 -19.610 91.930 ;
        RECT -20.430 91.680 -19.610 91.820 ;
        RECT -19.930 91.650 -19.610 91.680 ;
        RECT -17.250 91.820 -16.930 91.930 ;
        RECT -16.590 91.820 -16.430 92.610 ;
        RECT -14.990 92.460 -14.650 92.610 ;
        RECT -12.290 92.610 -10.350 92.760 ;
        RECT -12.290 92.460 -11.950 92.610 ;
        RECT -14.970 92.260 -14.650 92.290 ;
        RECT -17.250 91.680 -16.430 91.820 ;
        RECT -15.470 92.120 -14.650 92.260 ;
        RECT -17.250 91.650 -16.930 91.680 ;
        RECT -19.950 91.330 -19.610 91.480 ;
        RECT -21.550 91.180 -19.610 91.330 ;
        RECT -17.250 91.330 -16.910 91.480 ;
        RECT -15.470 91.330 -15.310 92.120 ;
        RECT -14.970 92.010 -14.650 92.120 ;
        RECT -12.290 92.260 -11.970 92.290 ;
        RECT -12.290 92.120 -11.470 92.260 ;
        RECT -12.290 92.010 -11.970 92.120 ;
        RECT -17.250 91.180 -15.310 91.330 ;
        RECT -11.630 91.330 -11.470 92.120 ;
        RECT -10.510 91.820 -10.350 92.610 ;
        RECT -6.670 92.610 -4.730 92.760 ;
        RECT -10.010 91.820 -9.690 91.930 ;
        RECT -10.510 91.680 -9.690 91.820 ;
        RECT -10.010 91.650 -9.690 91.680 ;
        RECT -7.330 91.820 -7.010 91.930 ;
        RECT -6.670 91.820 -6.510 92.610 ;
        RECT -5.070 92.460 -4.730 92.610 ;
        RECT -2.370 92.610 -0.430 92.760 ;
        RECT -2.370 92.460 -2.030 92.610 ;
        RECT -5.050 92.260 -4.730 92.290 ;
        RECT -7.330 91.680 -6.510 91.820 ;
        RECT -5.550 92.120 -4.730 92.260 ;
        RECT -7.330 91.650 -7.010 91.680 ;
        RECT -10.030 91.330 -9.690 91.480 ;
        RECT -11.630 91.180 -9.690 91.330 ;
        RECT -7.330 91.330 -6.990 91.480 ;
        RECT -5.550 91.330 -5.390 92.120 ;
        RECT -5.050 92.010 -4.730 92.120 ;
        RECT -2.370 92.260 -2.050 92.290 ;
        RECT -2.370 92.120 -1.550 92.260 ;
        RECT -2.370 92.010 -2.050 92.120 ;
        RECT -7.330 91.180 -5.390 91.330 ;
        RECT -1.710 91.330 -1.550 92.120 ;
        RECT -0.590 91.820 -0.430 92.610 ;
        RECT 3.250 92.610 5.190 92.760 ;
        RECT -0.090 91.820 0.230 91.930 ;
        RECT -0.590 91.680 0.230 91.820 ;
        RECT -0.090 91.650 0.230 91.680 ;
        RECT 2.590 91.820 2.910 91.930 ;
        RECT 3.250 91.820 3.410 92.610 ;
        RECT 4.850 92.460 5.190 92.610 ;
        RECT 7.550 92.610 9.490 92.760 ;
        RECT 7.550 92.460 7.890 92.610 ;
        RECT 4.870 92.260 5.190 92.290 ;
        RECT 2.590 91.680 3.410 91.820 ;
        RECT 4.370 92.120 5.190 92.260 ;
        RECT 2.590 91.650 2.910 91.680 ;
        RECT -0.110 91.330 0.230 91.480 ;
        RECT -1.710 91.180 0.230 91.330 ;
        RECT 2.590 91.330 2.930 91.480 ;
        RECT 4.370 91.330 4.530 92.120 ;
        RECT 4.870 92.010 5.190 92.120 ;
        RECT 7.550 92.260 7.870 92.290 ;
        RECT 7.550 92.120 8.370 92.260 ;
        RECT 7.550 92.010 7.870 92.120 ;
        RECT 2.590 91.180 4.530 91.330 ;
        RECT 8.210 91.330 8.370 92.120 ;
        RECT 9.330 91.820 9.490 92.610 ;
        RECT 13.170 92.610 15.110 92.760 ;
        RECT 9.830 91.820 10.150 91.930 ;
        RECT 9.330 91.680 10.150 91.820 ;
        RECT 9.830 91.650 10.150 91.680 ;
        RECT 12.510 91.820 12.830 91.930 ;
        RECT 13.170 91.820 13.330 92.610 ;
        RECT 14.770 92.460 15.110 92.610 ;
        RECT 17.470 92.610 19.410 92.760 ;
        RECT 17.470 92.460 17.810 92.610 ;
        RECT 14.790 92.260 15.110 92.290 ;
        RECT 12.510 91.680 13.330 91.820 ;
        RECT 14.290 92.120 15.110 92.260 ;
        RECT 12.510 91.650 12.830 91.680 ;
        RECT 9.810 91.330 10.150 91.480 ;
        RECT 8.210 91.180 10.150 91.330 ;
        RECT 12.510 91.330 12.850 91.480 ;
        RECT 14.290 91.330 14.450 92.120 ;
        RECT 14.790 92.010 15.110 92.120 ;
        RECT 17.470 92.260 17.790 92.290 ;
        RECT 17.470 92.120 18.290 92.260 ;
        RECT 17.470 92.010 17.790 92.120 ;
        RECT 12.510 91.180 14.450 91.330 ;
        RECT 18.130 91.330 18.290 92.120 ;
        RECT 19.250 91.820 19.410 92.610 ;
        RECT 23.090 92.610 25.030 92.760 ;
        RECT 19.750 91.820 20.070 91.930 ;
        RECT 19.250 91.680 20.070 91.820 ;
        RECT 19.750 91.650 20.070 91.680 ;
        RECT 22.430 91.820 22.750 91.930 ;
        RECT 23.090 91.820 23.250 92.610 ;
        RECT 24.690 92.460 25.030 92.610 ;
        RECT 24.710 92.260 25.030 92.290 ;
        RECT 22.430 91.680 23.250 91.820 ;
        RECT 24.210 92.120 25.030 92.260 ;
        RECT 22.430 91.650 22.750 91.680 ;
        RECT 19.730 91.330 20.070 91.480 ;
        RECT 18.130 91.180 20.070 91.330 ;
        RECT 22.430 91.330 22.770 91.480 ;
        RECT 24.210 91.330 24.370 92.120 ;
        RECT 24.710 92.010 25.030 92.120 ;
        RECT 22.430 91.180 24.370 91.330 ;
        RECT -291.460 90.370 -289.620 90.850 ;
        RECT -289.700 89.280 -289.220 90.180 ;
        RECT -288.400 90.050 -288.210 91.180 ;
        RECT -284.330 90.050 -284.140 91.180 ;
        RECT -278.480 90.050 -278.290 91.180 ;
        RECT -274.410 90.050 -274.220 91.180 ;
        RECT -268.560 90.050 -268.370 91.180 ;
        RECT -264.490 90.050 -264.300 91.180 ;
        RECT -258.640 90.050 -258.450 91.180 ;
        RECT -254.570 90.050 -254.380 91.180 ;
        RECT -248.720 90.050 -248.530 91.180 ;
        RECT -244.650 90.050 -244.460 91.180 ;
        RECT -238.800 90.050 -238.610 91.180 ;
        RECT -234.730 90.050 -234.540 91.180 ;
        RECT -228.880 90.050 -228.690 91.180 ;
        RECT -224.810 90.050 -224.620 91.180 ;
        RECT -218.960 90.050 -218.770 91.180 ;
        RECT -214.890 90.050 -214.700 91.180 ;
        RECT -209.040 90.050 -208.850 91.180 ;
        RECT -204.970 90.050 -204.780 91.180 ;
        RECT -199.120 90.050 -198.930 91.180 ;
        RECT -195.050 90.050 -194.860 91.180 ;
        RECT -189.200 90.050 -189.010 91.180 ;
        RECT -185.130 90.050 -184.940 91.180 ;
        RECT -179.280 90.050 -179.090 91.180 ;
        RECT -175.210 90.050 -175.020 91.180 ;
        RECT -169.360 90.050 -169.170 91.180 ;
        RECT -165.290 90.050 -165.100 91.180 ;
        RECT -159.440 90.050 -159.250 91.180 ;
        RECT -155.370 90.050 -155.180 91.180 ;
        RECT -149.520 90.050 -149.330 91.180 ;
        RECT -145.450 90.050 -145.260 91.180 ;
        RECT -139.600 90.050 -139.410 91.180 ;
        RECT -135.530 90.050 -135.340 91.180 ;
        RECT -129.680 90.050 -129.490 91.180 ;
        RECT -125.610 90.050 -125.420 91.180 ;
        RECT -119.760 90.050 -119.570 91.180 ;
        RECT -115.690 90.050 -115.500 91.180 ;
        RECT -109.840 90.050 -109.650 91.180 ;
        RECT -105.770 90.050 -105.580 91.180 ;
        RECT -99.920 90.050 -99.730 91.180 ;
        RECT -95.850 90.050 -95.660 91.180 ;
        RECT -90.000 90.050 -89.810 91.180 ;
        RECT -85.930 90.050 -85.740 91.180 ;
        RECT -80.080 90.050 -79.890 91.180 ;
        RECT -76.010 90.050 -75.820 91.180 ;
        RECT -70.160 90.050 -69.970 91.180 ;
        RECT -66.090 90.050 -65.900 91.180 ;
        RECT -60.240 90.050 -60.050 91.180 ;
        RECT -56.170 90.050 -55.980 91.180 ;
        RECT -50.320 90.050 -50.130 91.180 ;
        RECT -46.250 90.050 -46.060 91.180 ;
        RECT -40.400 90.050 -40.210 91.180 ;
        RECT -36.330 90.050 -36.140 91.180 ;
        RECT -30.480 90.050 -30.290 91.180 ;
        RECT -26.410 90.050 -26.220 91.180 ;
        RECT -20.560 90.050 -20.370 91.180 ;
        RECT -16.490 90.050 -16.300 91.180 ;
        RECT -10.640 90.050 -10.450 91.180 ;
        RECT -6.570 90.050 -6.380 91.180 ;
        RECT -0.720 90.050 -0.530 91.180 ;
        RECT 3.350 90.050 3.540 91.180 ;
        RECT 9.200 90.050 9.390 91.180 ;
        RECT 13.270 90.050 13.460 91.180 ;
        RECT 19.120 90.050 19.310 91.180 ;
        RECT 23.190 90.050 23.380 91.180 ;
        RECT -288.450 89.760 -288.130 90.050 ;
        RECT -284.410 89.760 -284.090 90.050 ;
        RECT -278.530 89.760 -278.210 90.050 ;
        RECT -274.490 89.760 -274.170 90.050 ;
        RECT -268.610 89.760 -268.290 90.050 ;
        RECT -264.570 89.760 -264.250 90.050 ;
        RECT -258.690 89.760 -258.370 90.050 ;
        RECT -254.650 89.760 -254.330 90.050 ;
        RECT -248.770 89.760 -248.450 90.050 ;
        RECT -244.730 89.760 -244.410 90.050 ;
        RECT -238.850 89.760 -238.530 90.050 ;
        RECT -234.810 89.760 -234.490 90.050 ;
        RECT -228.930 89.760 -228.610 90.050 ;
        RECT -224.890 89.760 -224.570 90.050 ;
        RECT -219.010 89.760 -218.690 90.050 ;
        RECT -214.970 89.760 -214.650 90.050 ;
        RECT -209.090 89.760 -208.770 90.050 ;
        RECT -205.050 89.760 -204.730 90.050 ;
        RECT -199.170 89.760 -198.850 90.050 ;
        RECT -195.130 89.760 -194.810 90.050 ;
        RECT -189.250 89.760 -188.930 90.050 ;
        RECT -185.210 89.760 -184.890 90.050 ;
        RECT -179.330 89.760 -179.010 90.050 ;
        RECT -175.290 89.760 -174.970 90.050 ;
        RECT -169.410 89.760 -169.090 90.050 ;
        RECT -165.370 89.760 -165.050 90.050 ;
        RECT -159.490 89.760 -159.170 90.050 ;
        RECT -155.450 89.760 -155.130 90.050 ;
        RECT -149.570 89.760 -149.250 90.050 ;
        RECT -145.530 89.760 -145.210 90.050 ;
        RECT -139.650 89.760 -139.330 90.050 ;
        RECT -135.610 89.760 -135.290 90.050 ;
        RECT -129.730 89.760 -129.410 90.050 ;
        RECT -125.690 89.760 -125.370 90.050 ;
        RECT -119.810 89.760 -119.490 90.050 ;
        RECT -115.770 89.760 -115.450 90.050 ;
        RECT -109.890 89.760 -109.570 90.050 ;
        RECT -105.850 89.760 -105.530 90.050 ;
        RECT -99.970 89.760 -99.650 90.050 ;
        RECT -95.930 89.760 -95.610 90.050 ;
        RECT -90.050 89.760 -89.730 90.050 ;
        RECT -86.010 89.760 -85.690 90.050 ;
        RECT -80.130 89.760 -79.810 90.050 ;
        RECT -76.090 89.760 -75.770 90.050 ;
        RECT -70.210 89.760 -69.890 90.050 ;
        RECT -66.170 89.760 -65.850 90.050 ;
        RECT -60.290 89.760 -59.970 90.050 ;
        RECT -56.250 89.760 -55.930 90.050 ;
        RECT -50.370 89.760 -50.050 90.050 ;
        RECT -46.330 89.760 -46.010 90.050 ;
        RECT -40.450 89.760 -40.130 90.050 ;
        RECT -36.410 89.760 -36.090 90.050 ;
        RECT -30.530 89.760 -30.210 90.050 ;
        RECT -26.490 89.760 -26.170 90.050 ;
        RECT -20.610 89.760 -20.290 90.050 ;
        RECT -16.570 89.760 -16.250 90.050 ;
        RECT -10.690 89.760 -10.370 90.050 ;
        RECT -6.650 89.760 -6.330 90.050 ;
        RECT -0.770 89.760 -0.450 90.050 ;
        RECT 3.270 89.760 3.590 90.050 ;
        RECT 9.150 89.760 9.470 90.050 ;
        RECT 13.190 89.760 13.510 90.050 ;
        RECT 19.070 89.760 19.390 90.050 ;
        RECT 23.110 89.760 23.430 90.050 ;
        RECT -290.160 88.800 -289.220 89.280 ;
        RECT 24.200 89.280 24.680 90.180 ;
        RECT -285.150 88.880 -283.460 89.180 ;
        RECT -275.230 88.880 -273.540 89.180 ;
        RECT -265.310 88.880 -263.620 89.180 ;
        RECT -255.390 88.880 -253.700 89.180 ;
        RECT -245.470 88.880 -243.780 89.180 ;
        RECT -235.550 88.880 -233.860 89.180 ;
        RECT -225.630 88.880 -223.940 89.180 ;
        RECT -215.710 88.880 -214.020 89.180 ;
        RECT -205.790 88.880 -204.100 89.180 ;
        RECT -195.870 88.880 -194.180 89.180 ;
        RECT -185.950 88.880 -184.260 89.180 ;
        RECT -176.030 88.880 -174.340 89.180 ;
        RECT -166.110 88.880 -164.420 89.180 ;
        RECT -156.190 88.880 -154.500 89.180 ;
        RECT -146.270 88.880 -144.580 89.180 ;
        RECT -136.350 88.880 -134.660 89.180 ;
        RECT -126.430 88.880 -124.740 89.180 ;
        RECT -116.510 88.880 -114.820 89.180 ;
        RECT -106.590 88.880 -104.900 89.180 ;
        RECT -96.670 88.880 -94.980 89.180 ;
        RECT -86.750 88.880 -85.060 89.180 ;
        RECT -76.830 88.880 -75.140 89.180 ;
        RECT -66.910 88.880 -65.220 89.180 ;
        RECT -56.990 88.880 -55.300 89.180 ;
        RECT -47.070 88.880 -45.380 89.180 ;
        RECT -37.150 88.880 -35.460 89.180 ;
        RECT -27.230 88.880 -25.540 89.180 ;
        RECT -17.310 88.880 -15.620 89.180 ;
        RECT -7.390 88.880 -5.700 89.180 ;
        RECT 2.530 88.880 4.220 89.180 ;
        RECT 12.450 88.880 14.140 89.180 ;
        RECT 22.370 88.880 24.060 89.180 ;
        RECT -284.640 88.180 -283.640 88.880 ;
        RECT -274.720 88.180 -273.720 88.880 ;
        RECT -264.800 88.180 -263.800 88.880 ;
        RECT -254.880 88.180 -253.880 88.880 ;
        RECT -244.960 88.180 -243.960 88.880 ;
        RECT -235.040 88.180 -234.040 88.880 ;
        RECT -225.120 88.180 -224.120 88.880 ;
        RECT -215.200 88.180 -214.200 88.880 ;
        RECT -205.280 88.180 -204.280 88.880 ;
        RECT -195.360 88.180 -194.360 88.880 ;
        RECT -185.440 88.180 -184.440 88.880 ;
        RECT -175.520 88.180 -174.520 88.880 ;
        RECT -165.600 88.180 -164.600 88.880 ;
        RECT -155.680 88.180 -154.680 88.880 ;
        RECT -145.760 88.180 -144.760 88.880 ;
        RECT -135.840 88.180 -134.840 88.880 ;
        RECT -125.920 88.180 -124.920 88.880 ;
        RECT -116.000 88.180 -115.000 88.880 ;
        RECT -106.080 88.180 -105.080 88.880 ;
        RECT -96.160 88.180 -95.160 88.880 ;
        RECT -86.240 88.180 -85.240 88.880 ;
        RECT -76.320 88.180 -75.320 88.880 ;
        RECT -66.400 88.180 -65.400 88.880 ;
        RECT -56.480 88.180 -55.480 88.880 ;
        RECT -46.560 88.180 -45.560 88.880 ;
        RECT -36.640 88.180 -35.640 88.880 ;
        RECT -26.720 88.180 -25.720 88.880 ;
        RECT -16.800 88.180 -15.800 88.880 ;
        RECT -6.880 88.180 -5.880 88.880 ;
        RECT 3.040 88.180 4.040 88.880 ;
        RECT 12.960 88.180 13.960 88.880 ;
        RECT 22.880 88.180 23.880 88.880 ;
        RECT 24.200 88.800 25.140 89.280 ;
        RECT -293.480 11.090 -293.020 11.095 ;
        RECT -293.480 10.615 -292.540 11.090 ;
        RECT -291.620 11.010 -290.620 11.710 ;
        RECT -281.700 11.010 -280.700 11.710 ;
        RECT -271.780 11.010 -270.780 11.710 ;
        RECT -261.860 11.010 -260.860 11.710 ;
        RECT -251.940 11.010 -250.940 11.710 ;
        RECT -242.020 11.010 -241.020 11.710 ;
        RECT -232.100 11.010 -231.100 11.710 ;
        RECT -222.180 11.010 -221.180 11.710 ;
        RECT -212.260 11.010 -211.260 11.710 ;
        RECT -202.340 11.010 -201.340 11.710 ;
        RECT -192.420 11.010 -191.420 11.710 ;
        RECT -182.500 11.010 -181.500 11.710 ;
        RECT -172.580 11.010 -171.580 11.710 ;
        RECT -162.660 11.010 -161.660 11.710 ;
        RECT -152.740 11.010 -151.740 11.710 ;
        RECT -142.820 11.010 -141.820 11.710 ;
        RECT -132.900 11.010 -131.900 11.710 ;
        RECT -122.980 11.010 -121.980 11.710 ;
        RECT -113.060 11.010 -112.060 11.710 ;
        RECT -103.140 11.010 -102.140 11.710 ;
        RECT -93.220 11.010 -92.220 11.710 ;
        RECT -83.300 11.010 -82.300 11.710 ;
        RECT -73.380 11.010 -72.380 11.710 ;
        RECT -63.460 11.010 -62.460 11.710 ;
        RECT -53.540 11.010 -52.540 11.710 ;
        RECT -43.620 11.010 -42.620 11.710 ;
        RECT -33.700 11.010 -32.700 11.710 ;
        RECT -23.780 11.010 -22.780 11.710 ;
        RECT -13.860 11.010 -12.860 11.710 ;
        RECT -3.940 11.010 -2.940 11.710 ;
        RECT 5.980 11.010 6.980 11.710 ;
        RECT 15.900 11.010 16.900 11.710 ;
        RECT -292.130 10.710 -290.440 11.010 ;
        RECT -282.210 10.710 -280.520 11.010 ;
        RECT -272.290 10.710 -270.600 11.010 ;
        RECT -262.370 10.710 -260.680 11.010 ;
        RECT -252.450 10.710 -250.760 11.010 ;
        RECT -242.530 10.710 -240.840 11.010 ;
        RECT -232.610 10.710 -230.920 11.010 ;
        RECT -222.690 10.710 -221.000 11.010 ;
        RECT -212.770 10.710 -211.080 11.010 ;
        RECT -202.850 10.710 -201.160 11.010 ;
        RECT -192.930 10.710 -191.240 11.010 ;
        RECT -183.010 10.710 -181.320 11.010 ;
        RECT -173.090 10.710 -171.400 11.010 ;
        RECT -163.170 10.710 -161.480 11.010 ;
        RECT -153.250 10.710 -151.560 11.010 ;
        RECT -143.330 10.710 -141.640 11.010 ;
        RECT -133.410 10.710 -131.720 11.010 ;
        RECT -123.490 10.710 -121.800 11.010 ;
        RECT -113.570 10.710 -111.880 11.010 ;
        RECT -103.650 10.710 -101.960 11.010 ;
        RECT -93.730 10.710 -92.040 11.010 ;
        RECT -83.810 10.710 -82.120 11.010 ;
        RECT -73.890 10.710 -72.200 11.010 ;
        RECT -63.970 10.710 -62.280 11.010 ;
        RECT -54.050 10.710 -52.360 11.010 ;
        RECT -44.130 10.710 -42.440 11.010 ;
        RECT -34.210 10.710 -32.520 11.010 ;
        RECT -24.290 10.710 -22.600 11.010 ;
        RECT -14.370 10.710 -12.680 11.010 ;
        RECT -4.450 10.710 -2.760 11.010 ;
        RECT 5.470 10.710 7.160 11.010 ;
        RECT 15.390 10.710 17.080 11.010 ;
        RECT -293.020 9.710 -292.540 10.615 ;
        RECT -291.390 9.840 -291.070 10.130 ;
        RECT -285.510 9.840 -285.190 10.130 ;
        RECT -281.470 9.840 -281.150 10.130 ;
        RECT -275.590 9.840 -275.270 10.130 ;
        RECT -271.550 9.840 -271.230 10.130 ;
        RECT -265.670 9.840 -265.350 10.130 ;
        RECT -261.630 9.840 -261.310 10.130 ;
        RECT -255.750 9.840 -255.430 10.130 ;
        RECT -251.710 9.840 -251.390 10.130 ;
        RECT -245.830 9.840 -245.510 10.130 ;
        RECT -241.790 9.840 -241.470 10.130 ;
        RECT -235.910 9.840 -235.590 10.130 ;
        RECT -231.870 9.840 -231.550 10.130 ;
        RECT -225.990 9.840 -225.670 10.130 ;
        RECT -221.950 9.840 -221.630 10.130 ;
        RECT -216.070 9.840 -215.750 10.130 ;
        RECT -212.030 9.840 -211.710 10.130 ;
        RECT -206.150 9.840 -205.830 10.130 ;
        RECT -202.110 9.840 -201.790 10.130 ;
        RECT -196.230 9.840 -195.910 10.130 ;
        RECT -192.190 9.840 -191.870 10.130 ;
        RECT -186.310 9.840 -185.990 10.130 ;
        RECT -182.270 9.840 -181.950 10.130 ;
        RECT -176.390 9.840 -176.070 10.130 ;
        RECT -172.350 9.840 -172.030 10.130 ;
        RECT -166.470 9.840 -166.150 10.130 ;
        RECT -162.430 9.840 -162.110 10.130 ;
        RECT -156.550 9.840 -156.230 10.130 ;
        RECT -152.510 9.840 -152.190 10.130 ;
        RECT -146.630 9.840 -146.310 10.130 ;
        RECT -142.590 9.840 -142.270 10.130 ;
        RECT -136.710 9.840 -136.390 10.130 ;
        RECT -132.670 9.840 -132.350 10.130 ;
        RECT -126.790 9.840 -126.470 10.130 ;
        RECT -122.750 9.840 -122.430 10.130 ;
        RECT -116.870 9.840 -116.550 10.130 ;
        RECT -112.830 9.840 -112.510 10.130 ;
        RECT -106.950 9.840 -106.630 10.130 ;
        RECT -102.910 9.840 -102.590 10.130 ;
        RECT -97.030 9.840 -96.710 10.130 ;
        RECT -92.990 9.840 -92.670 10.130 ;
        RECT -87.110 9.840 -86.790 10.130 ;
        RECT -83.070 9.840 -82.750 10.130 ;
        RECT -77.190 9.840 -76.870 10.130 ;
        RECT -73.150 9.840 -72.830 10.130 ;
        RECT -67.270 9.840 -66.950 10.130 ;
        RECT -63.230 9.840 -62.910 10.130 ;
        RECT -57.350 9.840 -57.030 10.130 ;
        RECT -53.310 9.840 -52.990 10.130 ;
        RECT -47.430 9.840 -47.110 10.130 ;
        RECT -43.390 9.840 -43.070 10.130 ;
        RECT -37.510 9.840 -37.190 10.130 ;
        RECT -33.470 9.840 -33.150 10.130 ;
        RECT -27.590 9.840 -27.270 10.130 ;
        RECT -23.550 9.840 -23.230 10.130 ;
        RECT -17.670 9.840 -17.350 10.130 ;
        RECT -13.630 9.840 -13.310 10.130 ;
        RECT -7.750 9.840 -7.430 10.130 ;
        RECT -3.710 9.840 -3.390 10.130 ;
        RECT 2.170 9.840 2.490 10.130 ;
        RECT 6.210 9.840 6.530 10.130 ;
        RECT 12.090 9.840 12.410 10.130 ;
        RECT 16.130 9.840 16.450 10.130 ;
        RECT 22.010 9.840 22.330 10.130 ;
        RECT -293.480 9.040 -291.640 9.520 ;
        RECT -291.310 8.710 -291.120 9.840 ;
        RECT -285.460 8.710 -285.270 9.840 ;
        RECT -281.390 8.710 -281.200 9.840 ;
        RECT -275.540 8.710 -275.350 9.840 ;
        RECT -271.470 8.710 -271.280 9.840 ;
        RECT -265.620 8.710 -265.430 9.840 ;
        RECT -261.550 8.710 -261.360 9.840 ;
        RECT -255.700 8.710 -255.510 9.840 ;
        RECT -251.630 8.710 -251.440 9.840 ;
        RECT -245.780 8.710 -245.590 9.840 ;
        RECT -241.710 8.710 -241.520 9.840 ;
        RECT -235.860 8.710 -235.670 9.840 ;
        RECT -231.790 8.710 -231.600 9.840 ;
        RECT -225.940 8.710 -225.750 9.840 ;
        RECT -221.870 8.710 -221.680 9.840 ;
        RECT -216.020 8.710 -215.830 9.840 ;
        RECT -211.950 8.710 -211.760 9.840 ;
        RECT -206.100 8.710 -205.910 9.840 ;
        RECT -202.030 8.710 -201.840 9.840 ;
        RECT -196.180 8.710 -195.990 9.840 ;
        RECT -192.110 8.710 -191.920 9.840 ;
        RECT -186.260 8.710 -186.070 9.840 ;
        RECT -182.190 8.710 -182.000 9.840 ;
        RECT -176.340 8.710 -176.150 9.840 ;
        RECT -172.270 8.710 -172.080 9.840 ;
        RECT -166.420 8.710 -166.230 9.840 ;
        RECT -162.350 8.710 -162.160 9.840 ;
        RECT -156.500 8.710 -156.310 9.840 ;
        RECT -152.430 8.710 -152.240 9.840 ;
        RECT -146.580 8.710 -146.390 9.840 ;
        RECT -142.510 8.710 -142.320 9.840 ;
        RECT -136.660 8.710 -136.470 9.840 ;
        RECT -132.590 8.710 -132.400 9.840 ;
        RECT -126.740 8.710 -126.550 9.840 ;
        RECT -122.670 8.710 -122.480 9.840 ;
        RECT -116.820 8.710 -116.630 9.840 ;
        RECT -112.750 8.710 -112.560 9.840 ;
        RECT -106.900 8.710 -106.710 9.840 ;
        RECT -102.830 8.710 -102.640 9.840 ;
        RECT -96.980 8.710 -96.790 9.840 ;
        RECT -92.910 8.710 -92.720 9.840 ;
        RECT -87.060 8.710 -86.870 9.840 ;
        RECT -82.990 8.710 -82.800 9.840 ;
        RECT -77.140 8.710 -76.950 9.840 ;
        RECT -73.070 8.710 -72.880 9.840 ;
        RECT -67.220 8.710 -67.030 9.840 ;
        RECT -63.150 8.710 -62.960 9.840 ;
        RECT -57.300 8.710 -57.110 9.840 ;
        RECT -53.230 8.710 -53.040 9.840 ;
        RECT -47.380 8.710 -47.190 9.840 ;
        RECT -43.310 8.710 -43.120 9.840 ;
        RECT -37.460 8.710 -37.270 9.840 ;
        RECT -33.390 8.710 -33.200 9.840 ;
        RECT -27.540 8.710 -27.350 9.840 ;
        RECT -23.470 8.710 -23.280 9.840 ;
        RECT -17.620 8.710 -17.430 9.840 ;
        RECT -13.550 8.710 -13.360 9.840 ;
        RECT -7.700 8.710 -7.510 9.840 ;
        RECT -3.630 8.710 -3.440 9.840 ;
        RECT 2.220 8.710 2.410 9.840 ;
        RECT 6.290 8.710 6.480 9.840 ;
        RECT 12.140 8.710 12.330 9.840 ;
        RECT 16.210 8.710 16.400 9.840 ;
        RECT 22.060 8.710 22.250 9.840 ;
        RECT 22.580 9.040 24.420 9.520 ;
        RECT -292.070 8.560 -290.130 8.710 ;
        RECT -292.070 8.410 -291.730 8.560 ;
        RECT -292.070 8.210 -291.750 8.240 ;
        RECT -292.070 8.070 -291.250 8.210 ;
        RECT -292.070 7.960 -291.750 8.070 ;
        RECT -291.410 7.280 -291.250 8.070 ;
        RECT -290.290 7.770 -290.130 8.560 ;
        RECT -286.450 8.560 -284.510 8.710 ;
        RECT -289.790 7.770 -289.470 7.880 ;
        RECT -290.290 7.630 -289.470 7.770 ;
        RECT -289.790 7.600 -289.470 7.630 ;
        RECT -287.110 7.770 -286.790 7.880 ;
        RECT -286.450 7.770 -286.290 8.560 ;
        RECT -284.850 8.410 -284.510 8.560 ;
        RECT -282.150 8.560 -280.210 8.710 ;
        RECT -282.150 8.410 -281.810 8.560 ;
        RECT -284.830 8.210 -284.510 8.240 ;
        RECT -287.110 7.630 -286.290 7.770 ;
        RECT -285.330 8.070 -284.510 8.210 ;
        RECT -287.110 7.600 -286.790 7.630 ;
        RECT -289.810 7.280 -289.470 7.430 ;
        RECT -291.410 7.130 -289.470 7.280 ;
        RECT -287.110 7.280 -286.770 7.430 ;
        RECT -285.330 7.280 -285.170 8.070 ;
        RECT -284.830 7.960 -284.510 8.070 ;
        RECT -282.150 8.210 -281.830 8.240 ;
        RECT -282.150 8.070 -281.330 8.210 ;
        RECT -282.150 7.960 -281.830 8.070 ;
        RECT -287.110 7.130 -285.170 7.280 ;
        RECT -281.490 7.280 -281.330 8.070 ;
        RECT -280.370 7.770 -280.210 8.560 ;
        RECT -276.530 8.560 -274.590 8.710 ;
        RECT -279.870 7.770 -279.550 7.880 ;
        RECT -280.370 7.630 -279.550 7.770 ;
        RECT -279.870 7.600 -279.550 7.630 ;
        RECT -277.190 7.770 -276.870 7.880 ;
        RECT -276.530 7.770 -276.370 8.560 ;
        RECT -274.930 8.410 -274.590 8.560 ;
        RECT -272.230 8.560 -270.290 8.710 ;
        RECT -272.230 8.410 -271.890 8.560 ;
        RECT -274.910 8.210 -274.590 8.240 ;
        RECT -277.190 7.630 -276.370 7.770 ;
        RECT -275.410 8.070 -274.590 8.210 ;
        RECT -277.190 7.600 -276.870 7.630 ;
        RECT -279.890 7.280 -279.550 7.430 ;
        RECT -281.490 7.130 -279.550 7.280 ;
        RECT -277.190 7.280 -276.850 7.430 ;
        RECT -275.410 7.280 -275.250 8.070 ;
        RECT -274.910 7.960 -274.590 8.070 ;
        RECT -272.230 8.210 -271.910 8.240 ;
        RECT -272.230 8.070 -271.410 8.210 ;
        RECT -272.230 7.960 -271.910 8.070 ;
        RECT -277.190 7.130 -275.250 7.280 ;
        RECT -271.570 7.280 -271.410 8.070 ;
        RECT -270.450 7.770 -270.290 8.560 ;
        RECT -266.610 8.560 -264.670 8.710 ;
        RECT -269.950 7.770 -269.630 7.880 ;
        RECT -270.450 7.630 -269.630 7.770 ;
        RECT -269.950 7.600 -269.630 7.630 ;
        RECT -267.270 7.770 -266.950 7.880 ;
        RECT -266.610 7.770 -266.450 8.560 ;
        RECT -265.010 8.410 -264.670 8.560 ;
        RECT -262.310 8.560 -260.370 8.710 ;
        RECT -262.310 8.410 -261.970 8.560 ;
        RECT -264.990 8.210 -264.670 8.240 ;
        RECT -267.270 7.630 -266.450 7.770 ;
        RECT -265.490 8.070 -264.670 8.210 ;
        RECT -267.270 7.600 -266.950 7.630 ;
        RECT -269.970 7.280 -269.630 7.430 ;
        RECT -271.570 7.130 -269.630 7.280 ;
        RECT -267.270 7.280 -266.930 7.430 ;
        RECT -265.490 7.280 -265.330 8.070 ;
        RECT -264.990 7.960 -264.670 8.070 ;
        RECT -262.310 8.210 -261.990 8.240 ;
        RECT -262.310 8.070 -261.490 8.210 ;
        RECT -262.310 7.960 -261.990 8.070 ;
        RECT -267.270 7.130 -265.330 7.280 ;
        RECT -261.650 7.280 -261.490 8.070 ;
        RECT -260.530 7.770 -260.370 8.560 ;
        RECT -256.690 8.560 -254.750 8.710 ;
        RECT -260.030 7.770 -259.710 7.880 ;
        RECT -260.530 7.630 -259.710 7.770 ;
        RECT -260.030 7.600 -259.710 7.630 ;
        RECT -257.350 7.770 -257.030 7.880 ;
        RECT -256.690 7.770 -256.530 8.560 ;
        RECT -255.090 8.410 -254.750 8.560 ;
        RECT -252.390 8.560 -250.450 8.710 ;
        RECT -252.390 8.410 -252.050 8.560 ;
        RECT -255.070 8.210 -254.750 8.240 ;
        RECT -257.350 7.630 -256.530 7.770 ;
        RECT -255.570 8.070 -254.750 8.210 ;
        RECT -257.350 7.600 -257.030 7.630 ;
        RECT -260.050 7.280 -259.710 7.430 ;
        RECT -261.650 7.130 -259.710 7.280 ;
        RECT -257.350 7.280 -257.010 7.430 ;
        RECT -255.570 7.280 -255.410 8.070 ;
        RECT -255.070 7.960 -254.750 8.070 ;
        RECT -252.390 8.210 -252.070 8.240 ;
        RECT -252.390 8.070 -251.570 8.210 ;
        RECT -252.390 7.960 -252.070 8.070 ;
        RECT -257.350 7.130 -255.410 7.280 ;
        RECT -251.730 7.280 -251.570 8.070 ;
        RECT -250.610 7.770 -250.450 8.560 ;
        RECT -246.770 8.560 -244.830 8.710 ;
        RECT -250.110 7.770 -249.790 7.880 ;
        RECT -250.610 7.630 -249.790 7.770 ;
        RECT -250.110 7.600 -249.790 7.630 ;
        RECT -247.430 7.770 -247.110 7.880 ;
        RECT -246.770 7.770 -246.610 8.560 ;
        RECT -245.170 8.410 -244.830 8.560 ;
        RECT -242.470 8.560 -240.530 8.710 ;
        RECT -242.470 8.410 -242.130 8.560 ;
        RECT -245.150 8.210 -244.830 8.240 ;
        RECT -247.430 7.630 -246.610 7.770 ;
        RECT -245.650 8.070 -244.830 8.210 ;
        RECT -247.430 7.600 -247.110 7.630 ;
        RECT -250.130 7.280 -249.790 7.430 ;
        RECT -251.730 7.130 -249.790 7.280 ;
        RECT -247.430 7.280 -247.090 7.430 ;
        RECT -245.650 7.280 -245.490 8.070 ;
        RECT -245.150 7.960 -244.830 8.070 ;
        RECT -242.470 8.210 -242.150 8.240 ;
        RECT -242.470 8.070 -241.650 8.210 ;
        RECT -242.470 7.960 -242.150 8.070 ;
        RECT -247.430 7.130 -245.490 7.280 ;
        RECT -241.810 7.280 -241.650 8.070 ;
        RECT -240.690 7.770 -240.530 8.560 ;
        RECT -236.850 8.560 -234.910 8.710 ;
        RECT -240.190 7.770 -239.870 7.880 ;
        RECT -240.690 7.630 -239.870 7.770 ;
        RECT -240.190 7.600 -239.870 7.630 ;
        RECT -237.510 7.770 -237.190 7.880 ;
        RECT -236.850 7.770 -236.690 8.560 ;
        RECT -235.250 8.410 -234.910 8.560 ;
        RECT -232.550 8.560 -230.610 8.710 ;
        RECT -232.550 8.410 -232.210 8.560 ;
        RECT -235.230 8.210 -234.910 8.240 ;
        RECT -237.510 7.630 -236.690 7.770 ;
        RECT -235.730 8.070 -234.910 8.210 ;
        RECT -237.510 7.600 -237.190 7.630 ;
        RECT -240.210 7.280 -239.870 7.430 ;
        RECT -241.810 7.130 -239.870 7.280 ;
        RECT -237.510 7.280 -237.170 7.430 ;
        RECT -235.730 7.280 -235.570 8.070 ;
        RECT -235.230 7.960 -234.910 8.070 ;
        RECT -232.550 8.210 -232.230 8.240 ;
        RECT -232.550 8.070 -231.730 8.210 ;
        RECT -232.550 7.960 -232.230 8.070 ;
        RECT -237.510 7.130 -235.570 7.280 ;
        RECT -231.890 7.280 -231.730 8.070 ;
        RECT -230.770 7.770 -230.610 8.560 ;
        RECT -226.930 8.560 -224.990 8.710 ;
        RECT -230.270 7.770 -229.950 7.880 ;
        RECT -230.770 7.630 -229.950 7.770 ;
        RECT -230.270 7.600 -229.950 7.630 ;
        RECT -227.590 7.770 -227.270 7.880 ;
        RECT -226.930 7.770 -226.770 8.560 ;
        RECT -225.330 8.410 -224.990 8.560 ;
        RECT -222.630 8.560 -220.690 8.710 ;
        RECT -222.630 8.410 -222.290 8.560 ;
        RECT -225.310 8.210 -224.990 8.240 ;
        RECT -227.590 7.630 -226.770 7.770 ;
        RECT -225.810 8.070 -224.990 8.210 ;
        RECT -227.590 7.600 -227.270 7.630 ;
        RECT -230.290 7.280 -229.950 7.430 ;
        RECT -231.890 7.130 -229.950 7.280 ;
        RECT -227.590 7.280 -227.250 7.430 ;
        RECT -225.810 7.280 -225.650 8.070 ;
        RECT -225.310 7.960 -224.990 8.070 ;
        RECT -222.630 8.210 -222.310 8.240 ;
        RECT -222.630 8.070 -221.810 8.210 ;
        RECT -222.630 7.960 -222.310 8.070 ;
        RECT -227.590 7.130 -225.650 7.280 ;
        RECT -221.970 7.280 -221.810 8.070 ;
        RECT -220.850 7.770 -220.690 8.560 ;
        RECT -217.010 8.560 -215.070 8.710 ;
        RECT -220.350 7.770 -220.030 7.880 ;
        RECT -220.850 7.630 -220.030 7.770 ;
        RECT -220.350 7.600 -220.030 7.630 ;
        RECT -217.670 7.770 -217.350 7.880 ;
        RECT -217.010 7.770 -216.850 8.560 ;
        RECT -215.410 8.410 -215.070 8.560 ;
        RECT -212.710 8.560 -210.770 8.710 ;
        RECT -212.710 8.410 -212.370 8.560 ;
        RECT -215.390 8.210 -215.070 8.240 ;
        RECT -217.670 7.630 -216.850 7.770 ;
        RECT -215.890 8.070 -215.070 8.210 ;
        RECT -217.670 7.600 -217.350 7.630 ;
        RECT -220.370 7.280 -220.030 7.430 ;
        RECT -221.970 7.130 -220.030 7.280 ;
        RECT -217.670 7.280 -217.330 7.430 ;
        RECT -215.890 7.280 -215.730 8.070 ;
        RECT -215.390 7.960 -215.070 8.070 ;
        RECT -212.710 8.210 -212.390 8.240 ;
        RECT -212.710 8.070 -211.890 8.210 ;
        RECT -212.710 7.960 -212.390 8.070 ;
        RECT -217.670 7.130 -215.730 7.280 ;
        RECT -212.050 7.280 -211.890 8.070 ;
        RECT -210.930 7.770 -210.770 8.560 ;
        RECT -207.090 8.560 -205.150 8.710 ;
        RECT -210.430 7.770 -210.110 7.880 ;
        RECT -210.930 7.630 -210.110 7.770 ;
        RECT -210.430 7.600 -210.110 7.630 ;
        RECT -207.750 7.770 -207.430 7.880 ;
        RECT -207.090 7.770 -206.930 8.560 ;
        RECT -205.490 8.410 -205.150 8.560 ;
        RECT -202.790 8.560 -200.850 8.710 ;
        RECT -202.790 8.410 -202.450 8.560 ;
        RECT -205.470 8.210 -205.150 8.240 ;
        RECT -207.750 7.630 -206.930 7.770 ;
        RECT -205.970 8.070 -205.150 8.210 ;
        RECT -207.750 7.600 -207.430 7.630 ;
        RECT -210.450 7.280 -210.110 7.430 ;
        RECT -212.050 7.130 -210.110 7.280 ;
        RECT -207.750 7.280 -207.410 7.430 ;
        RECT -205.970 7.280 -205.810 8.070 ;
        RECT -205.470 7.960 -205.150 8.070 ;
        RECT -202.790 8.210 -202.470 8.240 ;
        RECT -202.790 8.070 -201.970 8.210 ;
        RECT -202.790 7.960 -202.470 8.070 ;
        RECT -207.750 7.130 -205.810 7.280 ;
        RECT -202.130 7.280 -201.970 8.070 ;
        RECT -201.010 7.770 -200.850 8.560 ;
        RECT -197.170 8.560 -195.230 8.710 ;
        RECT -200.510 7.770 -200.190 7.880 ;
        RECT -201.010 7.630 -200.190 7.770 ;
        RECT -200.510 7.600 -200.190 7.630 ;
        RECT -197.830 7.770 -197.510 7.880 ;
        RECT -197.170 7.770 -197.010 8.560 ;
        RECT -195.570 8.410 -195.230 8.560 ;
        RECT -192.870 8.560 -190.930 8.710 ;
        RECT -192.870 8.410 -192.530 8.560 ;
        RECT -195.550 8.210 -195.230 8.240 ;
        RECT -197.830 7.630 -197.010 7.770 ;
        RECT -196.050 8.070 -195.230 8.210 ;
        RECT -197.830 7.600 -197.510 7.630 ;
        RECT -200.530 7.280 -200.190 7.430 ;
        RECT -202.130 7.130 -200.190 7.280 ;
        RECT -197.830 7.280 -197.490 7.430 ;
        RECT -196.050 7.280 -195.890 8.070 ;
        RECT -195.550 7.960 -195.230 8.070 ;
        RECT -192.870 8.210 -192.550 8.240 ;
        RECT -192.870 8.070 -192.050 8.210 ;
        RECT -192.870 7.960 -192.550 8.070 ;
        RECT -197.830 7.130 -195.890 7.280 ;
        RECT -192.210 7.280 -192.050 8.070 ;
        RECT -191.090 7.770 -190.930 8.560 ;
        RECT -187.250 8.560 -185.310 8.710 ;
        RECT -190.590 7.770 -190.270 7.880 ;
        RECT -191.090 7.630 -190.270 7.770 ;
        RECT -190.590 7.600 -190.270 7.630 ;
        RECT -187.910 7.770 -187.590 7.880 ;
        RECT -187.250 7.770 -187.090 8.560 ;
        RECT -185.650 8.410 -185.310 8.560 ;
        RECT -182.950 8.560 -181.010 8.710 ;
        RECT -182.950 8.410 -182.610 8.560 ;
        RECT -185.630 8.210 -185.310 8.240 ;
        RECT -187.910 7.630 -187.090 7.770 ;
        RECT -186.130 8.070 -185.310 8.210 ;
        RECT -187.910 7.600 -187.590 7.630 ;
        RECT -190.610 7.280 -190.270 7.430 ;
        RECT -192.210 7.130 -190.270 7.280 ;
        RECT -187.910 7.280 -187.570 7.430 ;
        RECT -186.130 7.280 -185.970 8.070 ;
        RECT -185.630 7.960 -185.310 8.070 ;
        RECT -182.950 8.210 -182.630 8.240 ;
        RECT -182.950 8.070 -182.130 8.210 ;
        RECT -182.950 7.960 -182.630 8.070 ;
        RECT -187.910 7.130 -185.970 7.280 ;
        RECT -182.290 7.280 -182.130 8.070 ;
        RECT -181.170 7.770 -181.010 8.560 ;
        RECT -177.330 8.560 -175.390 8.710 ;
        RECT -180.670 7.770 -180.350 7.880 ;
        RECT -181.170 7.630 -180.350 7.770 ;
        RECT -180.670 7.600 -180.350 7.630 ;
        RECT -177.990 7.770 -177.670 7.880 ;
        RECT -177.330 7.770 -177.170 8.560 ;
        RECT -175.730 8.410 -175.390 8.560 ;
        RECT -173.030 8.560 -171.090 8.710 ;
        RECT -173.030 8.410 -172.690 8.560 ;
        RECT -175.710 8.210 -175.390 8.240 ;
        RECT -177.990 7.630 -177.170 7.770 ;
        RECT -176.210 8.070 -175.390 8.210 ;
        RECT -177.990 7.600 -177.670 7.630 ;
        RECT -180.690 7.280 -180.350 7.430 ;
        RECT -182.290 7.130 -180.350 7.280 ;
        RECT -177.990 7.280 -177.650 7.430 ;
        RECT -176.210 7.280 -176.050 8.070 ;
        RECT -175.710 7.960 -175.390 8.070 ;
        RECT -173.030 8.210 -172.710 8.240 ;
        RECT -173.030 8.070 -172.210 8.210 ;
        RECT -173.030 7.960 -172.710 8.070 ;
        RECT -177.990 7.130 -176.050 7.280 ;
        RECT -172.370 7.280 -172.210 8.070 ;
        RECT -171.250 7.770 -171.090 8.560 ;
        RECT -167.410 8.560 -165.470 8.710 ;
        RECT -170.750 7.770 -170.430 7.880 ;
        RECT -171.250 7.630 -170.430 7.770 ;
        RECT -170.750 7.600 -170.430 7.630 ;
        RECT -168.070 7.770 -167.750 7.880 ;
        RECT -167.410 7.770 -167.250 8.560 ;
        RECT -165.810 8.410 -165.470 8.560 ;
        RECT -163.110 8.560 -161.170 8.710 ;
        RECT -163.110 8.410 -162.770 8.560 ;
        RECT -165.790 8.210 -165.470 8.240 ;
        RECT -168.070 7.630 -167.250 7.770 ;
        RECT -166.290 8.070 -165.470 8.210 ;
        RECT -168.070 7.600 -167.750 7.630 ;
        RECT -170.770 7.280 -170.430 7.430 ;
        RECT -172.370 7.130 -170.430 7.280 ;
        RECT -168.070 7.280 -167.730 7.430 ;
        RECT -166.290 7.280 -166.130 8.070 ;
        RECT -165.790 7.960 -165.470 8.070 ;
        RECT -163.110 8.210 -162.790 8.240 ;
        RECT -163.110 8.070 -162.290 8.210 ;
        RECT -163.110 7.960 -162.790 8.070 ;
        RECT -168.070 7.130 -166.130 7.280 ;
        RECT -162.450 7.280 -162.290 8.070 ;
        RECT -161.330 7.770 -161.170 8.560 ;
        RECT -157.490 8.560 -155.550 8.710 ;
        RECT -160.830 7.770 -160.510 7.880 ;
        RECT -161.330 7.630 -160.510 7.770 ;
        RECT -160.830 7.600 -160.510 7.630 ;
        RECT -158.150 7.770 -157.830 7.880 ;
        RECT -157.490 7.770 -157.330 8.560 ;
        RECT -155.890 8.410 -155.550 8.560 ;
        RECT -153.190 8.560 -151.250 8.710 ;
        RECT -153.190 8.410 -152.850 8.560 ;
        RECT -155.870 8.210 -155.550 8.240 ;
        RECT -158.150 7.630 -157.330 7.770 ;
        RECT -156.370 8.070 -155.550 8.210 ;
        RECT -158.150 7.600 -157.830 7.630 ;
        RECT -160.850 7.280 -160.510 7.430 ;
        RECT -162.450 7.130 -160.510 7.280 ;
        RECT -158.150 7.280 -157.810 7.430 ;
        RECT -156.370 7.280 -156.210 8.070 ;
        RECT -155.870 7.960 -155.550 8.070 ;
        RECT -153.190 8.210 -152.870 8.240 ;
        RECT -153.190 8.070 -152.370 8.210 ;
        RECT -153.190 7.960 -152.870 8.070 ;
        RECT -158.150 7.130 -156.210 7.280 ;
        RECT -152.530 7.280 -152.370 8.070 ;
        RECT -151.410 7.770 -151.250 8.560 ;
        RECT -147.570 8.560 -145.630 8.710 ;
        RECT -150.910 7.770 -150.590 7.880 ;
        RECT -151.410 7.630 -150.590 7.770 ;
        RECT -150.910 7.600 -150.590 7.630 ;
        RECT -148.230 7.770 -147.910 7.880 ;
        RECT -147.570 7.770 -147.410 8.560 ;
        RECT -145.970 8.410 -145.630 8.560 ;
        RECT -143.270 8.560 -141.330 8.710 ;
        RECT -143.270 8.410 -142.930 8.560 ;
        RECT -145.950 8.210 -145.630 8.240 ;
        RECT -148.230 7.630 -147.410 7.770 ;
        RECT -146.450 8.070 -145.630 8.210 ;
        RECT -148.230 7.600 -147.910 7.630 ;
        RECT -150.930 7.280 -150.590 7.430 ;
        RECT -152.530 7.130 -150.590 7.280 ;
        RECT -148.230 7.280 -147.890 7.430 ;
        RECT -146.450 7.280 -146.290 8.070 ;
        RECT -145.950 7.960 -145.630 8.070 ;
        RECT -143.270 8.210 -142.950 8.240 ;
        RECT -143.270 8.070 -142.450 8.210 ;
        RECT -143.270 7.960 -142.950 8.070 ;
        RECT -148.230 7.130 -146.290 7.280 ;
        RECT -142.610 7.280 -142.450 8.070 ;
        RECT -141.490 7.770 -141.330 8.560 ;
        RECT -137.650 8.560 -135.710 8.710 ;
        RECT -140.990 7.770 -140.670 7.880 ;
        RECT -141.490 7.630 -140.670 7.770 ;
        RECT -140.990 7.600 -140.670 7.630 ;
        RECT -138.310 7.770 -137.990 7.880 ;
        RECT -137.650 7.770 -137.490 8.560 ;
        RECT -136.050 8.410 -135.710 8.560 ;
        RECT -133.350 8.560 -131.410 8.710 ;
        RECT -133.350 8.410 -133.010 8.560 ;
        RECT -136.030 8.210 -135.710 8.240 ;
        RECT -138.310 7.630 -137.490 7.770 ;
        RECT -136.530 8.070 -135.710 8.210 ;
        RECT -138.310 7.600 -137.990 7.630 ;
        RECT -141.010 7.280 -140.670 7.430 ;
        RECT -142.610 7.130 -140.670 7.280 ;
        RECT -138.310 7.280 -137.970 7.430 ;
        RECT -136.530 7.280 -136.370 8.070 ;
        RECT -136.030 7.960 -135.710 8.070 ;
        RECT -133.350 8.210 -133.030 8.240 ;
        RECT -133.350 8.070 -132.530 8.210 ;
        RECT -133.350 7.960 -133.030 8.070 ;
        RECT -138.310 7.130 -136.370 7.280 ;
        RECT -132.690 7.280 -132.530 8.070 ;
        RECT -131.570 7.770 -131.410 8.560 ;
        RECT -127.730 8.560 -125.790 8.710 ;
        RECT -131.070 7.770 -130.750 7.880 ;
        RECT -131.570 7.630 -130.750 7.770 ;
        RECT -131.070 7.600 -130.750 7.630 ;
        RECT -128.390 7.770 -128.070 7.880 ;
        RECT -127.730 7.770 -127.570 8.560 ;
        RECT -126.130 8.410 -125.790 8.560 ;
        RECT -123.430 8.560 -121.490 8.710 ;
        RECT -123.430 8.410 -123.090 8.560 ;
        RECT -126.110 8.210 -125.790 8.240 ;
        RECT -128.390 7.630 -127.570 7.770 ;
        RECT -126.610 8.070 -125.790 8.210 ;
        RECT -128.390 7.600 -128.070 7.630 ;
        RECT -131.090 7.280 -130.750 7.430 ;
        RECT -132.690 7.130 -130.750 7.280 ;
        RECT -128.390 7.280 -128.050 7.430 ;
        RECT -126.610 7.280 -126.450 8.070 ;
        RECT -126.110 7.960 -125.790 8.070 ;
        RECT -123.430 8.210 -123.110 8.240 ;
        RECT -123.430 8.070 -122.610 8.210 ;
        RECT -123.430 7.960 -123.110 8.070 ;
        RECT -128.390 7.130 -126.450 7.280 ;
        RECT -122.770 7.280 -122.610 8.070 ;
        RECT -121.650 7.770 -121.490 8.560 ;
        RECT -117.810 8.560 -115.870 8.710 ;
        RECT -121.150 7.770 -120.830 7.880 ;
        RECT -121.650 7.630 -120.830 7.770 ;
        RECT -121.150 7.600 -120.830 7.630 ;
        RECT -118.470 7.770 -118.150 7.880 ;
        RECT -117.810 7.770 -117.650 8.560 ;
        RECT -116.210 8.410 -115.870 8.560 ;
        RECT -113.510 8.560 -111.570 8.710 ;
        RECT -113.510 8.410 -113.170 8.560 ;
        RECT -116.190 8.210 -115.870 8.240 ;
        RECT -118.470 7.630 -117.650 7.770 ;
        RECT -116.690 8.070 -115.870 8.210 ;
        RECT -118.470 7.600 -118.150 7.630 ;
        RECT -121.170 7.280 -120.830 7.430 ;
        RECT -122.770 7.130 -120.830 7.280 ;
        RECT -118.470 7.280 -118.130 7.430 ;
        RECT -116.690 7.280 -116.530 8.070 ;
        RECT -116.190 7.960 -115.870 8.070 ;
        RECT -113.510 8.210 -113.190 8.240 ;
        RECT -113.510 8.070 -112.690 8.210 ;
        RECT -113.510 7.960 -113.190 8.070 ;
        RECT -118.470 7.130 -116.530 7.280 ;
        RECT -112.850 7.280 -112.690 8.070 ;
        RECT -111.730 7.770 -111.570 8.560 ;
        RECT -107.890 8.560 -105.950 8.710 ;
        RECT -111.230 7.770 -110.910 7.880 ;
        RECT -111.730 7.630 -110.910 7.770 ;
        RECT -111.230 7.600 -110.910 7.630 ;
        RECT -108.550 7.770 -108.230 7.880 ;
        RECT -107.890 7.770 -107.730 8.560 ;
        RECT -106.290 8.410 -105.950 8.560 ;
        RECT -103.590 8.560 -101.650 8.710 ;
        RECT -103.590 8.410 -103.250 8.560 ;
        RECT -106.270 8.210 -105.950 8.240 ;
        RECT -108.550 7.630 -107.730 7.770 ;
        RECT -106.770 8.070 -105.950 8.210 ;
        RECT -108.550 7.600 -108.230 7.630 ;
        RECT -111.250 7.280 -110.910 7.430 ;
        RECT -112.850 7.130 -110.910 7.280 ;
        RECT -108.550 7.280 -108.210 7.430 ;
        RECT -106.770 7.280 -106.610 8.070 ;
        RECT -106.270 7.960 -105.950 8.070 ;
        RECT -103.590 8.210 -103.270 8.240 ;
        RECT -103.590 8.070 -102.770 8.210 ;
        RECT -103.590 7.960 -103.270 8.070 ;
        RECT -108.550 7.130 -106.610 7.280 ;
        RECT -102.930 7.280 -102.770 8.070 ;
        RECT -101.810 7.770 -101.650 8.560 ;
        RECT -97.970 8.560 -96.030 8.710 ;
        RECT -101.310 7.770 -100.990 7.880 ;
        RECT -101.810 7.630 -100.990 7.770 ;
        RECT -101.310 7.600 -100.990 7.630 ;
        RECT -98.630 7.770 -98.310 7.880 ;
        RECT -97.970 7.770 -97.810 8.560 ;
        RECT -96.370 8.410 -96.030 8.560 ;
        RECT -93.670 8.560 -91.730 8.710 ;
        RECT -93.670 8.410 -93.330 8.560 ;
        RECT -96.350 8.210 -96.030 8.240 ;
        RECT -98.630 7.630 -97.810 7.770 ;
        RECT -96.850 8.070 -96.030 8.210 ;
        RECT -98.630 7.600 -98.310 7.630 ;
        RECT -101.330 7.280 -100.990 7.430 ;
        RECT -102.930 7.130 -100.990 7.280 ;
        RECT -98.630 7.280 -98.290 7.430 ;
        RECT -96.850 7.280 -96.690 8.070 ;
        RECT -96.350 7.960 -96.030 8.070 ;
        RECT -93.670 8.210 -93.350 8.240 ;
        RECT -93.670 8.070 -92.850 8.210 ;
        RECT -93.670 7.960 -93.350 8.070 ;
        RECT -98.630 7.130 -96.690 7.280 ;
        RECT -93.010 7.280 -92.850 8.070 ;
        RECT -91.890 7.770 -91.730 8.560 ;
        RECT -88.050 8.560 -86.110 8.710 ;
        RECT -91.390 7.770 -91.070 7.880 ;
        RECT -91.890 7.630 -91.070 7.770 ;
        RECT -91.390 7.600 -91.070 7.630 ;
        RECT -88.710 7.770 -88.390 7.880 ;
        RECT -88.050 7.770 -87.890 8.560 ;
        RECT -86.450 8.410 -86.110 8.560 ;
        RECT -83.750 8.560 -81.810 8.710 ;
        RECT -83.750 8.410 -83.410 8.560 ;
        RECT -86.430 8.210 -86.110 8.240 ;
        RECT -88.710 7.630 -87.890 7.770 ;
        RECT -86.930 8.070 -86.110 8.210 ;
        RECT -88.710 7.600 -88.390 7.630 ;
        RECT -91.410 7.280 -91.070 7.430 ;
        RECT -93.010 7.130 -91.070 7.280 ;
        RECT -88.710 7.280 -88.370 7.430 ;
        RECT -86.930 7.280 -86.770 8.070 ;
        RECT -86.430 7.960 -86.110 8.070 ;
        RECT -83.750 8.210 -83.430 8.240 ;
        RECT -83.750 8.070 -82.930 8.210 ;
        RECT -83.750 7.960 -83.430 8.070 ;
        RECT -88.710 7.130 -86.770 7.280 ;
        RECT -83.090 7.280 -82.930 8.070 ;
        RECT -81.970 7.770 -81.810 8.560 ;
        RECT -78.130 8.560 -76.190 8.710 ;
        RECT -81.470 7.770 -81.150 7.880 ;
        RECT -81.970 7.630 -81.150 7.770 ;
        RECT -81.470 7.600 -81.150 7.630 ;
        RECT -78.790 7.770 -78.470 7.880 ;
        RECT -78.130 7.770 -77.970 8.560 ;
        RECT -76.530 8.410 -76.190 8.560 ;
        RECT -73.830 8.560 -71.890 8.710 ;
        RECT -73.830 8.410 -73.490 8.560 ;
        RECT -76.510 8.210 -76.190 8.240 ;
        RECT -78.790 7.630 -77.970 7.770 ;
        RECT -77.010 8.070 -76.190 8.210 ;
        RECT -78.790 7.600 -78.470 7.630 ;
        RECT -81.490 7.280 -81.150 7.430 ;
        RECT -83.090 7.130 -81.150 7.280 ;
        RECT -78.790 7.280 -78.450 7.430 ;
        RECT -77.010 7.280 -76.850 8.070 ;
        RECT -76.510 7.960 -76.190 8.070 ;
        RECT -73.830 8.210 -73.510 8.240 ;
        RECT -73.830 8.070 -73.010 8.210 ;
        RECT -73.830 7.960 -73.510 8.070 ;
        RECT -78.790 7.130 -76.850 7.280 ;
        RECT -73.170 7.280 -73.010 8.070 ;
        RECT -72.050 7.770 -71.890 8.560 ;
        RECT -68.210 8.560 -66.270 8.710 ;
        RECT -71.550 7.770 -71.230 7.880 ;
        RECT -72.050 7.630 -71.230 7.770 ;
        RECT -71.550 7.600 -71.230 7.630 ;
        RECT -68.870 7.770 -68.550 7.880 ;
        RECT -68.210 7.770 -68.050 8.560 ;
        RECT -66.610 8.410 -66.270 8.560 ;
        RECT -63.910 8.560 -61.970 8.710 ;
        RECT -63.910 8.410 -63.570 8.560 ;
        RECT -66.590 8.210 -66.270 8.240 ;
        RECT -68.870 7.630 -68.050 7.770 ;
        RECT -67.090 8.070 -66.270 8.210 ;
        RECT -68.870 7.600 -68.550 7.630 ;
        RECT -71.570 7.280 -71.230 7.430 ;
        RECT -73.170 7.130 -71.230 7.280 ;
        RECT -68.870 7.280 -68.530 7.430 ;
        RECT -67.090 7.280 -66.930 8.070 ;
        RECT -66.590 7.960 -66.270 8.070 ;
        RECT -63.910 8.210 -63.590 8.240 ;
        RECT -63.910 8.070 -63.090 8.210 ;
        RECT -63.910 7.960 -63.590 8.070 ;
        RECT -68.870 7.130 -66.930 7.280 ;
        RECT -63.250 7.280 -63.090 8.070 ;
        RECT -62.130 7.770 -61.970 8.560 ;
        RECT -58.290 8.560 -56.350 8.710 ;
        RECT -61.630 7.770 -61.310 7.880 ;
        RECT -62.130 7.630 -61.310 7.770 ;
        RECT -61.630 7.600 -61.310 7.630 ;
        RECT -58.950 7.770 -58.630 7.880 ;
        RECT -58.290 7.770 -58.130 8.560 ;
        RECT -56.690 8.410 -56.350 8.560 ;
        RECT -53.990 8.560 -52.050 8.710 ;
        RECT -53.990 8.410 -53.650 8.560 ;
        RECT -56.670 8.210 -56.350 8.240 ;
        RECT -58.950 7.630 -58.130 7.770 ;
        RECT -57.170 8.070 -56.350 8.210 ;
        RECT -58.950 7.600 -58.630 7.630 ;
        RECT -61.650 7.280 -61.310 7.430 ;
        RECT -63.250 7.130 -61.310 7.280 ;
        RECT -58.950 7.280 -58.610 7.430 ;
        RECT -57.170 7.280 -57.010 8.070 ;
        RECT -56.670 7.960 -56.350 8.070 ;
        RECT -53.990 8.210 -53.670 8.240 ;
        RECT -53.990 8.070 -53.170 8.210 ;
        RECT -53.990 7.960 -53.670 8.070 ;
        RECT -58.950 7.130 -57.010 7.280 ;
        RECT -53.330 7.280 -53.170 8.070 ;
        RECT -52.210 7.770 -52.050 8.560 ;
        RECT -48.370 8.560 -46.430 8.710 ;
        RECT -51.710 7.770 -51.390 7.880 ;
        RECT -52.210 7.630 -51.390 7.770 ;
        RECT -51.710 7.600 -51.390 7.630 ;
        RECT -49.030 7.770 -48.710 7.880 ;
        RECT -48.370 7.770 -48.210 8.560 ;
        RECT -46.770 8.410 -46.430 8.560 ;
        RECT -44.070 8.560 -42.130 8.710 ;
        RECT -44.070 8.410 -43.730 8.560 ;
        RECT -46.750 8.210 -46.430 8.240 ;
        RECT -49.030 7.630 -48.210 7.770 ;
        RECT -47.250 8.070 -46.430 8.210 ;
        RECT -49.030 7.600 -48.710 7.630 ;
        RECT -51.730 7.280 -51.390 7.430 ;
        RECT -53.330 7.130 -51.390 7.280 ;
        RECT -49.030 7.280 -48.690 7.430 ;
        RECT -47.250 7.280 -47.090 8.070 ;
        RECT -46.750 7.960 -46.430 8.070 ;
        RECT -44.070 8.210 -43.750 8.240 ;
        RECT -44.070 8.070 -43.250 8.210 ;
        RECT -44.070 7.960 -43.750 8.070 ;
        RECT -49.030 7.130 -47.090 7.280 ;
        RECT -43.410 7.280 -43.250 8.070 ;
        RECT -42.290 7.770 -42.130 8.560 ;
        RECT -38.450 8.560 -36.510 8.710 ;
        RECT -41.790 7.770 -41.470 7.880 ;
        RECT -42.290 7.630 -41.470 7.770 ;
        RECT -41.790 7.600 -41.470 7.630 ;
        RECT -39.110 7.770 -38.790 7.880 ;
        RECT -38.450 7.770 -38.290 8.560 ;
        RECT -36.850 8.410 -36.510 8.560 ;
        RECT -34.150 8.560 -32.210 8.710 ;
        RECT -34.150 8.410 -33.810 8.560 ;
        RECT -36.830 8.210 -36.510 8.240 ;
        RECT -39.110 7.630 -38.290 7.770 ;
        RECT -37.330 8.070 -36.510 8.210 ;
        RECT -39.110 7.600 -38.790 7.630 ;
        RECT -41.810 7.280 -41.470 7.430 ;
        RECT -43.410 7.130 -41.470 7.280 ;
        RECT -39.110 7.280 -38.770 7.430 ;
        RECT -37.330 7.280 -37.170 8.070 ;
        RECT -36.830 7.960 -36.510 8.070 ;
        RECT -34.150 8.210 -33.830 8.240 ;
        RECT -34.150 8.070 -33.330 8.210 ;
        RECT -34.150 7.960 -33.830 8.070 ;
        RECT -39.110 7.130 -37.170 7.280 ;
        RECT -33.490 7.280 -33.330 8.070 ;
        RECT -32.370 7.770 -32.210 8.560 ;
        RECT -28.530 8.560 -26.590 8.710 ;
        RECT -31.870 7.770 -31.550 7.880 ;
        RECT -32.370 7.630 -31.550 7.770 ;
        RECT -31.870 7.600 -31.550 7.630 ;
        RECT -29.190 7.770 -28.870 7.880 ;
        RECT -28.530 7.770 -28.370 8.560 ;
        RECT -26.930 8.410 -26.590 8.560 ;
        RECT -24.230 8.560 -22.290 8.710 ;
        RECT -24.230 8.410 -23.890 8.560 ;
        RECT -26.910 8.210 -26.590 8.240 ;
        RECT -29.190 7.630 -28.370 7.770 ;
        RECT -27.410 8.070 -26.590 8.210 ;
        RECT -29.190 7.600 -28.870 7.630 ;
        RECT -31.890 7.280 -31.550 7.430 ;
        RECT -33.490 7.130 -31.550 7.280 ;
        RECT -29.190 7.280 -28.850 7.430 ;
        RECT -27.410 7.280 -27.250 8.070 ;
        RECT -26.910 7.960 -26.590 8.070 ;
        RECT -24.230 8.210 -23.910 8.240 ;
        RECT -24.230 8.070 -23.410 8.210 ;
        RECT -24.230 7.960 -23.910 8.070 ;
        RECT -29.190 7.130 -27.250 7.280 ;
        RECT -23.570 7.280 -23.410 8.070 ;
        RECT -22.450 7.770 -22.290 8.560 ;
        RECT -18.610 8.560 -16.670 8.710 ;
        RECT -21.950 7.770 -21.630 7.880 ;
        RECT -22.450 7.630 -21.630 7.770 ;
        RECT -21.950 7.600 -21.630 7.630 ;
        RECT -19.270 7.770 -18.950 7.880 ;
        RECT -18.610 7.770 -18.450 8.560 ;
        RECT -17.010 8.410 -16.670 8.560 ;
        RECT -14.310 8.560 -12.370 8.710 ;
        RECT -14.310 8.410 -13.970 8.560 ;
        RECT -16.990 8.210 -16.670 8.240 ;
        RECT -19.270 7.630 -18.450 7.770 ;
        RECT -17.490 8.070 -16.670 8.210 ;
        RECT -19.270 7.600 -18.950 7.630 ;
        RECT -21.970 7.280 -21.630 7.430 ;
        RECT -23.570 7.130 -21.630 7.280 ;
        RECT -19.270 7.280 -18.930 7.430 ;
        RECT -17.490 7.280 -17.330 8.070 ;
        RECT -16.990 7.960 -16.670 8.070 ;
        RECT -14.310 8.210 -13.990 8.240 ;
        RECT -14.310 8.070 -13.490 8.210 ;
        RECT -14.310 7.960 -13.990 8.070 ;
        RECT -19.270 7.130 -17.330 7.280 ;
        RECT -13.650 7.280 -13.490 8.070 ;
        RECT -12.530 7.770 -12.370 8.560 ;
        RECT -8.690 8.560 -6.750 8.710 ;
        RECT -12.030 7.770 -11.710 7.880 ;
        RECT -12.530 7.630 -11.710 7.770 ;
        RECT -12.030 7.600 -11.710 7.630 ;
        RECT -9.350 7.770 -9.030 7.880 ;
        RECT -8.690 7.770 -8.530 8.560 ;
        RECT -7.090 8.410 -6.750 8.560 ;
        RECT -4.390 8.560 -2.450 8.710 ;
        RECT -4.390 8.410 -4.050 8.560 ;
        RECT -7.070 8.210 -6.750 8.240 ;
        RECT -9.350 7.630 -8.530 7.770 ;
        RECT -7.570 8.070 -6.750 8.210 ;
        RECT -9.350 7.600 -9.030 7.630 ;
        RECT -12.050 7.280 -11.710 7.430 ;
        RECT -13.650 7.130 -11.710 7.280 ;
        RECT -9.350 7.280 -9.010 7.430 ;
        RECT -7.570 7.280 -7.410 8.070 ;
        RECT -7.070 7.960 -6.750 8.070 ;
        RECT -4.390 8.210 -4.070 8.240 ;
        RECT -4.390 8.070 -3.570 8.210 ;
        RECT -4.390 7.960 -4.070 8.070 ;
        RECT -9.350 7.130 -7.410 7.280 ;
        RECT -3.730 7.280 -3.570 8.070 ;
        RECT -2.610 7.770 -2.450 8.560 ;
        RECT 1.230 8.560 3.170 8.710 ;
        RECT -2.110 7.770 -1.790 7.880 ;
        RECT -2.610 7.630 -1.790 7.770 ;
        RECT -2.110 7.600 -1.790 7.630 ;
        RECT 0.570 7.770 0.890 7.880 ;
        RECT 1.230 7.770 1.390 8.560 ;
        RECT 2.830 8.410 3.170 8.560 ;
        RECT 5.530 8.560 7.470 8.710 ;
        RECT 5.530 8.410 5.870 8.560 ;
        RECT 2.850 8.210 3.170 8.240 ;
        RECT 0.570 7.630 1.390 7.770 ;
        RECT 2.350 8.070 3.170 8.210 ;
        RECT 0.570 7.600 0.890 7.630 ;
        RECT -2.130 7.280 -1.790 7.430 ;
        RECT -3.730 7.130 -1.790 7.280 ;
        RECT 0.570 7.280 0.910 7.430 ;
        RECT 2.350 7.280 2.510 8.070 ;
        RECT 2.850 7.960 3.170 8.070 ;
        RECT 5.530 8.210 5.850 8.240 ;
        RECT 5.530 8.070 6.350 8.210 ;
        RECT 5.530 7.960 5.850 8.070 ;
        RECT 0.570 7.130 2.510 7.280 ;
        RECT 6.190 7.280 6.350 8.070 ;
        RECT 7.310 7.770 7.470 8.560 ;
        RECT 11.150 8.560 13.090 8.710 ;
        RECT 7.810 7.770 8.130 7.880 ;
        RECT 7.310 7.630 8.130 7.770 ;
        RECT 7.810 7.600 8.130 7.630 ;
        RECT 10.490 7.770 10.810 7.880 ;
        RECT 11.150 7.770 11.310 8.560 ;
        RECT 12.750 8.410 13.090 8.560 ;
        RECT 15.450 8.560 17.390 8.710 ;
        RECT 15.450 8.410 15.790 8.560 ;
        RECT 12.770 8.210 13.090 8.240 ;
        RECT 10.490 7.630 11.310 7.770 ;
        RECT 12.270 8.070 13.090 8.210 ;
        RECT 10.490 7.600 10.810 7.630 ;
        RECT 7.790 7.280 8.130 7.430 ;
        RECT 6.190 7.130 8.130 7.280 ;
        RECT 10.490 7.280 10.830 7.430 ;
        RECT 12.270 7.280 12.430 8.070 ;
        RECT 12.770 7.960 13.090 8.070 ;
        RECT 15.450 8.210 15.770 8.240 ;
        RECT 15.450 8.070 16.270 8.210 ;
        RECT 15.450 7.960 15.770 8.070 ;
        RECT 10.490 7.130 12.430 7.280 ;
        RECT 16.110 7.280 16.270 8.070 ;
        RECT 17.230 7.770 17.390 8.560 ;
        RECT 21.070 8.560 23.010 8.710 ;
        RECT 17.730 7.770 18.050 7.880 ;
        RECT 17.230 7.630 18.050 7.770 ;
        RECT 17.730 7.600 18.050 7.630 ;
        RECT 20.410 7.770 20.730 7.880 ;
        RECT 21.070 7.770 21.230 8.560 ;
        RECT 22.670 8.410 23.010 8.560 ;
        RECT 22.690 8.210 23.010 8.240 ;
        RECT 20.410 7.630 21.230 7.770 ;
        RECT 22.190 8.070 23.010 8.210 ;
        RECT 20.410 7.600 20.730 7.630 ;
        RECT 17.710 7.280 18.050 7.430 ;
        RECT 16.110 7.130 18.050 7.280 ;
        RECT 20.410 7.280 20.750 7.430 ;
        RECT 22.190 7.280 22.350 8.070 ;
        RECT 22.690 7.960 23.010 8.070 ;
        RECT 20.410 7.130 22.350 7.280 ;
        RECT -293.480 6.320 -291.640 6.800 ;
        RECT -291.720 5.230 -291.240 6.130 ;
        RECT -290.420 6.000 -290.230 7.130 ;
        RECT -286.350 6.000 -286.160 7.130 ;
        RECT -280.500 6.000 -280.310 7.130 ;
        RECT -276.430 6.000 -276.240 7.130 ;
        RECT -270.580 6.000 -270.390 7.130 ;
        RECT -266.510 6.000 -266.320 7.130 ;
        RECT -260.660 6.000 -260.470 7.130 ;
        RECT -256.590 6.000 -256.400 7.130 ;
        RECT -250.740 6.000 -250.550 7.130 ;
        RECT -246.670 6.000 -246.480 7.130 ;
        RECT -240.820 6.000 -240.630 7.130 ;
        RECT -236.750 6.000 -236.560 7.130 ;
        RECT -230.900 6.000 -230.710 7.130 ;
        RECT -226.830 6.000 -226.640 7.130 ;
        RECT -220.980 6.000 -220.790 7.130 ;
        RECT -216.910 6.000 -216.720 7.130 ;
        RECT -211.060 6.000 -210.870 7.130 ;
        RECT -206.990 6.000 -206.800 7.130 ;
        RECT -201.140 6.000 -200.950 7.130 ;
        RECT -197.070 6.000 -196.880 7.130 ;
        RECT -191.220 6.000 -191.030 7.130 ;
        RECT -187.150 6.000 -186.960 7.130 ;
        RECT -181.300 6.000 -181.110 7.130 ;
        RECT -177.230 6.000 -177.040 7.130 ;
        RECT -171.380 6.000 -171.190 7.130 ;
        RECT -167.310 6.000 -167.120 7.130 ;
        RECT -161.460 6.000 -161.270 7.130 ;
        RECT -157.390 6.000 -157.200 7.130 ;
        RECT -151.540 6.000 -151.350 7.130 ;
        RECT -147.470 6.000 -147.280 7.130 ;
        RECT -141.620 6.000 -141.430 7.130 ;
        RECT -137.550 6.000 -137.360 7.130 ;
        RECT -131.700 6.000 -131.510 7.130 ;
        RECT -127.630 6.000 -127.440 7.130 ;
        RECT -121.780 6.000 -121.590 7.130 ;
        RECT -117.710 6.000 -117.520 7.130 ;
        RECT -111.860 6.000 -111.670 7.130 ;
        RECT -107.790 6.000 -107.600 7.130 ;
        RECT -101.940 6.000 -101.750 7.130 ;
        RECT -97.870 6.000 -97.680 7.130 ;
        RECT -92.020 6.000 -91.830 7.130 ;
        RECT -87.950 6.000 -87.760 7.130 ;
        RECT -82.100 6.000 -81.910 7.130 ;
        RECT -78.030 6.000 -77.840 7.130 ;
        RECT -72.180 6.000 -71.990 7.130 ;
        RECT -68.110 6.000 -67.920 7.130 ;
        RECT -62.260 6.000 -62.070 7.130 ;
        RECT -58.190 6.000 -58.000 7.130 ;
        RECT -52.340 6.000 -52.150 7.130 ;
        RECT -48.270 6.000 -48.080 7.130 ;
        RECT -42.420 6.000 -42.230 7.130 ;
        RECT -38.350 6.000 -38.160 7.130 ;
        RECT -32.500 6.000 -32.310 7.130 ;
        RECT -28.430 6.000 -28.240 7.130 ;
        RECT -22.580 6.000 -22.390 7.130 ;
        RECT -18.510 6.000 -18.320 7.130 ;
        RECT -12.660 6.000 -12.470 7.130 ;
        RECT -8.590 6.000 -8.400 7.130 ;
        RECT -2.740 6.000 -2.550 7.130 ;
        RECT 1.330 6.000 1.520 7.130 ;
        RECT 7.180 6.000 7.370 7.130 ;
        RECT 11.250 6.000 11.440 7.130 ;
        RECT 17.100 6.000 17.290 7.130 ;
        RECT 21.170 6.000 21.360 7.130 ;
        RECT -290.470 5.710 -290.150 6.000 ;
        RECT -286.430 5.710 -286.110 6.000 ;
        RECT -280.550 5.710 -280.230 6.000 ;
        RECT -276.510 5.710 -276.190 6.000 ;
        RECT -270.630 5.710 -270.310 6.000 ;
        RECT -266.590 5.710 -266.270 6.000 ;
        RECT -260.710 5.710 -260.390 6.000 ;
        RECT -256.670 5.710 -256.350 6.000 ;
        RECT -250.790 5.710 -250.470 6.000 ;
        RECT -246.750 5.710 -246.430 6.000 ;
        RECT -240.870 5.710 -240.550 6.000 ;
        RECT -236.830 5.710 -236.510 6.000 ;
        RECT -230.950 5.710 -230.630 6.000 ;
        RECT -226.910 5.710 -226.590 6.000 ;
        RECT -221.030 5.710 -220.710 6.000 ;
        RECT -216.990 5.710 -216.670 6.000 ;
        RECT -211.110 5.710 -210.790 6.000 ;
        RECT -207.070 5.710 -206.750 6.000 ;
        RECT -201.190 5.710 -200.870 6.000 ;
        RECT -197.150 5.710 -196.830 6.000 ;
        RECT -191.270 5.710 -190.950 6.000 ;
        RECT -187.230 5.710 -186.910 6.000 ;
        RECT -181.350 5.710 -181.030 6.000 ;
        RECT -177.310 5.710 -176.990 6.000 ;
        RECT -171.430 5.710 -171.110 6.000 ;
        RECT -167.390 5.710 -167.070 6.000 ;
        RECT -161.510 5.710 -161.190 6.000 ;
        RECT -157.470 5.710 -157.150 6.000 ;
        RECT -151.590 5.710 -151.270 6.000 ;
        RECT -147.550 5.710 -147.230 6.000 ;
        RECT -141.670 5.710 -141.350 6.000 ;
        RECT -137.630 5.710 -137.310 6.000 ;
        RECT -131.750 5.710 -131.430 6.000 ;
        RECT -127.710 5.710 -127.390 6.000 ;
        RECT -121.830 5.710 -121.510 6.000 ;
        RECT -117.790 5.710 -117.470 6.000 ;
        RECT -111.910 5.710 -111.590 6.000 ;
        RECT -107.870 5.710 -107.550 6.000 ;
        RECT -101.990 5.710 -101.670 6.000 ;
        RECT -97.950 5.710 -97.630 6.000 ;
        RECT -92.070 5.710 -91.750 6.000 ;
        RECT -88.030 5.710 -87.710 6.000 ;
        RECT -82.150 5.710 -81.830 6.000 ;
        RECT -78.110 5.710 -77.790 6.000 ;
        RECT -72.230 5.710 -71.910 6.000 ;
        RECT -68.190 5.710 -67.870 6.000 ;
        RECT -62.310 5.710 -61.990 6.000 ;
        RECT -58.270 5.710 -57.950 6.000 ;
        RECT -52.390 5.710 -52.070 6.000 ;
        RECT -48.350 5.710 -48.030 6.000 ;
        RECT -42.470 5.710 -42.150 6.000 ;
        RECT -38.430 5.710 -38.110 6.000 ;
        RECT -32.550 5.710 -32.230 6.000 ;
        RECT -28.510 5.710 -28.190 6.000 ;
        RECT -22.630 5.710 -22.310 6.000 ;
        RECT -18.590 5.710 -18.270 6.000 ;
        RECT -12.710 5.710 -12.390 6.000 ;
        RECT -8.670 5.710 -8.350 6.000 ;
        RECT -2.790 5.710 -2.470 6.000 ;
        RECT 1.250 5.710 1.570 6.000 ;
        RECT 7.130 5.710 7.450 6.000 ;
        RECT 11.170 5.710 11.490 6.000 ;
        RECT 17.050 5.710 17.370 6.000 ;
        RECT 21.090 5.710 21.410 6.000 ;
        RECT -292.180 4.750 -291.240 5.230 ;
        RECT 22.180 5.230 22.660 6.130 ;
        RECT -287.170 4.830 -285.480 5.130 ;
        RECT -277.250 4.830 -275.560 5.130 ;
        RECT -267.330 4.830 -265.640 5.130 ;
        RECT -257.410 4.830 -255.720 5.130 ;
        RECT -247.490 4.830 -245.800 5.130 ;
        RECT -237.570 4.830 -235.880 5.130 ;
        RECT -227.650 4.830 -225.960 5.130 ;
        RECT -217.730 4.830 -216.040 5.130 ;
        RECT -207.810 4.830 -206.120 5.130 ;
        RECT -197.890 4.830 -196.200 5.130 ;
        RECT -187.970 4.830 -186.280 5.130 ;
        RECT -178.050 4.830 -176.360 5.130 ;
        RECT -168.130 4.830 -166.440 5.130 ;
        RECT -158.210 4.830 -156.520 5.130 ;
        RECT -148.290 4.830 -146.600 5.130 ;
        RECT -138.370 4.830 -136.680 5.130 ;
        RECT -128.450 4.830 -126.760 5.130 ;
        RECT -118.530 4.830 -116.840 5.130 ;
        RECT -108.610 4.830 -106.920 5.130 ;
        RECT -98.690 4.830 -97.000 5.130 ;
        RECT -88.770 4.830 -87.080 5.130 ;
        RECT -78.850 4.830 -77.160 5.130 ;
        RECT -68.930 4.830 -67.240 5.130 ;
        RECT -59.010 4.830 -57.320 5.130 ;
        RECT -49.090 4.830 -47.400 5.130 ;
        RECT -39.170 4.830 -37.480 5.130 ;
        RECT -29.250 4.830 -27.560 5.130 ;
        RECT -19.330 4.830 -17.640 5.130 ;
        RECT -9.410 4.830 -7.720 5.130 ;
        RECT 0.510 4.830 2.200 5.130 ;
        RECT 10.430 4.830 12.120 5.130 ;
        RECT 20.350 4.830 22.040 5.130 ;
        RECT -286.660 4.130 -285.660 4.830 ;
        RECT -276.740 4.130 -275.740 4.830 ;
        RECT -266.820 4.130 -265.820 4.830 ;
        RECT -256.900 4.130 -255.900 4.830 ;
        RECT -246.980 4.130 -245.980 4.830 ;
        RECT -237.060 4.130 -236.060 4.830 ;
        RECT -227.140 4.130 -226.140 4.830 ;
        RECT -217.220 4.130 -216.220 4.830 ;
        RECT -207.300 4.130 -206.300 4.830 ;
        RECT -197.380 4.130 -196.380 4.830 ;
        RECT -187.460 4.130 -186.460 4.830 ;
        RECT -177.540 4.130 -176.540 4.830 ;
        RECT -167.620 4.130 -166.620 4.830 ;
        RECT -157.700 4.130 -156.700 4.830 ;
        RECT -147.780 4.130 -146.780 4.830 ;
        RECT -137.860 4.130 -136.860 4.830 ;
        RECT -127.940 4.130 -126.940 4.830 ;
        RECT -118.020 4.130 -117.020 4.830 ;
        RECT -108.100 4.130 -107.100 4.830 ;
        RECT -98.180 4.130 -97.180 4.830 ;
        RECT -88.260 4.130 -87.260 4.830 ;
        RECT -78.340 4.130 -77.340 4.830 ;
        RECT -68.420 4.130 -67.420 4.830 ;
        RECT -58.500 4.130 -57.500 4.830 ;
        RECT -48.580 4.130 -47.580 4.830 ;
        RECT -38.660 4.130 -37.660 4.830 ;
        RECT -28.740 4.130 -27.740 4.830 ;
        RECT -18.820 4.130 -17.820 4.830 ;
        RECT -8.900 4.130 -7.900 4.830 ;
        RECT 1.020 4.130 2.020 4.830 ;
        RECT 10.940 4.130 11.940 4.830 ;
        RECT 20.860 4.130 21.860 4.830 ;
        RECT 22.180 4.750 23.120 5.230 ;
        RECT -293.120 -77.860 -292.660 -77.855 ;
        RECT -293.120 -78.335 -292.180 -77.860 ;
        RECT -291.260 -77.940 -290.260 -77.240 ;
        RECT -281.340 -77.940 -280.340 -77.240 ;
        RECT -271.420 -77.940 -270.420 -77.240 ;
        RECT -261.500 -77.940 -260.500 -77.240 ;
        RECT -251.580 -77.940 -250.580 -77.240 ;
        RECT -241.660 -77.940 -240.660 -77.240 ;
        RECT -231.740 -77.940 -230.740 -77.240 ;
        RECT -221.820 -77.940 -220.820 -77.240 ;
        RECT -211.900 -77.940 -210.900 -77.240 ;
        RECT -201.980 -77.940 -200.980 -77.240 ;
        RECT -192.060 -77.940 -191.060 -77.240 ;
        RECT -182.140 -77.940 -181.140 -77.240 ;
        RECT -172.220 -77.940 -171.220 -77.240 ;
        RECT -162.300 -77.940 -161.300 -77.240 ;
        RECT -152.380 -77.940 -151.380 -77.240 ;
        RECT -142.460 -77.940 -141.460 -77.240 ;
        RECT -132.540 -77.940 -131.540 -77.240 ;
        RECT -122.620 -77.940 -121.620 -77.240 ;
        RECT -112.700 -77.940 -111.700 -77.240 ;
        RECT -102.780 -77.940 -101.780 -77.240 ;
        RECT -92.860 -77.940 -91.860 -77.240 ;
        RECT -82.940 -77.940 -81.940 -77.240 ;
        RECT -73.020 -77.940 -72.020 -77.240 ;
        RECT -63.100 -77.940 -62.100 -77.240 ;
        RECT -53.180 -77.940 -52.180 -77.240 ;
        RECT -43.260 -77.940 -42.260 -77.240 ;
        RECT -33.340 -77.940 -32.340 -77.240 ;
        RECT -23.420 -77.940 -22.420 -77.240 ;
        RECT -13.500 -77.940 -12.500 -77.240 ;
        RECT -3.580 -77.940 -2.580 -77.240 ;
        RECT 6.340 -77.940 7.340 -77.240 ;
        RECT 16.260 -77.940 17.260 -77.240 ;
        RECT -291.770 -78.240 -290.080 -77.940 ;
        RECT -281.850 -78.240 -280.160 -77.940 ;
        RECT -271.930 -78.240 -270.240 -77.940 ;
        RECT -262.010 -78.240 -260.320 -77.940 ;
        RECT -252.090 -78.240 -250.400 -77.940 ;
        RECT -242.170 -78.240 -240.480 -77.940 ;
        RECT -232.250 -78.240 -230.560 -77.940 ;
        RECT -222.330 -78.240 -220.640 -77.940 ;
        RECT -212.410 -78.240 -210.720 -77.940 ;
        RECT -202.490 -78.240 -200.800 -77.940 ;
        RECT -192.570 -78.240 -190.880 -77.940 ;
        RECT -182.650 -78.240 -180.960 -77.940 ;
        RECT -172.730 -78.240 -171.040 -77.940 ;
        RECT -162.810 -78.240 -161.120 -77.940 ;
        RECT -152.890 -78.240 -151.200 -77.940 ;
        RECT -142.970 -78.240 -141.280 -77.940 ;
        RECT -133.050 -78.240 -131.360 -77.940 ;
        RECT -123.130 -78.240 -121.440 -77.940 ;
        RECT -113.210 -78.240 -111.520 -77.940 ;
        RECT -103.290 -78.240 -101.600 -77.940 ;
        RECT -93.370 -78.240 -91.680 -77.940 ;
        RECT -83.450 -78.240 -81.760 -77.940 ;
        RECT -73.530 -78.240 -71.840 -77.940 ;
        RECT -63.610 -78.240 -61.920 -77.940 ;
        RECT -53.690 -78.240 -52.000 -77.940 ;
        RECT -43.770 -78.240 -42.080 -77.940 ;
        RECT -33.850 -78.240 -32.160 -77.940 ;
        RECT -23.930 -78.240 -22.240 -77.940 ;
        RECT -14.010 -78.240 -12.320 -77.940 ;
        RECT -4.090 -78.240 -2.400 -77.940 ;
        RECT 5.830 -78.240 7.520 -77.940 ;
        RECT 15.750 -78.240 17.440 -77.940 ;
        RECT -292.660 -79.240 -292.180 -78.335 ;
        RECT -291.030 -79.110 -290.710 -78.820 ;
        RECT -285.150 -79.110 -284.830 -78.820 ;
        RECT -281.110 -79.110 -280.790 -78.820 ;
        RECT -275.230 -79.110 -274.910 -78.820 ;
        RECT -271.190 -79.110 -270.870 -78.820 ;
        RECT -265.310 -79.110 -264.990 -78.820 ;
        RECT -261.270 -79.110 -260.950 -78.820 ;
        RECT -255.390 -79.110 -255.070 -78.820 ;
        RECT -251.350 -79.110 -251.030 -78.820 ;
        RECT -245.470 -79.110 -245.150 -78.820 ;
        RECT -241.430 -79.110 -241.110 -78.820 ;
        RECT -235.550 -79.110 -235.230 -78.820 ;
        RECT -231.510 -79.110 -231.190 -78.820 ;
        RECT -225.630 -79.110 -225.310 -78.820 ;
        RECT -221.590 -79.110 -221.270 -78.820 ;
        RECT -215.710 -79.110 -215.390 -78.820 ;
        RECT -211.670 -79.110 -211.350 -78.820 ;
        RECT -205.790 -79.110 -205.470 -78.820 ;
        RECT -201.750 -79.110 -201.430 -78.820 ;
        RECT -195.870 -79.110 -195.550 -78.820 ;
        RECT -191.830 -79.110 -191.510 -78.820 ;
        RECT -185.950 -79.110 -185.630 -78.820 ;
        RECT -181.910 -79.110 -181.590 -78.820 ;
        RECT -176.030 -79.110 -175.710 -78.820 ;
        RECT -171.990 -79.110 -171.670 -78.820 ;
        RECT -166.110 -79.110 -165.790 -78.820 ;
        RECT -162.070 -79.110 -161.750 -78.820 ;
        RECT -156.190 -79.110 -155.870 -78.820 ;
        RECT -152.150 -79.110 -151.830 -78.820 ;
        RECT -146.270 -79.110 -145.950 -78.820 ;
        RECT -142.230 -79.110 -141.910 -78.820 ;
        RECT -136.350 -79.110 -136.030 -78.820 ;
        RECT -132.310 -79.110 -131.990 -78.820 ;
        RECT -126.430 -79.110 -126.110 -78.820 ;
        RECT -122.390 -79.110 -122.070 -78.820 ;
        RECT -116.510 -79.110 -116.190 -78.820 ;
        RECT -112.470 -79.110 -112.150 -78.820 ;
        RECT -106.590 -79.110 -106.270 -78.820 ;
        RECT -102.550 -79.110 -102.230 -78.820 ;
        RECT -96.670 -79.110 -96.350 -78.820 ;
        RECT -92.630 -79.110 -92.310 -78.820 ;
        RECT -86.750 -79.110 -86.430 -78.820 ;
        RECT -82.710 -79.110 -82.390 -78.820 ;
        RECT -76.830 -79.110 -76.510 -78.820 ;
        RECT -72.790 -79.110 -72.470 -78.820 ;
        RECT -66.910 -79.110 -66.590 -78.820 ;
        RECT -62.870 -79.110 -62.550 -78.820 ;
        RECT -56.990 -79.110 -56.670 -78.820 ;
        RECT -52.950 -79.110 -52.630 -78.820 ;
        RECT -47.070 -79.110 -46.750 -78.820 ;
        RECT -43.030 -79.110 -42.710 -78.820 ;
        RECT -37.150 -79.110 -36.830 -78.820 ;
        RECT -33.110 -79.110 -32.790 -78.820 ;
        RECT -27.230 -79.110 -26.910 -78.820 ;
        RECT -23.190 -79.110 -22.870 -78.820 ;
        RECT -17.310 -79.110 -16.990 -78.820 ;
        RECT -13.270 -79.110 -12.950 -78.820 ;
        RECT -7.390 -79.110 -7.070 -78.820 ;
        RECT -3.350 -79.110 -3.030 -78.820 ;
        RECT 2.530 -79.110 2.850 -78.820 ;
        RECT 6.570 -79.110 6.890 -78.820 ;
        RECT 12.450 -79.110 12.770 -78.820 ;
        RECT 16.490 -79.110 16.810 -78.820 ;
        RECT 22.370 -79.110 22.690 -78.820 ;
        RECT -293.120 -79.910 -291.280 -79.430 ;
        RECT -290.950 -80.240 -290.760 -79.110 ;
        RECT -285.100 -80.240 -284.910 -79.110 ;
        RECT -281.030 -80.240 -280.840 -79.110 ;
        RECT -275.180 -80.240 -274.990 -79.110 ;
        RECT -271.110 -80.240 -270.920 -79.110 ;
        RECT -265.260 -80.240 -265.070 -79.110 ;
        RECT -261.190 -80.240 -261.000 -79.110 ;
        RECT -255.340 -80.240 -255.150 -79.110 ;
        RECT -251.270 -80.240 -251.080 -79.110 ;
        RECT -245.420 -80.240 -245.230 -79.110 ;
        RECT -241.350 -80.240 -241.160 -79.110 ;
        RECT -235.500 -80.240 -235.310 -79.110 ;
        RECT -231.430 -80.240 -231.240 -79.110 ;
        RECT -225.580 -80.240 -225.390 -79.110 ;
        RECT -221.510 -80.240 -221.320 -79.110 ;
        RECT -215.660 -80.240 -215.470 -79.110 ;
        RECT -211.590 -80.240 -211.400 -79.110 ;
        RECT -205.740 -80.240 -205.550 -79.110 ;
        RECT -201.670 -80.240 -201.480 -79.110 ;
        RECT -195.820 -80.240 -195.630 -79.110 ;
        RECT -191.750 -80.240 -191.560 -79.110 ;
        RECT -185.900 -80.240 -185.710 -79.110 ;
        RECT -181.830 -80.240 -181.640 -79.110 ;
        RECT -175.980 -80.240 -175.790 -79.110 ;
        RECT -171.910 -80.240 -171.720 -79.110 ;
        RECT -166.060 -80.240 -165.870 -79.110 ;
        RECT -161.990 -80.240 -161.800 -79.110 ;
        RECT -156.140 -80.240 -155.950 -79.110 ;
        RECT -152.070 -80.240 -151.880 -79.110 ;
        RECT -146.220 -80.240 -146.030 -79.110 ;
        RECT -142.150 -80.240 -141.960 -79.110 ;
        RECT -136.300 -80.240 -136.110 -79.110 ;
        RECT -132.230 -80.240 -132.040 -79.110 ;
        RECT -126.380 -80.240 -126.190 -79.110 ;
        RECT -122.310 -80.240 -122.120 -79.110 ;
        RECT -116.460 -80.240 -116.270 -79.110 ;
        RECT -112.390 -80.240 -112.200 -79.110 ;
        RECT -106.540 -80.240 -106.350 -79.110 ;
        RECT -102.470 -80.240 -102.280 -79.110 ;
        RECT -96.620 -80.240 -96.430 -79.110 ;
        RECT -92.550 -80.240 -92.360 -79.110 ;
        RECT -86.700 -80.240 -86.510 -79.110 ;
        RECT -82.630 -80.240 -82.440 -79.110 ;
        RECT -76.780 -80.240 -76.590 -79.110 ;
        RECT -72.710 -80.240 -72.520 -79.110 ;
        RECT -66.860 -80.240 -66.670 -79.110 ;
        RECT -62.790 -80.240 -62.600 -79.110 ;
        RECT -56.940 -80.240 -56.750 -79.110 ;
        RECT -52.870 -80.240 -52.680 -79.110 ;
        RECT -47.020 -80.240 -46.830 -79.110 ;
        RECT -42.950 -80.240 -42.760 -79.110 ;
        RECT -37.100 -80.240 -36.910 -79.110 ;
        RECT -33.030 -80.240 -32.840 -79.110 ;
        RECT -27.180 -80.240 -26.990 -79.110 ;
        RECT -23.110 -80.240 -22.920 -79.110 ;
        RECT -17.260 -80.240 -17.070 -79.110 ;
        RECT -13.190 -80.240 -13.000 -79.110 ;
        RECT -7.340 -80.240 -7.150 -79.110 ;
        RECT -3.270 -80.240 -3.080 -79.110 ;
        RECT 2.580 -80.240 2.770 -79.110 ;
        RECT 6.650 -80.240 6.840 -79.110 ;
        RECT 12.500 -80.240 12.690 -79.110 ;
        RECT 16.570 -80.240 16.760 -79.110 ;
        RECT 22.420 -80.240 22.610 -79.110 ;
        RECT 22.940 -79.910 24.780 -79.430 ;
        RECT -291.710 -80.390 -289.770 -80.240 ;
        RECT -291.710 -80.540 -291.370 -80.390 ;
        RECT -291.710 -80.740 -291.390 -80.710 ;
        RECT -291.710 -80.880 -290.890 -80.740 ;
        RECT -291.710 -80.990 -291.390 -80.880 ;
        RECT -291.050 -81.670 -290.890 -80.880 ;
        RECT -289.930 -81.180 -289.770 -80.390 ;
        RECT -286.090 -80.390 -284.150 -80.240 ;
        RECT -289.430 -81.180 -289.110 -81.070 ;
        RECT -289.930 -81.320 -289.110 -81.180 ;
        RECT -289.430 -81.350 -289.110 -81.320 ;
        RECT -286.750 -81.180 -286.430 -81.070 ;
        RECT -286.090 -81.180 -285.930 -80.390 ;
        RECT -284.490 -80.540 -284.150 -80.390 ;
        RECT -281.790 -80.390 -279.850 -80.240 ;
        RECT -281.790 -80.540 -281.450 -80.390 ;
        RECT -284.470 -80.740 -284.150 -80.710 ;
        RECT -286.750 -81.320 -285.930 -81.180 ;
        RECT -284.970 -80.880 -284.150 -80.740 ;
        RECT -286.750 -81.350 -286.430 -81.320 ;
        RECT -289.450 -81.670 -289.110 -81.520 ;
        RECT -291.050 -81.820 -289.110 -81.670 ;
        RECT -286.750 -81.670 -286.410 -81.520 ;
        RECT -284.970 -81.670 -284.810 -80.880 ;
        RECT -284.470 -80.990 -284.150 -80.880 ;
        RECT -281.790 -80.740 -281.470 -80.710 ;
        RECT -281.790 -80.880 -280.970 -80.740 ;
        RECT -281.790 -80.990 -281.470 -80.880 ;
        RECT -286.750 -81.820 -284.810 -81.670 ;
        RECT -281.130 -81.670 -280.970 -80.880 ;
        RECT -280.010 -81.180 -279.850 -80.390 ;
        RECT -276.170 -80.390 -274.230 -80.240 ;
        RECT -279.510 -81.180 -279.190 -81.070 ;
        RECT -280.010 -81.320 -279.190 -81.180 ;
        RECT -279.510 -81.350 -279.190 -81.320 ;
        RECT -276.830 -81.180 -276.510 -81.070 ;
        RECT -276.170 -81.180 -276.010 -80.390 ;
        RECT -274.570 -80.540 -274.230 -80.390 ;
        RECT -271.870 -80.390 -269.930 -80.240 ;
        RECT -271.870 -80.540 -271.530 -80.390 ;
        RECT -274.550 -80.740 -274.230 -80.710 ;
        RECT -276.830 -81.320 -276.010 -81.180 ;
        RECT -275.050 -80.880 -274.230 -80.740 ;
        RECT -276.830 -81.350 -276.510 -81.320 ;
        RECT -279.530 -81.670 -279.190 -81.520 ;
        RECT -281.130 -81.820 -279.190 -81.670 ;
        RECT -276.830 -81.670 -276.490 -81.520 ;
        RECT -275.050 -81.670 -274.890 -80.880 ;
        RECT -274.550 -80.990 -274.230 -80.880 ;
        RECT -271.870 -80.740 -271.550 -80.710 ;
        RECT -271.870 -80.880 -271.050 -80.740 ;
        RECT -271.870 -80.990 -271.550 -80.880 ;
        RECT -276.830 -81.820 -274.890 -81.670 ;
        RECT -271.210 -81.670 -271.050 -80.880 ;
        RECT -270.090 -81.180 -269.930 -80.390 ;
        RECT -266.250 -80.390 -264.310 -80.240 ;
        RECT -269.590 -81.180 -269.270 -81.070 ;
        RECT -270.090 -81.320 -269.270 -81.180 ;
        RECT -269.590 -81.350 -269.270 -81.320 ;
        RECT -266.910 -81.180 -266.590 -81.070 ;
        RECT -266.250 -81.180 -266.090 -80.390 ;
        RECT -264.650 -80.540 -264.310 -80.390 ;
        RECT -261.950 -80.390 -260.010 -80.240 ;
        RECT -261.950 -80.540 -261.610 -80.390 ;
        RECT -264.630 -80.740 -264.310 -80.710 ;
        RECT -266.910 -81.320 -266.090 -81.180 ;
        RECT -265.130 -80.880 -264.310 -80.740 ;
        RECT -266.910 -81.350 -266.590 -81.320 ;
        RECT -269.610 -81.670 -269.270 -81.520 ;
        RECT -271.210 -81.820 -269.270 -81.670 ;
        RECT -266.910 -81.670 -266.570 -81.520 ;
        RECT -265.130 -81.670 -264.970 -80.880 ;
        RECT -264.630 -80.990 -264.310 -80.880 ;
        RECT -261.950 -80.740 -261.630 -80.710 ;
        RECT -261.950 -80.880 -261.130 -80.740 ;
        RECT -261.950 -80.990 -261.630 -80.880 ;
        RECT -266.910 -81.820 -264.970 -81.670 ;
        RECT -261.290 -81.670 -261.130 -80.880 ;
        RECT -260.170 -81.180 -260.010 -80.390 ;
        RECT -256.330 -80.390 -254.390 -80.240 ;
        RECT -259.670 -81.180 -259.350 -81.070 ;
        RECT -260.170 -81.320 -259.350 -81.180 ;
        RECT -259.670 -81.350 -259.350 -81.320 ;
        RECT -256.990 -81.180 -256.670 -81.070 ;
        RECT -256.330 -81.180 -256.170 -80.390 ;
        RECT -254.730 -80.540 -254.390 -80.390 ;
        RECT -252.030 -80.390 -250.090 -80.240 ;
        RECT -252.030 -80.540 -251.690 -80.390 ;
        RECT -254.710 -80.740 -254.390 -80.710 ;
        RECT -256.990 -81.320 -256.170 -81.180 ;
        RECT -255.210 -80.880 -254.390 -80.740 ;
        RECT -256.990 -81.350 -256.670 -81.320 ;
        RECT -259.690 -81.670 -259.350 -81.520 ;
        RECT -261.290 -81.820 -259.350 -81.670 ;
        RECT -256.990 -81.670 -256.650 -81.520 ;
        RECT -255.210 -81.670 -255.050 -80.880 ;
        RECT -254.710 -80.990 -254.390 -80.880 ;
        RECT -252.030 -80.740 -251.710 -80.710 ;
        RECT -252.030 -80.880 -251.210 -80.740 ;
        RECT -252.030 -80.990 -251.710 -80.880 ;
        RECT -256.990 -81.820 -255.050 -81.670 ;
        RECT -251.370 -81.670 -251.210 -80.880 ;
        RECT -250.250 -81.180 -250.090 -80.390 ;
        RECT -246.410 -80.390 -244.470 -80.240 ;
        RECT -249.750 -81.180 -249.430 -81.070 ;
        RECT -250.250 -81.320 -249.430 -81.180 ;
        RECT -249.750 -81.350 -249.430 -81.320 ;
        RECT -247.070 -81.180 -246.750 -81.070 ;
        RECT -246.410 -81.180 -246.250 -80.390 ;
        RECT -244.810 -80.540 -244.470 -80.390 ;
        RECT -242.110 -80.390 -240.170 -80.240 ;
        RECT -242.110 -80.540 -241.770 -80.390 ;
        RECT -244.790 -80.740 -244.470 -80.710 ;
        RECT -247.070 -81.320 -246.250 -81.180 ;
        RECT -245.290 -80.880 -244.470 -80.740 ;
        RECT -247.070 -81.350 -246.750 -81.320 ;
        RECT -249.770 -81.670 -249.430 -81.520 ;
        RECT -251.370 -81.820 -249.430 -81.670 ;
        RECT -247.070 -81.670 -246.730 -81.520 ;
        RECT -245.290 -81.670 -245.130 -80.880 ;
        RECT -244.790 -80.990 -244.470 -80.880 ;
        RECT -242.110 -80.740 -241.790 -80.710 ;
        RECT -242.110 -80.880 -241.290 -80.740 ;
        RECT -242.110 -80.990 -241.790 -80.880 ;
        RECT -247.070 -81.820 -245.130 -81.670 ;
        RECT -241.450 -81.670 -241.290 -80.880 ;
        RECT -240.330 -81.180 -240.170 -80.390 ;
        RECT -236.490 -80.390 -234.550 -80.240 ;
        RECT -239.830 -81.180 -239.510 -81.070 ;
        RECT -240.330 -81.320 -239.510 -81.180 ;
        RECT -239.830 -81.350 -239.510 -81.320 ;
        RECT -237.150 -81.180 -236.830 -81.070 ;
        RECT -236.490 -81.180 -236.330 -80.390 ;
        RECT -234.890 -80.540 -234.550 -80.390 ;
        RECT -232.190 -80.390 -230.250 -80.240 ;
        RECT -232.190 -80.540 -231.850 -80.390 ;
        RECT -234.870 -80.740 -234.550 -80.710 ;
        RECT -237.150 -81.320 -236.330 -81.180 ;
        RECT -235.370 -80.880 -234.550 -80.740 ;
        RECT -237.150 -81.350 -236.830 -81.320 ;
        RECT -239.850 -81.670 -239.510 -81.520 ;
        RECT -241.450 -81.820 -239.510 -81.670 ;
        RECT -237.150 -81.670 -236.810 -81.520 ;
        RECT -235.370 -81.670 -235.210 -80.880 ;
        RECT -234.870 -80.990 -234.550 -80.880 ;
        RECT -232.190 -80.740 -231.870 -80.710 ;
        RECT -232.190 -80.880 -231.370 -80.740 ;
        RECT -232.190 -80.990 -231.870 -80.880 ;
        RECT -237.150 -81.820 -235.210 -81.670 ;
        RECT -231.530 -81.670 -231.370 -80.880 ;
        RECT -230.410 -81.180 -230.250 -80.390 ;
        RECT -226.570 -80.390 -224.630 -80.240 ;
        RECT -229.910 -81.180 -229.590 -81.070 ;
        RECT -230.410 -81.320 -229.590 -81.180 ;
        RECT -229.910 -81.350 -229.590 -81.320 ;
        RECT -227.230 -81.180 -226.910 -81.070 ;
        RECT -226.570 -81.180 -226.410 -80.390 ;
        RECT -224.970 -80.540 -224.630 -80.390 ;
        RECT -222.270 -80.390 -220.330 -80.240 ;
        RECT -222.270 -80.540 -221.930 -80.390 ;
        RECT -224.950 -80.740 -224.630 -80.710 ;
        RECT -227.230 -81.320 -226.410 -81.180 ;
        RECT -225.450 -80.880 -224.630 -80.740 ;
        RECT -227.230 -81.350 -226.910 -81.320 ;
        RECT -229.930 -81.670 -229.590 -81.520 ;
        RECT -231.530 -81.820 -229.590 -81.670 ;
        RECT -227.230 -81.670 -226.890 -81.520 ;
        RECT -225.450 -81.670 -225.290 -80.880 ;
        RECT -224.950 -80.990 -224.630 -80.880 ;
        RECT -222.270 -80.740 -221.950 -80.710 ;
        RECT -222.270 -80.880 -221.450 -80.740 ;
        RECT -222.270 -80.990 -221.950 -80.880 ;
        RECT -227.230 -81.820 -225.290 -81.670 ;
        RECT -221.610 -81.670 -221.450 -80.880 ;
        RECT -220.490 -81.180 -220.330 -80.390 ;
        RECT -216.650 -80.390 -214.710 -80.240 ;
        RECT -219.990 -81.180 -219.670 -81.070 ;
        RECT -220.490 -81.320 -219.670 -81.180 ;
        RECT -219.990 -81.350 -219.670 -81.320 ;
        RECT -217.310 -81.180 -216.990 -81.070 ;
        RECT -216.650 -81.180 -216.490 -80.390 ;
        RECT -215.050 -80.540 -214.710 -80.390 ;
        RECT -212.350 -80.390 -210.410 -80.240 ;
        RECT -212.350 -80.540 -212.010 -80.390 ;
        RECT -215.030 -80.740 -214.710 -80.710 ;
        RECT -217.310 -81.320 -216.490 -81.180 ;
        RECT -215.530 -80.880 -214.710 -80.740 ;
        RECT -217.310 -81.350 -216.990 -81.320 ;
        RECT -220.010 -81.670 -219.670 -81.520 ;
        RECT -221.610 -81.820 -219.670 -81.670 ;
        RECT -217.310 -81.670 -216.970 -81.520 ;
        RECT -215.530 -81.670 -215.370 -80.880 ;
        RECT -215.030 -80.990 -214.710 -80.880 ;
        RECT -212.350 -80.740 -212.030 -80.710 ;
        RECT -212.350 -80.880 -211.530 -80.740 ;
        RECT -212.350 -80.990 -212.030 -80.880 ;
        RECT -217.310 -81.820 -215.370 -81.670 ;
        RECT -211.690 -81.670 -211.530 -80.880 ;
        RECT -210.570 -81.180 -210.410 -80.390 ;
        RECT -206.730 -80.390 -204.790 -80.240 ;
        RECT -210.070 -81.180 -209.750 -81.070 ;
        RECT -210.570 -81.320 -209.750 -81.180 ;
        RECT -210.070 -81.350 -209.750 -81.320 ;
        RECT -207.390 -81.180 -207.070 -81.070 ;
        RECT -206.730 -81.180 -206.570 -80.390 ;
        RECT -205.130 -80.540 -204.790 -80.390 ;
        RECT -202.430 -80.390 -200.490 -80.240 ;
        RECT -202.430 -80.540 -202.090 -80.390 ;
        RECT -205.110 -80.740 -204.790 -80.710 ;
        RECT -207.390 -81.320 -206.570 -81.180 ;
        RECT -205.610 -80.880 -204.790 -80.740 ;
        RECT -207.390 -81.350 -207.070 -81.320 ;
        RECT -210.090 -81.670 -209.750 -81.520 ;
        RECT -211.690 -81.820 -209.750 -81.670 ;
        RECT -207.390 -81.670 -207.050 -81.520 ;
        RECT -205.610 -81.670 -205.450 -80.880 ;
        RECT -205.110 -80.990 -204.790 -80.880 ;
        RECT -202.430 -80.740 -202.110 -80.710 ;
        RECT -202.430 -80.880 -201.610 -80.740 ;
        RECT -202.430 -80.990 -202.110 -80.880 ;
        RECT -207.390 -81.820 -205.450 -81.670 ;
        RECT -201.770 -81.670 -201.610 -80.880 ;
        RECT -200.650 -81.180 -200.490 -80.390 ;
        RECT -196.810 -80.390 -194.870 -80.240 ;
        RECT -200.150 -81.180 -199.830 -81.070 ;
        RECT -200.650 -81.320 -199.830 -81.180 ;
        RECT -200.150 -81.350 -199.830 -81.320 ;
        RECT -197.470 -81.180 -197.150 -81.070 ;
        RECT -196.810 -81.180 -196.650 -80.390 ;
        RECT -195.210 -80.540 -194.870 -80.390 ;
        RECT -192.510 -80.390 -190.570 -80.240 ;
        RECT -192.510 -80.540 -192.170 -80.390 ;
        RECT -195.190 -80.740 -194.870 -80.710 ;
        RECT -197.470 -81.320 -196.650 -81.180 ;
        RECT -195.690 -80.880 -194.870 -80.740 ;
        RECT -197.470 -81.350 -197.150 -81.320 ;
        RECT -200.170 -81.670 -199.830 -81.520 ;
        RECT -201.770 -81.820 -199.830 -81.670 ;
        RECT -197.470 -81.670 -197.130 -81.520 ;
        RECT -195.690 -81.670 -195.530 -80.880 ;
        RECT -195.190 -80.990 -194.870 -80.880 ;
        RECT -192.510 -80.740 -192.190 -80.710 ;
        RECT -192.510 -80.880 -191.690 -80.740 ;
        RECT -192.510 -80.990 -192.190 -80.880 ;
        RECT -197.470 -81.820 -195.530 -81.670 ;
        RECT -191.850 -81.670 -191.690 -80.880 ;
        RECT -190.730 -81.180 -190.570 -80.390 ;
        RECT -186.890 -80.390 -184.950 -80.240 ;
        RECT -190.230 -81.180 -189.910 -81.070 ;
        RECT -190.730 -81.320 -189.910 -81.180 ;
        RECT -190.230 -81.350 -189.910 -81.320 ;
        RECT -187.550 -81.180 -187.230 -81.070 ;
        RECT -186.890 -81.180 -186.730 -80.390 ;
        RECT -185.290 -80.540 -184.950 -80.390 ;
        RECT -182.590 -80.390 -180.650 -80.240 ;
        RECT -182.590 -80.540 -182.250 -80.390 ;
        RECT -185.270 -80.740 -184.950 -80.710 ;
        RECT -187.550 -81.320 -186.730 -81.180 ;
        RECT -185.770 -80.880 -184.950 -80.740 ;
        RECT -187.550 -81.350 -187.230 -81.320 ;
        RECT -190.250 -81.670 -189.910 -81.520 ;
        RECT -191.850 -81.820 -189.910 -81.670 ;
        RECT -187.550 -81.670 -187.210 -81.520 ;
        RECT -185.770 -81.670 -185.610 -80.880 ;
        RECT -185.270 -80.990 -184.950 -80.880 ;
        RECT -182.590 -80.740 -182.270 -80.710 ;
        RECT -182.590 -80.880 -181.770 -80.740 ;
        RECT -182.590 -80.990 -182.270 -80.880 ;
        RECT -187.550 -81.820 -185.610 -81.670 ;
        RECT -181.930 -81.670 -181.770 -80.880 ;
        RECT -180.810 -81.180 -180.650 -80.390 ;
        RECT -176.970 -80.390 -175.030 -80.240 ;
        RECT -180.310 -81.180 -179.990 -81.070 ;
        RECT -180.810 -81.320 -179.990 -81.180 ;
        RECT -180.310 -81.350 -179.990 -81.320 ;
        RECT -177.630 -81.180 -177.310 -81.070 ;
        RECT -176.970 -81.180 -176.810 -80.390 ;
        RECT -175.370 -80.540 -175.030 -80.390 ;
        RECT -172.670 -80.390 -170.730 -80.240 ;
        RECT -172.670 -80.540 -172.330 -80.390 ;
        RECT -175.350 -80.740 -175.030 -80.710 ;
        RECT -177.630 -81.320 -176.810 -81.180 ;
        RECT -175.850 -80.880 -175.030 -80.740 ;
        RECT -177.630 -81.350 -177.310 -81.320 ;
        RECT -180.330 -81.670 -179.990 -81.520 ;
        RECT -181.930 -81.820 -179.990 -81.670 ;
        RECT -177.630 -81.670 -177.290 -81.520 ;
        RECT -175.850 -81.670 -175.690 -80.880 ;
        RECT -175.350 -80.990 -175.030 -80.880 ;
        RECT -172.670 -80.740 -172.350 -80.710 ;
        RECT -172.670 -80.880 -171.850 -80.740 ;
        RECT -172.670 -80.990 -172.350 -80.880 ;
        RECT -177.630 -81.820 -175.690 -81.670 ;
        RECT -172.010 -81.670 -171.850 -80.880 ;
        RECT -170.890 -81.180 -170.730 -80.390 ;
        RECT -167.050 -80.390 -165.110 -80.240 ;
        RECT -170.390 -81.180 -170.070 -81.070 ;
        RECT -170.890 -81.320 -170.070 -81.180 ;
        RECT -170.390 -81.350 -170.070 -81.320 ;
        RECT -167.710 -81.180 -167.390 -81.070 ;
        RECT -167.050 -81.180 -166.890 -80.390 ;
        RECT -165.450 -80.540 -165.110 -80.390 ;
        RECT -162.750 -80.390 -160.810 -80.240 ;
        RECT -162.750 -80.540 -162.410 -80.390 ;
        RECT -165.430 -80.740 -165.110 -80.710 ;
        RECT -167.710 -81.320 -166.890 -81.180 ;
        RECT -165.930 -80.880 -165.110 -80.740 ;
        RECT -167.710 -81.350 -167.390 -81.320 ;
        RECT -170.410 -81.670 -170.070 -81.520 ;
        RECT -172.010 -81.820 -170.070 -81.670 ;
        RECT -167.710 -81.670 -167.370 -81.520 ;
        RECT -165.930 -81.670 -165.770 -80.880 ;
        RECT -165.430 -80.990 -165.110 -80.880 ;
        RECT -162.750 -80.740 -162.430 -80.710 ;
        RECT -162.750 -80.880 -161.930 -80.740 ;
        RECT -162.750 -80.990 -162.430 -80.880 ;
        RECT -167.710 -81.820 -165.770 -81.670 ;
        RECT -162.090 -81.670 -161.930 -80.880 ;
        RECT -160.970 -81.180 -160.810 -80.390 ;
        RECT -157.130 -80.390 -155.190 -80.240 ;
        RECT -160.470 -81.180 -160.150 -81.070 ;
        RECT -160.970 -81.320 -160.150 -81.180 ;
        RECT -160.470 -81.350 -160.150 -81.320 ;
        RECT -157.790 -81.180 -157.470 -81.070 ;
        RECT -157.130 -81.180 -156.970 -80.390 ;
        RECT -155.530 -80.540 -155.190 -80.390 ;
        RECT -152.830 -80.390 -150.890 -80.240 ;
        RECT -152.830 -80.540 -152.490 -80.390 ;
        RECT -155.510 -80.740 -155.190 -80.710 ;
        RECT -157.790 -81.320 -156.970 -81.180 ;
        RECT -156.010 -80.880 -155.190 -80.740 ;
        RECT -157.790 -81.350 -157.470 -81.320 ;
        RECT -160.490 -81.670 -160.150 -81.520 ;
        RECT -162.090 -81.820 -160.150 -81.670 ;
        RECT -157.790 -81.670 -157.450 -81.520 ;
        RECT -156.010 -81.670 -155.850 -80.880 ;
        RECT -155.510 -80.990 -155.190 -80.880 ;
        RECT -152.830 -80.740 -152.510 -80.710 ;
        RECT -152.830 -80.880 -152.010 -80.740 ;
        RECT -152.830 -80.990 -152.510 -80.880 ;
        RECT -157.790 -81.820 -155.850 -81.670 ;
        RECT -152.170 -81.670 -152.010 -80.880 ;
        RECT -151.050 -81.180 -150.890 -80.390 ;
        RECT -147.210 -80.390 -145.270 -80.240 ;
        RECT -150.550 -81.180 -150.230 -81.070 ;
        RECT -151.050 -81.320 -150.230 -81.180 ;
        RECT -150.550 -81.350 -150.230 -81.320 ;
        RECT -147.870 -81.180 -147.550 -81.070 ;
        RECT -147.210 -81.180 -147.050 -80.390 ;
        RECT -145.610 -80.540 -145.270 -80.390 ;
        RECT -142.910 -80.390 -140.970 -80.240 ;
        RECT -142.910 -80.540 -142.570 -80.390 ;
        RECT -145.590 -80.740 -145.270 -80.710 ;
        RECT -147.870 -81.320 -147.050 -81.180 ;
        RECT -146.090 -80.880 -145.270 -80.740 ;
        RECT -147.870 -81.350 -147.550 -81.320 ;
        RECT -150.570 -81.670 -150.230 -81.520 ;
        RECT -152.170 -81.820 -150.230 -81.670 ;
        RECT -147.870 -81.670 -147.530 -81.520 ;
        RECT -146.090 -81.670 -145.930 -80.880 ;
        RECT -145.590 -80.990 -145.270 -80.880 ;
        RECT -142.910 -80.740 -142.590 -80.710 ;
        RECT -142.910 -80.880 -142.090 -80.740 ;
        RECT -142.910 -80.990 -142.590 -80.880 ;
        RECT -147.870 -81.820 -145.930 -81.670 ;
        RECT -142.250 -81.670 -142.090 -80.880 ;
        RECT -141.130 -81.180 -140.970 -80.390 ;
        RECT -137.290 -80.390 -135.350 -80.240 ;
        RECT -140.630 -81.180 -140.310 -81.070 ;
        RECT -141.130 -81.320 -140.310 -81.180 ;
        RECT -140.630 -81.350 -140.310 -81.320 ;
        RECT -137.950 -81.180 -137.630 -81.070 ;
        RECT -137.290 -81.180 -137.130 -80.390 ;
        RECT -135.690 -80.540 -135.350 -80.390 ;
        RECT -132.990 -80.390 -131.050 -80.240 ;
        RECT -132.990 -80.540 -132.650 -80.390 ;
        RECT -135.670 -80.740 -135.350 -80.710 ;
        RECT -137.950 -81.320 -137.130 -81.180 ;
        RECT -136.170 -80.880 -135.350 -80.740 ;
        RECT -137.950 -81.350 -137.630 -81.320 ;
        RECT -140.650 -81.670 -140.310 -81.520 ;
        RECT -142.250 -81.820 -140.310 -81.670 ;
        RECT -137.950 -81.670 -137.610 -81.520 ;
        RECT -136.170 -81.670 -136.010 -80.880 ;
        RECT -135.670 -80.990 -135.350 -80.880 ;
        RECT -132.990 -80.740 -132.670 -80.710 ;
        RECT -132.990 -80.880 -132.170 -80.740 ;
        RECT -132.990 -80.990 -132.670 -80.880 ;
        RECT -137.950 -81.820 -136.010 -81.670 ;
        RECT -132.330 -81.670 -132.170 -80.880 ;
        RECT -131.210 -81.180 -131.050 -80.390 ;
        RECT -127.370 -80.390 -125.430 -80.240 ;
        RECT -130.710 -81.180 -130.390 -81.070 ;
        RECT -131.210 -81.320 -130.390 -81.180 ;
        RECT -130.710 -81.350 -130.390 -81.320 ;
        RECT -128.030 -81.180 -127.710 -81.070 ;
        RECT -127.370 -81.180 -127.210 -80.390 ;
        RECT -125.770 -80.540 -125.430 -80.390 ;
        RECT -123.070 -80.390 -121.130 -80.240 ;
        RECT -123.070 -80.540 -122.730 -80.390 ;
        RECT -125.750 -80.740 -125.430 -80.710 ;
        RECT -128.030 -81.320 -127.210 -81.180 ;
        RECT -126.250 -80.880 -125.430 -80.740 ;
        RECT -128.030 -81.350 -127.710 -81.320 ;
        RECT -130.730 -81.670 -130.390 -81.520 ;
        RECT -132.330 -81.820 -130.390 -81.670 ;
        RECT -128.030 -81.670 -127.690 -81.520 ;
        RECT -126.250 -81.670 -126.090 -80.880 ;
        RECT -125.750 -80.990 -125.430 -80.880 ;
        RECT -123.070 -80.740 -122.750 -80.710 ;
        RECT -123.070 -80.880 -122.250 -80.740 ;
        RECT -123.070 -80.990 -122.750 -80.880 ;
        RECT -128.030 -81.820 -126.090 -81.670 ;
        RECT -122.410 -81.670 -122.250 -80.880 ;
        RECT -121.290 -81.180 -121.130 -80.390 ;
        RECT -117.450 -80.390 -115.510 -80.240 ;
        RECT -120.790 -81.180 -120.470 -81.070 ;
        RECT -121.290 -81.320 -120.470 -81.180 ;
        RECT -120.790 -81.350 -120.470 -81.320 ;
        RECT -118.110 -81.180 -117.790 -81.070 ;
        RECT -117.450 -81.180 -117.290 -80.390 ;
        RECT -115.850 -80.540 -115.510 -80.390 ;
        RECT -113.150 -80.390 -111.210 -80.240 ;
        RECT -113.150 -80.540 -112.810 -80.390 ;
        RECT -115.830 -80.740 -115.510 -80.710 ;
        RECT -118.110 -81.320 -117.290 -81.180 ;
        RECT -116.330 -80.880 -115.510 -80.740 ;
        RECT -118.110 -81.350 -117.790 -81.320 ;
        RECT -120.810 -81.670 -120.470 -81.520 ;
        RECT -122.410 -81.820 -120.470 -81.670 ;
        RECT -118.110 -81.670 -117.770 -81.520 ;
        RECT -116.330 -81.670 -116.170 -80.880 ;
        RECT -115.830 -80.990 -115.510 -80.880 ;
        RECT -113.150 -80.740 -112.830 -80.710 ;
        RECT -113.150 -80.880 -112.330 -80.740 ;
        RECT -113.150 -80.990 -112.830 -80.880 ;
        RECT -118.110 -81.820 -116.170 -81.670 ;
        RECT -112.490 -81.670 -112.330 -80.880 ;
        RECT -111.370 -81.180 -111.210 -80.390 ;
        RECT -107.530 -80.390 -105.590 -80.240 ;
        RECT -110.870 -81.180 -110.550 -81.070 ;
        RECT -111.370 -81.320 -110.550 -81.180 ;
        RECT -110.870 -81.350 -110.550 -81.320 ;
        RECT -108.190 -81.180 -107.870 -81.070 ;
        RECT -107.530 -81.180 -107.370 -80.390 ;
        RECT -105.930 -80.540 -105.590 -80.390 ;
        RECT -103.230 -80.390 -101.290 -80.240 ;
        RECT -103.230 -80.540 -102.890 -80.390 ;
        RECT -105.910 -80.740 -105.590 -80.710 ;
        RECT -108.190 -81.320 -107.370 -81.180 ;
        RECT -106.410 -80.880 -105.590 -80.740 ;
        RECT -108.190 -81.350 -107.870 -81.320 ;
        RECT -110.890 -81.670 -110.550 -81.520 ;
        RECT -112.490 -81.820 -110.550 -81.670 ;
        RECT -108.190 -81.670 -107.850 -81.520 ;
        RECT -106.410 -81.670 -106.250 -80.880 ;
        RECT -105.910 -80.990 -105.590 -80.880 ;
        RECT -103.230 -80.740 -102.910 -80.710 ;
        RECT -103.230 -80.880 -102.410 -80.740 ;
        RECT -103.230 -80.990 -102.910 -80.880 ;
        RECT -108.190 -81.820 -106.250 -81.670 ;
        RECT -102.570 -81.670 -102.410 -80.880 ;
        RECT -101.450 -81.180 -101.290 -80.390 ;
        RECT -97.610 -80.390 -95.670 -80.240 ;
        RECT -100.950 -81.180 -100.630 -81.070 ;
        RECT -101.450 -81.320 -100.630 -81.180 ;
        RECT -100.950 -81.350 -100.630 -81.320 ;
        RECT -98.270 -81.180 -97.950 -81.070 ;
        RECT -97.610 -81.180 -97.450 -80.390 ;
        RECT -96.010 -80.540 -95.670 -80.390 ;
        RECT -93.310 -80.390 -91.370 -80.240 ;
        RECT -93.310 -80.540 -92.970 -80.390 ;
        RECT -95.990 -80.740 -95.670 -80.710 ;
        RECT -98.270 -81.320 -97.450 -81.180 ;
        RECT -96.490 -80.880 -95.670 -80.740 ;
        RECT -98.270 -81.350 -97.950 -81.320 ;
        RECT -100.970 -81.670 -100.630 -81.520 ;
        RECT -102.570 -81.820 -100.630 -81.670 ;
        RECT -98.270 -81.670 -97.930 -81.520 ;
        RECT -96.490 -81.670 -96.330 -80.880 ;
        RECT -95.990 -80.990 -95.670 -80.880 ;
        RECT -93.310 -80.740 -92.990 -80.710 ;
        RECT -93.310 -80.880 -92.490 -80.740 ;
        RECT -93.310 -80.990 -92.990 -80.880 ;
        RECT -98.270 -81.820 -96.330 -81.670 ;
        RECT -92.650 -81.670 -92.490 -80.880 ;
        RECT -91.530 -81.180 -91.370 -80.390 ;
        RECT -87.690 -80.390 -85.750 -80.240 ;
        RECT -91.030 -81.180 -90.710 -81.070 ;
        RECT -91.530 -81.320 -90.710 -81.180 ;
        RECT -91.030 -81.350 -90.710 -81.320 ;
        RECT -88.350 -81.180 -88.030 -81.070 ;
        RECT -87.690 -81.180 -87.530 -80.390 ;
        RECT -86.090 -80.540 -85.750 -80.390 ;
        RECT -83.390 -80.390 -81.450 -80.240 ;
        RECT -83.390 -80.540 -83.050 -80.390 ;
        RECT -86.070 -80.740 -85.750 -80.710 ;
        RECT -88.350 -81.320 -87.530 -81.180 ;
        RECT -86.570 -80.880 -85.750 -80.740 ;
        RECT -88.350 -81.350 -88.030 -81.320 ;
        RECT -91.050 -81.670 -90.710 -81.520 ;
        RECT -92.650 -81.820 -90.710 -81.670 ;
        RECT -88.350 -81.670 -88.010 -81.520 ;
        RECT -86.570 -81.670 -86.410 -80.880 ;
        RECT -86.070 -80.990 -85.750 -80.880 ;
        RECT -83.390 -80.740 -83.070 -80.710 ;
        RECT -83.390 -80.880 -82.570 -80.740 ;
        RECT -83.390 -80.990 -83.070 -80.880 ;
        RECT -88.350 -81.820 -86.410 -81.670 ;
        RECT -82.730 -81.670 -82.570 -80.880 ;
        RECT -81.610 -81.180 -81.450 -80.390 ;
        RECT -77.770 -80.390 -75.830 -80.240 ;
        RECT -81.110 -81.180 -80.790 -81.070 ;
        RECT -81.610 -81.320 -80.790 -81.180 ;
        RECT -81.110 -81.350 -80.790 -81.320 ;
        RECT -78.430 -81.180 -78.110 -81.070 ;
        RECT -77.770 -81.180 -77.610 -80.390 ;
        RECT -76.170 -80.540 -75.830 -80.390 ;
        RECT -73.470 -80.390 -71.530 -80.240 ;
        RECT -73.470 -80.540 -73.130 -80.390 ;
        RECT -76.150 -80.740 -75.830 -80.710 ;
        RECT -78.430 -81.320 -77.610 -81.180 ;
        RECT -76.650 -80.880 -75.830 -80.740 ;
        RECT -78.430 -81.350 -78.110 -81.320 ;
        RECT -81.130 -81.670 -80.790 -81.520 ;
        RECT -82.730 -81.820 -80.790 -81.670 ;
        RECT -78.430 -81.670 -78.090 -81.520 ;
        RECT -76.650 -81.670 -76.490 -80.880 ;
        RECT -76.150 -80.990 -75.830 -80.880 ;
        RECT -73.470 -80.740 -73.150 -80.710 ;
        RECT -73.470 -80.880 -72.650 -80.740 ;
        RECT -73.470 -80.990 -73.150 -80.880 ;
        RECT -78.430 -81.820 -76.490 -81.670 ;
        RECT -72.810 -81.670 -72.650 -80.880 ;
        RECT -71.690 -81.180 -71.530 -80.390 ;
        RECT -67.850 -80.390 -65.910 -80.240 ;
        RECT -71.190 -81.180 -70.870 -81.070 ;
        RECT -71.690 -81.320 -70.870 -81.180 ;
        RECT -71.190 -81.350 -70.870 -81.320 ;
        RECT -68.510 -81.180 -68.190 -81.070 ;
        RECT -67.850 -81.180 -67.690 -80.390 ;
        RECT -66.250 -80.540 -65.910 -80.390 ;
        RECT -63.550 -80.390 -61.610 -80.240 ;
        RECT -63.550 -80.540 -63.210 -80.390 ;
        RECT -66.230 -80.740 -65.910 -80.710 ;
        RECT -68.510 -81.320 -67.690 -81.180 ;
        RECT -66.730 -80.880 -65.910 -80.740 ;
        RECT -68.510 -81.350 -68.190 -81.320 ;
        RECT -71.210 -81.670 -70.870 -81.520 ;
        RECT -72.810 -81.820 -70.870 -81.670 ;
        RECT -68.510 -81.670 -68.170 -81.520 ;
        RECT -66.730 -81.670 -66.570 -80.880 ;
        RECT -66.230 -80.990 -65.910 -80.880 ;
        RECT -63.550 -80.740 -63.230 -80.710 ;
        RECT -63.550 -80.880 -62.730 -80.740 ;
        RECT -63.550 -80.990 -63.230 -80.880 ;
        RECT -68.510 -81.820 -66.570 -81.670 ;
        RECT -62.890 -81.670 -62.730 -80.880 ;
        RECT -61.770 -81.180 -61.610 -80.390 ;
        RECT -57.930 -80.390 -55.990 -80.240 ;
        RECT -61.270 -81.180 -60.950 -81.070 ;
        RECT -61.770 -81.320 -60.950 -81.180 ;
        RECT -61.270 -81.350 -60.950 -81.320 ;
        RECT -58.590 -81.180 -58.270 -81.070 ;
        RECT -57.930 -81.180 -57.770 -80.390 ;
        RECT -56.330 -80.540 -55.990 -80.390 ;
        RECT -53.630 -80.390 -51.690 -80.240 ;
        RECT -53.630 -80.540 -53.290 -80.390 ;
        RECT -56.310 -80.740 -55.990 -80.710 ;
        RECT -58.590 -81.320 -57.770 -81.180 ;
        RECT -56.810 -80.880 -55.990 -80.740 ;
        RECT -58.590 -81.350 -58.270 -81.320 ;
        RECT -61.290 -81.670 -60.950 -81.520 ;
        RECT -62.890 -81.820 -60.950 -81.670 ;
        RECT -58.590 -81.670 -58.250 -81.520 ;
        RECT -56.810 -81.670 -56.650 -80.880 ;
        RECT -56.310 -80.990 -55.990 -80.880 ;
        RECT -53.630 -80.740 -53.310 -80.710 ;
        RECT -53.630 -80.880 -52.810 -80.740 ;
        RECT -53.630 -80.990 -53.310 -80.880 ;
        RECT -58.590 -81.820 -56.650 -81.670 ;
        RECT -52.970 -81.670 -52.810 -80.880 ;
        RECT -51.850 -81.180 -51.690 -80.390 ;
        RECT -48.010 -80.390 -46.070 -80.240 ;
        RECT -51.350 -81.180 -51.030 -81.070 ;
        RECT -51.850 -81.320 -51.030 -81.180 ;
        RECT -51.350 -81.350 -51.030 -81.320 ;
        RECT -48.670 -81.180 -48.350 -81.070 ;
        RECT -48.010 -81.180 -47.850 -80.390 ;
        RECT -46.410 -80.540 -46.070 -80.390 ;
        RECT -43.710 -80.390 -41.770 -80.240 ;
        RECT -43.710 -80.540 -43.370 -80.390 ;
        RECT -46.390 -80.740 -46.070 -80.710 ;
        RECT -48.670 -81.320 -47.850 -81.180 ;
        RECT -46.890 -80.880 -46.070 -80.740 ;
        RECT -48.670 -81.350 -48.350 -81.320 ;
        RECT -51.370 -81.670 -51.030 -81.520 ;
        RECT -52.970 -81.820 -51.030 -81.670 ;
        RECT -48.670 -81.670 -48.330 -81.520 ;
        RECT -46.890 -81.670 -46.730 -80.880 ;
        RECT -46.390 -80.990 -46.070 -80.880 ;
        RECT -43.710 -80.740 -43.390 -80.710 ;
        RECT -43.710 -80.880 -42.890 -80.740 ;
        RECT -43.710 -80.990 -43.390 -80.880 ;
        RECT -48.670 -81.820 -46.730 -81.670 ;
        RECT -43.050 -81.670 -42.890 -80.880 ;
        RECT -41.930 -81.180 -41.770 -80.390 ;
        RECT -38.090 -80.390 -36.150 -80.240 ;
        RECT -41.430 -81.180 -41.110 -81.070 ;
        RECT -41.930 -81.320 -41.110 -81.180 ;
        RECT -41.430 -81.350 -41.110 -81.320 ;
        RECT -38.750 -81.180 -38.430 -81.070 ;
        RECT -38.090 -81.180 -37.930 -80.390 ;
        RECT -36.490 -80.540 -36.150 -80.390 ;
        RECT -33.790 -80.390 -31.850 -80.240 ;
        RECT -33.790 -80.540 -33.450 -80.390 ;
        RECT -36.470 -80.740 -36.150 -80.710 ;
        RECT -38.750 -81.320 -37.930 -81.180 ;
        RECT -36.970 -80.880 -36.150 -80.740 ;
        RECT -38.750 -81.350 -38.430 -81.320 ;
        RECT -41.450 -81.670 -41.110 -81.520 ;
        RECT -43.050 -81.820 -41.110 -81.670 ;
        RECT -38.750 -81.670 -38.410 -81.520 ;
        RECT -36.970 -81.670 -36.810 -80.880 ;
        RECT -36.470 -80.990 -36.150 -80.880 ;
        RECT -33.790 -80.740 -33.470 -80.710 ;
        RECT -33.790 -80.880 -32.970 -80.740 ;
        RECT -33.790 -80.990 -33.470 -80.880 ;
        RECT -38.750 -81.820 -36.810 -81.670 ;
        RECT -33.130 -81.670 -32.970 -80.880 ;
        RECT -32.010 -81.180 -31.850 -80.390 ;
        RECT -28.170 -80.390 -26.230 -80.240 ;
        RECT -31.510 -81.180 -31.190 -81.070 ;
        RECT -32.010 -81.320 -31.190 -81.180 ;
        RECT -31.510 -81.350 -31.190 -81.320 ;
        RECT -28.830 -81.180 -28.510 -81.070 ;
        RECT -28.170 -81.180 -28.010 -80.390 ;
        RECT -26.570 -80.540 -26.230 -80.390 ;
        RECT -23.870 -80.390 -21.930 -80.240 ;
        RECT -23.870 -80.540 -23.530 -80.390 ;
        RECT -26.550 -80.740 -26.230 -80.710 ;
        RECT -28.830 -81.320 -28.010 -81.180 ;
        RECT -27.050 -80.880 -26.230 -80.740 ;
        RECT -28.830 -81.350 -28.510 -81.320 ;
        RECT -31.530 -81.670 -31.190 -81.520 ;
        RECT -33.130 -81.820 -31.190 -81.670 ;
        RECT -28.830 -81.670 -28.490 -81.520 ;
        RECT -27.050 -81.670 -26.890 -80.880 ;
        RECT -26.550 -80.990 -26.230 -80.880 ;
        RECT -23.870 -80.740 -23.550 -80.710 ;
        RECT -23.870 -80.880 -23.050 -80.740 ;
        RECT -23.870 -80.990 -23.550 -80.880 ;
        RECT -28.830 -81.820 -26.890 -81.670 ;
        RECT -23.210 -81.670 -23.050 -80.880 ;
        RECT -22.090 -81.180 -21.930 -80.390 ;
        RECT -18.250 -80.390 -16.310 -80.240 ;
        RECT -21.590 -81.180 -21.270 -81.070 ;
        RECT -22.090 -81.320 -21.270 -81.180 ;
        RECT -21.590 -81.350 -21.270 -81.320 ;
        RECT -18.910 -81.180 -18.590 -81.070 ;
        RECT -18.250 -81.180 -18.090 -80.390 ;
        RECT -16.650 -80.540 -16.310 -80.390 ;
        RECT -13.950 -80.390 -12.010 -80.240 ;
        RECT -13.950 -80.540 -13.610 -80.390 ;
        RECT -16.630 -80.740 -16.310 -80.710 ;
        RECT -18.910 -81.320 -18.090 -81.180 ;
        RECT -17.130 -80.880 -16.310 -80.740 ;
        RECT -18.910 -81.350 -18.590 -81.320 ;
        RECT -21.610 -81.670 -21.270 -81.520 ;
        RECT -23.210 -81.820 -21.270 -81.670 ;
        RECT -18.910 -81.670 -18.570 -81.520 ;
        RECT -17.130 -81.670 -16.970 -80.880 ;
        RECT -16.630 -80.990 -16.310 -80.880 ;
        RECT -13.950 -80.740 -13.630 -80.710 ;
        RECT -13.950 -80.880 -13.130 -80.740 ;
        RECT -13.950 -80.990 -13.630 -80.880 ;
        RECT -18.910 -81.820 -16.970 -81.670 ;
        RECT -13.290 -81.670 -13.130 -80.880 ;
        RECT -12.170 -81.180 -12.010 -80.390 ;
        RECT -8.330 -80.390 -6.390 -80.240 ;
        RECT -11.670 -81.180 -11.350 -81.070 ;
        RECT -12.170 -81.320 -11.350 -81.180 ;
        RECT -11.670 -81.350 -11.350 -81.320 ;
        RECT -8.990 -81.180 -8.670 -81.070 ;
        RECT -8.330 -81.180 -8.170 -80.390 ;
        RECT -6.730 -80.540 -6.390 -80.390 ;
        RECT -4.030 -80.390 -2.090 -80.240 ;
        RECT -4.030 -80.540 -3.690 -80.390 ;
        RECT -6.710 -80.740 -6.390 -80.710 ;
        RECT -8.990 -81.320 -8.170 -81.180 ;
        RECT -7.210 -80.880 -6.390 -80.740 ;
        RECT -8.990 -81.350 -8.670 -81.320 ;
        RECT -11.690 -81.670 -11.350 -81.520 ;
        RECT -13.290 -81.820 -11.350 -81.670 ;
        RECT -8.990 -81.670 -8.650 -81.520 ;
        RECT -7.210 -81.670 -7.050 -80.880 ;
        RECT -6.710 -80.990 -6.390 -80.880 ;
        RECT -4.030 -80.740 -3.710 -80.710 ;
        RECT -4.030 -80.880 -3.210 -80.740 ;
        RECT -4.030 -80.990 -3.710 -80.880 ;
        RECT -8.990 -81.820 -7.050 -81.670 ;
        RECT -3.370 -81.670 -3.210 -80.880 ;
        RECT -2.250 -81.180 -2.090 -80.390 ;
        RECT 1.590 -80.390 3.530 -80.240 ;
        RECT -1.750 -81.180 -1.430 -81.070 ;
        RECT -2.250 -81.320 -1.430 -81.180 ;
        RECT -1.750 -81.350 -1.430 -81.320 ;
        RECT 0.930 -81.180 1.250 -81.070 ;
        RECT 1.590 -81.180 1.750 -80.390 ;
        RECT 3.190 -80.540 3.530 -80.390 ;
        RECT 5.890 -80.390 7.830 -80.240 ;
        RECT 5.890 -80.540 6.230 -80.390 ;
        RECT 3.210 -80.740 3.530 -80.710 ;
        RECT 0.930 -81.320 1.750 -81.180 ;
        RECT 2.710 -80.880 3.530 -80.740 ;
        RECT 0.930 -81.350 1.250 -81.320 ;
        RECT -1.770 -81.670 -1.430 -81.520 ;
        RECT -3.370 -81.820 -1.430 -81.670 ;
        RECT 0.930 -81.670 1.270 -81.520 ;
        RECT 2.710 -81.670 2.870 -80.880 ;
        RECT 3.210 -80.990 3.530 -80.880 ;
        RECT 5.890 -80.740 6.210 -80.710 ;
        RECT 5.890 -80.880 6.710 -80.740 ;
        RECT 5.890 -80.990 6.210 -80.880 ;
        RECT 0.930 -81.820 2.870 -81.670 ;
        RECT 6.550 -81.670 6.710 -80.880 ;
        RECT 7.670 -81.180 7.830 -80.390 ;
        RECT 11.510 -80.390 13.450 -80.240 ;
        RECT 8.170 -81.180 8.490 -81.070 ;
        RECT 7.670 -81.320 8.490 -81.180 ;
        RECT 8.170 -81.350 8.490 -81.320 ;
        RECT 10.850 -81.180 11.170 -81.070 ;
        RECT 11.510 -81.180 11.670 -80.390 ;
        RECT 13.110 -80.540 13.450 -80.390 ;
        RECT 15.810 -80.390 17.750 -80.240 ;
        RECT 15.810 -80.540 16.150 -80.390 ;
        RECT 13.130 -80.740 13.450 -80.710 ;
        RECT 10.850 -81.320 11.670 -81.180 ;
        RECT 12.630 -80.880 13.450 -80.740 ;
        RECT 10.850 -81.350 11.170 -81.320 ;
        RECT 8.150 -81.670 8.490 -81.520 ;
        RECT 6.550 -81.820 8.490 -81.670 ;
        RECT 10.850 -81.670 11.190 -81.520 ;
        RECT 12.630 -81.670 12.790 -80.880 ;
        RECT 13.130 -80.990 13.450 -80.880 ;
        RECT 15.810 -80.740 16.130 -80.710 ;
        RECT 15.810 -80.880 16.630 -80.740 ;
        RECT 15.810 -80.990 16.130 -80.880 ;
        RECT 10.850 -81.820 12.790 -81.670 ;
        RECT 16.470 -81.670 16.630 -80.880 ;
        RECT 17.590 -81.180 17.750 -80.390 ;
        RECT 21.430 -80.390 23.370 -80.240 ;
        RECT 18.090 -81.180 18.410 -81.070 ;
        RECT 17.590 -81.320 18.410 -81.180 ;
        RECT 18.090 -81.350 18.410 -81.320 ;
        RECT 20.770 -81.180 21.090 -81.070 ;
        RECT 21.430 -81.180 21.590 -80.390 ;
        RECT 23.030 -80.540 23.370 -80.390 ;
        RECT 23.050 -80.740 23.370 -80.710 ;
        RECT 20.770 -81.320 21.590 -81.180 ;
        RECT 22.550 -80.880 23.370 -80.740 ;
        RECT 20.770 -81.350 21.090 -81.320 ;
        RECT 18.070 -81.670 18.410 -81.520 ;
        RECT 16.470 -81.820 18.410 -81.670 ;
        RECT 20.770 -81.670 21.110 -81.520 ;
        RECT 22.550 -81.670 22.710 -80.880 ;
        RECT 23.050 -80.990 23.370 -80.880 ;
        RECT 20.770 -81.820 22.710 -81.670 ;
        RECT -293.120 -82.630 -291.280 -82.150 ;
        RECT -291.360 -83.720 -290.880 -82.820 ;
        RECT -290.060 -82.950 -289.870 -81.820 ;
        RECT -285.990 -82.950 -285.800 -81.820 ;
        RECT -280.140 -82.950 -279.950 -81.820 ;
        RECT -276.070 -82.950 -275.880 -81.820 ;
        RECT -270.220 -82.950 -270.030 -81.820 ;
        RECT -266.150 -82.950 -265.960 -81.820 ;
        RECT -260.300 -82.950 -260.110 -81.820 ;
        RECT -256.230 -82.950 -256.040 -81.820 ;
        RECT -250.380 -82.950 -250.190 -81.820 ;
        RECT -246.310 -82.950 -246.120 -81.820 ;
        RECT -240.460 -82.950 -240.270 -81.820 ;
        RECT -236.390 -82.950 -236.200 -81.820 ;
        RECT -230.540 -82.950 -230.350 -81.820 ;
        RECT -226.470 -82.950 -226.280 -81.820 ;
        RECT -220.620 -82.950 -220.430 -81.820 ;
        RECT -216.550 -82.950 -216.360 -81.820 ;
        RECT -210.700 -82.950 -210.510 -81.820 ;
        RECT -206.630 -82.950 -206.440 -81.820 ;
        RECT -200.780 -82.950 -200.590 -81.820 ;
        RECT -196.710 -82.950 -196.520 -81.820 ;
        RECT -190.860 -82.950 -190.670 -81.820 ;
        RECT -186.790 -82.950 -186.600 -81.820 ;
        RECT -180.940 -82.950 -180.750 -81.820 ;
        RECT -176.870 -82.950 -176.680 -81.820 ;
        RECT -171.020 -82.950 -170.830 -81.820 ;
        RECT -166.950 -82.950 -166.760 -81.820 ;
        RECT -161.100 -82.950 -160.910 -81.820 ;
        RECT -157.030 -82.950 -156.840 -81.820 ;
        RECT -151.180 -82.950 -150.990 -81.820 ;
        RECT -147.110 -82.950 -146.920 -81.820 ;
        RECT -141.260 -82.950 -141.070 -81.820 ;
        RECT -137.190 -82.950 -137.000 -81.820 ;
        RECT -131.340 -82.950 -131.150 -81.820 ;
        RECT -127.270 -82.950 -127.080 -81.820 ;
        RECT -121.420 -82.950 -121.230 -81.820 ;
        RECT -117.350 -82.950 -117.160 -81.820 ;
        RECT -111.500 -82.950 -111.310 -81.820 ;
        RECT -107.430 -82.950 -107.240 -81.820 ;
        RECT -101.580 -82.950 -101.390 -81.820 ;
        RECT -97.510 -82.950 -97.320 -81.820 ;
        RECT -91.660 -82.950 -91.470 -81.820 ;
        RECT -87.590 -82.950 -87.400 -81.820 ;
        RECT -81.740 -82.950 -81.550 -81.820 ;
        RECT -77.670 -82.950 -77.480 -81.820 ;
        RECT -71.820 -82.950 -71.630 -81.820 ;
        RECT -67.750 -82.950 -67.560 -81.820 ;
        RECT -61.900 -82.950 -61.710 -81.820 ;
        RECT -57.830 -82.950 -57.640 -81.820 ;
        RECT -51.980 -82.950 -51.790 -81.820 ;
        RECT -47.910 -82.950 -47.720 -81.820 ;
        RECT -42.060 -82.950 -41.870 -81.820 ;
        RECT -37.990 -82.950 -37.800 -81.820 ;
        RECT -32.140 -82.950 -31.950 -81.820 ;
        RECT -28.070 -82.950 -27.880 -81.820 ;
        RECT -22.220 -82.950 -22.030 -81.820 ;
        RECT -18.150 -82.950 -17.960 -81.820 ;
        RECT -12.300 -82.950 -12.110 -81.820 ;
        RECT -8.230 -82.950 -8.040 -81.820 ;
        RECT -2.380 -82.950 -2.190 -81.820 ;
        RECT 1.690 -82.950 1.880 -81.820 ;
        RECT 7.540 -82.950 7.730 -81.820 ;
        RECT 11.610 -82.950 11.800 -81.820 ;
        RECT 17.460 -82.950 17.650 -81.820 ;
        RECT 21.530 -82.950 21.720 -81.820 ;
        RECT -290.110 -83.240 -289.790 -82.950 ;
        RECT -286.070 -83.240 -285.750 -82.950 ;
        RECT -280.190 -83.240 -279.870 -82.950 ;
        RECT -276.150 -83.240 -275.830 -82.950 ;
        RECT -270.270 -83.240 -269.950 -82.950 ;
        RECT -266.230 -83.240 -265.910 -82.950 ;
        RECT -260.350 -83.240 -260.030 -82.950 ;
        RECT -256.310 -83.240 -255.990 -82.950 ;
        RECT -250.430 -83.240 -250.110 -82.950 ;
        RECT -246.390 -83.240 -246.070 -82.950 ;
        RECT -240.510 -83.240 -240.190 -82.950 ;
        RECT -236.470 -83.240 -236.150 -82.950 ;
        RECT -230.590 -83.240 -230.270 -82.950 ;
        RECT -226.550 -83.240 -226.230 -82.950 ;
        RECT -220.670 -83.240 -220.350 -82.950 ;
        RECT -216.630 -83.240 -216.310 -82.950 ;
        RECT -210.750 -83.240 -210.430 -82.950 ;
        RECT -206.710 -83.240 -206.390 -82.950 ;
        RECT -200.830 -83.240 -200.510 -82.950 ;
        RECT -196.790 -83.240 -196.470 -82.950 ;
        RECT -190.910 -83.240 -190.590 -82.950 ;
        RECT -186.870 -83.240 -186.550 -82.950 ;
        RECT -180.990 -83.240 -180.670 -82.950 ;
        RECT -176.950 -83.240 -176.630 -82.950 ;
        RECT -171.070 -83.240 -170.750 -82.950 ;
        RECT -167.030 -83.240 -166.710 -82.950 ;
        RECT -161.150 -83.240 -160.830 -82.950 ;
        RECT -157.110 -83.240 -156.790 -82.950 ;
        RECT -151.230 -83.240 -150.910 -82.950 ;
        RECT -147.190 -83.240 -146.870 -82.950 ;
        RECT -141.310 -83.240 -140.990 -82.950 ;
        RECT -137.270 -83.240 -136.950 -82.950 ;
        RECT -131.390 -83.240 -131.070 -82.950 ;
        RECT -127.350 -83.240 -127.030 -82.950 ;
        RECT -121.470 -83.240 -121.150 -82.950 ;
        RECT -117.430 -83.240 -117.110 -82.950 ;
        RECT -111.550 -83.240 -111.230 -82.950 ;
        RECT -107.510 -83.240 -107.190 -82.950 ;
        RECT -101.630 -83.240 -101.310 -82.950 ;
        RECT -97.590 -83.240 -97.270 -82.950 ;
        RECT -91.710 -83.240 -91.390 -82.950 ;
        RECT -87.670 -83.240 -87.350 -82.950 ;
        RECT -81.790 -83.240 -81.470 -82.950 ;
        RECT -77.750 -83.240 -77.430 -82.950 ;
        RECT -71.870 -83.240 -71.550 -82.950 ;
        RECT -67.830 -83.240 -67.510 -82.950 ;
        RECT -61.950 -83.240 -61.630 -82.950 ;
        RECT -57.910 -83.240 -57.590 -82.950 ;
        RECT -52.030 -83.240 -51.710 -82.950 ;
        RECT -47.990 -83.240 -47.670 -82.950 ;
        RECT -42.110 -83.240 -41.790 -82.950 ;
        RECT -38.070 -83.240 -37.750 -82.950 ;
        RECT -32.190 -83.240 -31.870 -82.950 ;
        RECT -28.150 -83.240 -27.830 -82.950 ;
        RECT -22.270 -83.240 -21.950 -82.950 ;
        RECT -18.230 -83.240 -17.910 -82.950 ;
        RECT -12.350 -83.240 -12.030 -82.950 ;
        RECT -8.310 -83.240 -7.990 -82.950 ;
        RECT -2.430 -83.240 -2.110 -82.950 ;
        RECT 1.610 -83.240 1.930 -82.950 ;
        RECT 7.490 -83.240 7.810 -82.950 ;
        RECT 11.530 -83.240 11.850 -82.950 ;
        RECT 17.410 -83.240 17.730 -82.950 ;
        RECT 21.450 -83.240 21.770 -82.950 ;
        RECT -291.820 -84.200 -290.880 -83.720 ;
        RECT 22.540 -83.720 23.020 -82.820 ;
        RECT -286.810 -84.120 -285.120 -83.820 ;
        RECT -276.890 -84.120 -275.200 -83.820 ;
        RECT -266.970 -84.120 -265.280 -83.820 ;
        RECT -257.050 -84.120 -255.360 -83.820 ;
        RECT -247.130 -84.120 -245.440 -83.820 ;
        RECT -237.210 -84.120 -235.520 -83.820 ;
        RECT -227.290 -84.120 -225.600 -83.820 ;
        RECT -217.370 -84.120 -215.680 -83.820 ;
        RECT -207.450 -84.120 -205.760 -83.820 ;
        RECT -197.530 -84.120 -195.840 -83.820 ;
        RECT -187.610 -84.120 -185.920 -83.820 ;
        RECT -177.690 -84.120 -176.000 -83.820 ;
        RECT -167.770 -84.120 -166.080 -83.820 ;
        RECT -157.850 -84.120 -156.160 -83.820 ;
        RECT -147.930 -84.120 -146.240 -83.820 ;
        RECT -138.010 -84.120 -136.320 -83.820 ;
        RECT -128.090 -84.120 -126.400 -83.820 ;
        RECT -118.170 -84.120 -116.480 -83.820 ;
        RECT -108.250 -84.120 -106.560 -83.820 ;
        RECT -98.330 -84.120 -96.640 -83.820 ;
        RECT -88.410 -84.120 -86.720 -83.820 ;
        RECT -78.490 -84.120 -76.800 -83.820 ;
        RECT -68.570 -84.120 -66.880 -83.820 ;
        RECT -58.650 -84.120 -56.960 -83.820 ;
        RECT -48.730 -84.120 -47.040 -83.820 ;
        RECT -38.810 -84.120 -37.120 -83.820 ;
        RECT -28.890 -84.120 -27.200 -83.820 ;
        RECT -18.970 -84.120 -17.280 -83.820 ;
        RECT -9.050 -84.120 -7.360 -83.820 ;
        RECT 0.870 -84.120 2.560 -83.820 ;
        RECT 10.790 -84.120 12.480 -83.820 ;
        RECT 20.710 -84.120 22.400 -83.820 ;
        RECT -286.300 -84.820 -285.300 -84.120 ;
        RECT -276.380 -84.820 -275.380 -84.120 ;
        RECT -266.460 -84.820 -265.460 -84.120 ;
        RECT -256.540 -84.820 -255.540 -84.120 ;
        RECT -246.620 -84.820 -245.620 -84.120 ;
        RECT -236.700 -84.820 -235.700 -84.120 ;
        RECT -226.780 -84.820 -225.780 -84.120 ;
        RECT -216.860 -84.820 -215.860 -84.120 ;
        RECT -206.940 -84.820 -205.940 -84.120 ;
        RECT -197.020 -84.820 -196.020 -84.120 ;
        RECT -187.100 -84.820 -186.100 -84.120 ;
        RECT -177.180 -84.820 -176.180 -84.120 ;
        RECT -167.260 -84.820 -166.260 -84.120 ;
        RECT -157.340 -84.820 -156.340 -84.120 ;
        RECT -147.420 -84.820 -146.420 -84.120 ;
        RECT -137.500 -84.820 -136.500 -84.120 ;
        RECT -127.580 -84.820 -126.580 -84.120 ;
        RECT -117.660 -84.820 -116.660 -84.120 ;
        RECT -107.740 -84.820 -106.740 -84.120 ;
        RECT -97.820 -84.820 -96.820 -84.120 ;
        RECT -87.900 -84.820 -86.900 -84.120 ;
        RECT -77.980 -84.820 -76.980 -84.120 ;
        RECT -68.060 -84.820 -67.060 -84.120 ;
        RECT -58.140 -84.820 -57.140 -84.120 ;
        RECT -48.220 -84.820 -47.220 -84.120 ;
        RECT -38.300 -84.820 -37.300 -84.120 ;
        RECT -28.380 -84.820 -27.380 -84.120 ;
        RECT -18.460 -84.820 -17.460 -84.120 ;
        RECT -8.540 -84.820 -7.540 -84.120 ;
        RECT 1.380 -84.820 2.380 -84.120 ;
        RECT 11.300 -84.820 12.300 -84.120 ;
        RECT 21.220 -84.820 22.220 -84.120 ;
        RECT 22.540 -84.200 23.480 -83.720 ;
        RECT -294.880 -172.440 -294.420 -172.435 ;
        RECT -294.880 -172.915 -293.940 -172.440 ;
        RECT -293.020 -172.520 -292.020 -171.820 ;
        RECT -283.100 -172.520 -282.100 -171.820 ;
        RECT -273.180 -172.520 -272.180 -171.820 ;
        RECT -263.260 -172.520 -262.260 -171.820 ;
        RECT -253.340 -172.520 -252.340 -171.820 ;
        RECT -243.420 -172.520 -242.420 -171.820 ;
        RECT -233.500 -172.520 -232.500 -171.820 ;
        RECT -223.580 -172.520 -222.580 -171.820 ;
        RECT -213.660 -172.520 -212.660 -171.820 ;
        RECT -203.740 -172.520 -202.740 -171.820 ;
        RECT -193.820 -172.520 -192.820 -171.820 ;
        RECT -183.900 -172.520 -182.900 -171.820 ;
        RECT -173.980 -172.520 -172.980 -171.820 ;
        RECT -164.060 -172.520 -163.060 -171.820 ;
        RECT -154.140 -172.520 -153.140 -171.820 ;
        RECT -144.220 -172.520 -143.220 -171.820 ;
        RECT -134.300 -172.520 -133.300 -171.820 ;
        RECT -124.380 -172.520 -123.380 -171.820 ;
        RECT -114.460 -172.520 -113.460 -171.820 ;
        RECT -104.540 -172.520 -103.540 -171.820 ;
        RECT -94.620 -172.520 -93.620 -171.820 ;
        RECT -84.700 -172.520 -83.700 -171.820 ;
        RECT -74.780 -172.520 -73.780 -171.820 ;
        RECT -64.860 -172.520 -63.860 -171.820 ;
        RECT -54.940 -172.520 -53.940 -171.820 ;
        RECT -45.020 -172.520 -44.020 -171.820 ;
        RECT -35.100 -172.520 -34.100 -171.820 ;
        RECT -25.180 -172.520 -24.180 -171.820 ;
        RECT -15.260 -172.520 -14.260 -171.820 ;
        RECT -5.340 -172.520 -4.340 -171.820 ;
        RECT 4.580 -172.520 5.580 -171.820 ;
        RECT 14.500 -172.520 15.500 -171.820 ;
        RECT -293.530 -172.820 -291.840 -172.520 ;
        RECT -283.610 -172.820 -281.920 -172.520 ;
        RECT -273.690 -172.820 -272.000 -172.520 ;
        RECT -263.770 -172.820 -262.080 -172.520 ;
        RECT -253.850 -172.820 -252.160 -172.520 ;
        RECT -243.930 -172.820 -242.240 -172.520 ;
        RECT -234.010 -172.820 -232.320 -172.520 ;
        RECT -224.090 -172.820 -222.400 -172.520 ;
        RECT -214.170 -172.820 -212.480 -172.520 ;
        RECT -204.250 -172.820 -202.560 -172.520 ;
        RECT -194.330 -172.820 -192.640 -172.520 ;
        RECT -184.410 -172.820 -182.720 -172.520 ;
        RECT -174.490 -172.820 -172.800 -172.520 ;
        RECT -164.570 -172.820 -162.880 -172.520 ;
        RECT -154.650 -172.820 -152.960 -172.520 ;
        RECT -144.730 -172.820 -143.040 -172.520 ;
        RECT -134.810 -172.820 -133.120 -172.520 ;
        RECT -124.890 -172.820 -123.200 -172.520 ;
        RECT -114.970 -172.820 -113.280 -172.520 ;
        RECT -105.050 -172.820 -103.360 -172.520 ;
        RECT -95.130 -172.820 -93.440 -172.520 ;
        RECT -85.210 -172.820 -83.520 -172.520 ;
        RECT -75.290 -172.820 -73.600 -172.520 ;
        RECT -65.370 -172.820 -63.680 -172.520 ;
        RECT -55.450 -172.820 -53.760 -172.520 ;
        RECT -45.530 -172.820 -43.840 -172.520 ;
        RECT -35.610 -172.820 -33.920 -172.520 ;
        RECT -25.690 -172.820 -24.000 -172.520 ;
        RECT -15.770 -172.820 -14.080 -172.520 ;
        RECT -5.850 -172.820 -4.160 -172.520 ;
        RECT 4.070 -172.820 5.760 -172.520 ;
        RECT 13.990 -172.820 15.680 -172.520 ;
        RECT -294.420 -173.820 -293.940 -172.915 ;
        RECT -292.790 -173.690 -292.470 -173.400 ;
        RECT -286.910 -173.690 -286.590 -173.400 ;
        RECT -282.870 -173.690 -282.550 -173.400 ;
        RECT -276.990 -173.690 -276.670 -173.400 ;
        RECT -272.950 -173.690 -272.630 -173.400 ;
        RECT -267.070 -173.690 -266.750 -173.400 ;
        RECT -263.030 -173.690 -262.710 -173.400 ;
        RECT -257.150 -173.690 -256.830 -173.400 ;
        RECT -253.110 -173.690 -252.790 -173.400 ;
        RECT -247.230 -173.690 -246.910 -173.400 ;
        RECT -243.190 -173.690 -242.870 -173.400 ;
        RECT -237.310 -173.690 -236.990 -173.400 ;
        RECT -233.270 -173.690 -232.950 -173.400 ;
        RECT -227.390 -173.690 -227.070 -173.400 ;
        RECT -223.350 -173.690 -223.030 -173.400 ;
        RECT -217.470 -173.690 -217.150 -173.400 ;
        RECT -213.430 -173.690 -213.110 -173.400 ;
        RECT -207.550 -173.690 -207.230 -173.400 ;
        RECT -203.510 -173.690 -203.190 -173.400 ;
        RECT -197.630 -173.690 -197.310 -173.400 ;
        RECT -193.590 -173.690 -193.270 -173.400 ;
        RECT -187.710 -173.690 -187.390 -173.400 ;
        RECT -183.670 -173.690 -183.350 -173.400 ;
        RECT -177.790 -173.690 -177.470 -173.400 ;
        RECT -173.750 -173.690 -173.430 -173.400 ;
        RECT -167.870 -173.690 -167.550 -173.400 ;
        RECT -163.830 -173.690 -163.510 -173.400 ;
        RECT -157.950 -173.690 -157.630 -173.400 ;
        RECT -153.910 -173.690 -153.590 -173.400 ;
        RECT -148.030 -173.690 -147.710 -173.400 ;
        RECT -143.990 -173.690 -143.670 -173.400 ;
        RECT -138.110 -173.690 -137.790 -173.400 ;
        RECT -134.070 -173.690 -133.750 -173.400 ;
        RECT -128.190 -173.690 -127.870 -173.400 ;
        RECT -124.150 -173.690 -123.830 -173.400 ;
        RECT -118.270 -173.690 -117.950 -173.400 ;
        RECT -114.230 -173.690 -113.910 -173.400 ;
        RECT -108.350 -173.690 -108.030 -173.400 ;
        RECT -104.310 -173.690 -103.990 -173.400 ;
        RECT -98.430 -173.690 -98.110 -173.400 ;
        RECT -94.390 -173.690 -94.070 -173.400 ;
        RECT -88.510 -173.690 -88.190 -173.400 ;
        RECT -84.470 -173.690 -84.150 -173.400 ;
        RECT -78.590 -173.690 -78.270 -173.400 ;
        RECT -74.550 -173.690 -74.230 -173.400 ;
        RECT -68.670 -173.690 -68.350 -173.400 ;
        RECT -64.630 -173.690 -64.310 -173.400 ;
        RECT -58.750 -173.690 -58.430 -173.400 ;
        RECT -54.710 -173.690 -54.390 -173.400 ;
        RECT -48.830 -173.690 -48.510 -173.400 ;
        RECT -44.790 -173.690 -44.470 -173.400 ;
        RECT -38.910 -173.690 -38.590 -173.400 ;
        RECT -34.870 -173.690 -34.550 -173.400 ;
        RECT -28.990 -173.690 -28.670 -173.400 ;
        RECT -24.950 -173.690 -24.630 -173.400 ;
        RECT -19.070 -173.690 -18.750 -173.400 ;
        RECT -15.030 -173.690 -14.710 -173.400 ;
        RECT -9.150 -173.690 -8.830 -173.400 ;
        RECT -5.110 -173.690 -4.790 -173.400 ;
        RECT 0.770 -173.690 1.090 -173.400 ;
        RECT 4.810 -173.690 5.130 -173.400 ;
        RECT 10.690 -173.690 11.010 -173.400 ;
        RECT 14.730 -173.690 15.050 -173.400 ;
        RECT 20.610 -173.690 20.930 -173.400 ;
        RECT -294.880 -174.490 -293.040 -174.010 ;
        RECT -292.710 -174.820 -292.520 -173.690 ;
        RECT -286.860 -174.820 -286.670 -173.690 ;
        RECT -282.790 -174.820 -282.600 -173.690 ;
        RECT -276.940 -174.820 -276.750 -173.690 ;
        RECT -272.870 -174.820 -272.680 -173.690 ;
        RECT -267.020 -174.820 -266.830 -173.690 ;
        RECT -262.950 -174.820 -262.760 -173.690 ;
        RECT -257.100 -174.820 -256.910 -173.690 ;
        RECT -253.030 -174.820 -252.840 -173.690 ;
        RECT -247.180 -174.820 -246.990 -173.690 ;
        RECT -243.110 -174.820 -242.920 -173.690 ;
        RECT -237.260 -174.820 -237.070 -173.690 ;
        RECT -233.190 -174.820 -233.000 -173.690 ;
        RECT -227.340 -174.820 -227.150 -173.690 ;
        RECT -223.270 -174.820 -223.080 -173.690 ;
        RECT -217.420 -174.820 -217.230 -173.690 ;
        RECT -213.350 -174.820 -213.160 -173.690 ;
        RECT -207.500 -174.820 -207.310 -173.690 ;
        RECT -203.430 -174.820 -203.240 -173.690 ;
        RECT -197.580 -174.820 -197.390 -173.690 ;
        RECT -193.510 -174.820 -193.320 -173.690 ;
        RECT -187.660 -174.820 -187.470 -173.690 ;
        RECT -183.590 -174.820 -183.400 -173.690 ;
        RECT -177.740 -174.820 -177.550 -173.690 ;
        RECT -173.670 -174.820 -173.480 -173.690 ;
        RECT -167.820 -174.820 -167.630 -173.690 ;
        RECT -163.750 -174.820 -163.560 -173.690 ;
        RECT -157.900 -174.820 -157.710 -173.690 ;
        RECT -153.830 -174.820 -153.640 -173.690 ;
        RECT -147.980 -174.820 -147.790 -173.690 ;
        RECT -143.910 -174.820 -143.720 -173.690 ;
        RECT -138.060 -174.820 -137.870 -173.690 ;
        RECT -133.990 -174.820 -133.800 -173.690 ;
        RECT -128.140 -174.820 -127.950 -173.690 ;
        RECT -124.070 -174.820 -123.880 -173.690 ;
        RECT -118.220 -174.820 -118.030 -173.690 ;
        RECT -114.150 -174.820 -113.960 -173.690 ;
        RECT -108.300 -174.820 -108.110 -173.690 ;
        RECT -104.230 -174.820 -104.040 -173.690 ;
        RECT -98.380 -174.820 -98.190 -173.690 ;
        RECT -94.310 -174.820 -94.120 -173.690 ;
        RECT -88.460 -174.820 -88.270 -173.690 ;
        RECT -84.390 -174.820 -84.200 -173.690 ;
        RECT -78.540 -174.820 -78.350 -173.690 ;
        RECT -74.470 -174.820 -74.280 -173.690 ;
        RECT -68.620 -174.820 -68.430 -173.690 ;
        RECT -64.550 -174.820 -64.360 -173.690 ;
        RECT -58.700 -174.820 -58.510 -173.690 ;
        RECT -54.630 -174.820 -54.440 -173.690 ;
        RECT -48.780 -174.820 -48.590 -173.690 ;
        RECT -44.710 -174.820 -44.520 -173.690 ;
        RECT -38.860 -174.820 -38.670 -173.690 ;
        RECT -34.790 -174.820 -34.600 -173.690 ;
        RECT -28.940 -174.820 -28.750 -173.690 ;
        RECT -24.870 -174.820 -24.680 -173.690 ;
        RECT -19.020 -174.820 -18.830 -173.690 ;
        RECT -14.950 -174.820 -14.760 -173.690 ;
        RECT -9.100 -174.820 -8.910 -173.690 ;
        RECT -5.030 -174.820 -4.840 -173.690 ;
        RECT 0.820 -174.820 1.010 -173.690 ;
        RECT 4.890 -174.820 5.080 -173.690 ;
        RECT 10.740 -174.820 10.930 -173.690 ;
        RECT 14.810 -174.820 15.000 -173.690 ;
        RECT 20.660 -174.820 20.850 -173.690 ;
        RECT 21.180 -174.490 23.020 -174.010 ;
        RECT -293.470 -174.970 -291.530 -174.820 ;
        RECT -293.470 -175.120 -293.130 -174.970 ;
        RECT -293.470 -175.320 -293.150 -175.290 ;
        RECT -293.470 -175.460 -292.650 -175.320 ;
        RECT -293.470 -175.570 -293.150 -175.460 ;
        RECT -292.810 -176.250 -292.650 -175.460 ;
        RECT -291.690 -175.760 -291.530 -174.970 ;
        RECT -287.850 -174.970 -285.910 -174.820 ;
        RECT -291.190 -175.760 -290.870 -175.650 ;
        RECT -291.690 -175.900 -290.870 -175.760 ;
        RECT -291.190 -175.930 -290.870 -175.900 ;
        RECT -288.510 -175.760 -288.190 -175.650 ;
        RECT -287.850 -175.760 -287.690 -174.970 ;
        RECT -286.250 -175.120 -285.910 -174.970 ;
        RECT -283.550 -174.970 -281.610 -174.820 ;
        RECT -283.550 -175.120 -283.210 -174.970 ;
        RECT -286.230 -175.320 -285.910 -175.290 ;
        RECT -288.510 -175.900 -287.690 -175.760 ;
        RECT -286.730 -175.460 -285.910 -175.320 ;
        RECT -288.510 -175.930 -288.190 -175.900 ;
        RECT -291.210 -176.250 -290.870 -176.100 ;
        RECT -292.810 -176.400 -290.870 -176.250 ;
        RECT -288.510 -176.250 -288.170 -176.100 ;
        RECT -286.730 -176.250 -286.570 -175.460 ;
        RECT -286.230 -175.570 -285.910 -175.460 ;
        RECT -283.550 -175.320 -283.230 -175.290 ;
        RECT -283.550 -175.460 -282.730 -175.320 ;
        RECT -283.550 -175.570 -283.230 -175.460 ;
        RECT -288.510 -176.400 -286.570 -176.250 ;
        RECT -282.890 -176.250 -282.730 -175.460 ;
        RECT -281.770 -175.760 -281.610 -174.970 ;
        RECT -277.930 -174.970 -275.990 -174.820 ;
        RECT -281.270 -175.760 -280.950 -175.650 ;
        RECT -281.770 -175.900 -280.950 -175.760 ;
        RECT -281.270 -175.930 -280.950 -175.900 ;
        RECT -278.590 -175.760 -278.270 -175.650 ;
        RECT -277.930 -175.760 -277.770 -174.970 ;
        RECT -276.330 -175.120 -275.990 -174.970 ;
        RECT -273.630 -174.970 -271.690 -174.820 ;
        RECT -273.630 -175.120 -273.290 -174.970 ;
        RECT -276.310 -175.320 -275.990 -175.290 ;
        RECT -278.590 -175.900 -277.770 -175.760 ;
        RECT -276.810 -175.460 -275.990 -175.320 ;
        RECT -278.590 -175.930 -278.270 -175.900 ;
        RECT -281.290 -176.250 -280.950 -176.100 ;
        RECT -282.890 -176.400 -280.950 -176.250 ;
        RECT -278.590 -176.250 -278.250 -176.100 ;
        RECT -276.810 -176.250 -276.650 -175.460 ;
        RECT -276.310 -175.570 -275.990 -175.460 ;
        RECT -273.630 -175.320 -273.310 -175.290 ;
        RECT -273.630 -175.460 -272.810 -175.320 ;
        RECT -273.630 -175.570 -273.310 -175.460 ;
        RECT -278.590 -176.400 -276.650 -176.250 ;
        RECT -272.970 -176.250 -272.810 -175.460 ;
        RECT -271.850 -175.760 -271.690 -174.970 ;
        RECT -268.010 -174.970 -266.070 -174.820 ;
        RECT -271.350 -175.760 -271.030 -175.650 ;
        RECT -271.850 -175.900 -271.030 -175.760 ;
        RECT -271.350 -175.930 -271.030 -175.900 ;
        RECT -268.670 -175.760 -268.350 -175.650 ;
        RECT -268.010 -175.760 -267.850 -174.970 ;
        RECT -266.410 -175.120 -266.070 -174.970 ;
        RECT -263.710 -174.970 -261.770 -174.820 ;
        RECT -263.710 -175.120 -263.370 -174.970 ;
        RECT -266.390 -175.320 -266.070 -175.290 ;
        RECT -268.670 -175.900 -267.850 -175.760 ;
        RECT -266.890 -175.460 -266.070 -175.320 ;
        RECT -268.670 -175.930 -268.350 -175.900 ;
        RECT -271.370 -176.250 -271.030 -176.100 ;
        RECT -272.970 -176.400 -271.030 -176.250 ;
        RECT -268.670 -176.250 -268.330 -176.100 ;
        RECT -266.890 -176.250 -266.730 -175.460 ;
        RECT -266.390 -175.570 -266.070 -175.460 ;
        RECT -263.710 -175.320 -263.390 -175.290 ;
        RECT -263.710 -175.460 -262.890 -175.320 ;
        RECT -263.710 -175.570 -263.390 -175.460 ;
        RECT -268.670 -176.400 -266.730 -176.250 ;
        RECT -263.050 -176.250 -262.890 -175.460 ;
        RECT -261.930 -175.760 -261.770 -174.970 ;
        RECT -258.090 -174.970 -256.150 -174.820 ;
        RECT -261.430 -175.760 -261.110 -175.650 ;
        RECT -261.930 -175.900 -261.110 -175.760 ;
        RECT -261.430 -175.930 -261.110 -175.900 ;
        RECT -258.750 -175.760 -258.430 -175.650 ;
        RECT -258.090 -175.760 -257.930 -174.970 ;
        RECT -256.490 -175.120 -256.150 -174.970 ;
        RECT -253.790 -174.970 -251.850 -174.820 ;
        RECT -253.790 -175.120 -253.450 -174.970 ;
        RECT -256.470 -175.320 -256.150 -175.290 ;
        RECT -258.750 -175.900 -257.930 -175.760 ;
        RECT -256.970 -175.460 -256.150 -175.320 ;
        RECT -258.750 -175.930 -258.430 -175.900 ;
        RECT -261.450 -176.250 -261.110 -176.100 ;
        RECT -263.050 -176.400 -261.110 -176.250 ;
        RECT -258.750 -176.250 -258.410 -176.100 ;
        RECT -256.970 -176.250 -256.810 -175.460 ;
        RECT -256.470 -175.570 -256.150 -175.460 ;
        RECT -253.790 -175.320 -253.470 -175.290 ;
        RECT -253.790 -175.460 -252.970 -175.320 ;
        RECT -253.790 -175.570 -253.470 -175.460 ;
        RECT -258.750 -176.400 -256.810 -176.250 ;
        RECT -253.130 -176.250 -252.970 -175.460 ;
        RECT -252.010 -175.760 -251.850 -174.970 ;
        RECT -248.170 -174.970 -246.230 -174.820 ;
        RECT -251.510 -175.760 -251.190 -175.650 ;
        RECT -252.010 -175.900 -251.190 -175.760 ;
        RECT -251.510 -175.930 -251.190 -175.900 ;
        RECT -248.830 -175.760 -248.510 -175.650 ;
        RECT -248.170 -175.760 -248.010 -174.970 ;
        RECT -246.570 -175.120 -246.230 -174.970 ;
        RECT -243.870 -174.970 -241.930 -174.820 ;
        RECT -243.870 -175.120 -243.530 -174.970 ;
        RECT -246.550 -175.320 -246.230 -175.290 ;
        RECT -248.830 -175.900 -248.010 -175.760 ;
        RECT -247.050 -175.460 -246.230 -175.320 ;
        RECT -248.830 -175.930 -248.510 -175.900 ;
        RECT -251.530 -176.250 -251.190 -176.100 ;
        RECT -253.130 -176.400 -251.190 -176.250 ;
        RECT -248.830 -176.250 -248.490 -176.100 ;
        RECT -247.050 -176.250 -246.890 -175.460 ;
        RECT -246.550 -175.570 -246.230 -175.460 ;
        RECT -243.870 -175.320 -243.550 -175.290 ;
        RECT -243.870 -175.460 -243.050 -175.320 ;
        RECT -243.870 -175.570 -243.550 -175.460 ;
        RECT -248.830 -176.400 -246.890 -176.250 ;
        RECT -243.210 -176.250 -243.050 -175.460 ;
        RECT -242.090 -175.760 -241.930 -174.970 ;
        RECT -238.250 -174.970 -236.310 -174.820 ;
        RECT -241.590 -175.760 -241.270 -175.650 ;
        RECT -242.090 -175.900 -241.270 -175.760 ;
        RECT -241.590 -175.930 -241.270 -175.900 ;
        RECT -238.910 -175.760 -238.590 -175.650 ;
        RECT -238.250 -175.760 -238.090 -174.970 ;
        RECT -236.650 -175.120 -236.310 -174.970 ;
        RECT -233.950 -174.970 -232.010 -174.820 ;
        RECT -233.950 -175.120 -233.610 -174.970 ;
        RECT -236.630 -175.320 -236.310 -175.290 ;
        RECT -238.910 -175.900 -238.090 -175.760 ;
        RECT -237.130 -175.460 -236.310 -175.320 ;
        RECT -238.910 -175.930 -238.590 -175.900 ;
        RECT -241.610 -176.250 -241.270 -176.100 ;
        RECT -243.210 -176.400 -241.270 -176.250 ;
        RECT -238.910 -176.250 -238.570 -176.100 ;
        RECT -237.130 -176.250 -236.970 -175.460 ;
        RECT -236.630 -175.570 -236.310 -175.460 ;
        RECT -233.950 -175.320 -233.630 -175.290 ;
        RECT -233.950 -175.460 -233.130 -175.320 ;
        RECT -233.950 -175.570 -233.630 -175.460 ;
        RECT -238.910 -176.400 -236.970 -176.250 ;
        RECT -233.290 -176.250 -233.130 -175.460 ;
        RECT -232.170 -175.760 -232.010 -174.970 ;
        RECT -228.330 -174.970 -226.390 -174.820 ;
        RECT -231.670 -175.760 -231.350 -175.650 ;
        RECT -232.170 -175.900 -231.350 -175.760 ;
        RECT -231.670 -175.930 -231.350 -175.900 ;
        RECT -228.990 -175.760 -228.670 -175.650 ;
        RECT -228.330 -175.760 -228.170 -174.970 ;
        RECT -226.730 -175.120 -226.390 -174.970 ;
        RECT -224.030 -174.970 -222.090 -174.820 ;
        RECT -224.030 -175.120 -223.690 -174.970 ;
        RECT -226.710 -175.320 -226.390 -175.290 ;
        RECT -228.990 -175.900 -228.170 -175.760 ;
        RECT -227.210 -175.460 -226.390 -175.320 ;
        RECT -228.990 -175.930 -228.670 -175.900 ;
        RECT -231.690 -176.250 -231.350 -176.100 ;
        RECT -233.290 -176.400 -231.350 -176.250 ;
        RECT -228.990 -176.250 -228.650 -176.100 ;
        RECT -227.210 -176.250 -227.050 -175.460 ;
        RECT -226.710 -175.570 -226.390 -175.460 ;
        RECT -224.030 -175.320 -223.710 -175.290 ;
        RECT -224.030 -175.460 -223.210 -175.320 ;
        RECT -224.030 -175.570 -223.710 -175.460 ;
        RECT -228.990 -176.400 -227.050 -176.250 ;
        RECT -223.370 -176.250 -223.210 -175.460 ;
        RECT -222.250 -175.760 -222.090 -174.970 ;
        RECT -218.410 -174.970 -216.470 -174.820 ;
        RECT -221.750 -175.760 -221.430 -175.650 ;
        RECT -222.250 -175.900 -221.430 -175.760 ;
        RECT -221.750 -175.930 -221.430 -175.900 ;
        RECT -219.070 -175.760 -218.750 -175.650 ;
        RECT -218.410 -175.760 -218.250 -174.970 ;
        RECT -216.810 -175.120 -216.470 -174.970 ;
        RECT -214.110 -174.970 -212.170 -174.820 ;
        RECT -214.110 -175.120 -213.770 -174.970 ;
        RECT -216.790 -175.320 -216.470 -175.290 ;
        RECT -219.070 -175.900 -218.250 -175.760 ;
        RECT -217.290 -175.460 -216.470 -175.320 ;
        RECT -219.070 -175.930 -218.750 -175.900 ;
        RECT -221.770 -176.250 -221.430 -176.100 ;
        RECT -223.370 -176.400 -221.430 -176.250 ;
        RECT -219.070 -176.250 -218.730 -176.100 ;
        RECT -217.290 -176.250 -217.130 -175.460 ;
        RECT -216.790 -175.570 -216.470 -175.460 ;
        RECT -214.110 -175.320 -213.790 -175.290 ;
        RECT -214.110 -175.460 -213.290 -175.320 ;
        RECT -214.110 -175.570 -213.790 -175.460 ;
        RECT -219.070 -176.400 -217.130 -176.250 ;
        RECT -213.450 -176.250 -213.290 -175.460 ;
        RECT -212.330 -175.760 -212.170 -174.970 ;
        RECT -208.490 -174.970 -206.550 -174.820 ;
        RECT -211.830 -175.760 -211.510 -175.650 ;
        RECT -212.330 -175.900 -211.510 -175.760 ;
        RECT -211.830 -175.930 -211.510 -175.900 ;
        RECT -209.150 -175.760 -208.830 -175.650 ;
        RECT -208.490 -175.760 -208.330 -174.970 ;
        RECT -206.890 -175.120 -206.550 -174.970 ;
        RECT -204.190 -174.970 -202.250 -174.820 ;
        RECT -204.190 -175.120 -203.850 -174.970 ;
        RECT -206.870 -175.320 -206.550 -175.290 ;
        RECT -209.150 -175.900 -208.330 -175.760 ;
        RECT -207.370 -175.460 -206.550 -175.320 ;
        RECT -209.150 -175.930 -208.830 -175.900 ;
        RECT -211.850 -176.250 -211.510 -176.100 ;
        RECT -213.450 -176.400 -211.510 -176.250 ;
        RECT -209.150 -176.250 -208.810 -176.100 ;
        RECT -207.370 -176.250 -207.210 -175.460 ;
        RECT -206.870 -175.570 -206.550 -175.460 ;
        RECT -204.190 -175.320 -203.870 -175.290 ;
        RECT -204.190 -175.460 -203.370 -175.320 ;
        RECT -204.190 -175.570 -203.870 -175.460 ;
        RECT -209.150 -176.400 -207.210 -176.250 ;
        RECT -203.530 -176.250 -203.370 -175.460 ;
        RECT -202.410 -175.760 -202.250 -174.970 ;
        RECT -198.570 -174.970 -196.630 -174.820 ;
        RECT -201.910 -175.760 -201.590 -175.650 ;
        RECT -202.410 -175.900 -201.590 -175.760 ;
        RECT -201.910 -175.930 -201.590 -175.900 ;
        RECT -199.230 -175.760 -198.910 -175.650 ;
        RECT -198.570 -175.760 -198.410 -174.970 ;
        RECT -196.970 -175.120 -196.630 -174.970 ;
        RECT -194.270 -174.970 -192.330 -174.820 ;
        RECT -194.270 -175.120 -193.930 -174.970 ;
        RECT -196.950 -175.320 -196.630 -175.290 ;
        RECT -199.230 -175.900 -198.410 -175.760 ;
        RECT -197.450 -175.460 -196.630 -175.320 ;
        RECT -199.230 -175.930 -198.910 -175.900 ;
        RECT -201.930 -176.250 -201.590 -176.100 ;
        RECT -203.530 -176.400 -201.590 -176.250 ;
        RECT -199.230 -176.250 -198.890 -176.100 ;
        RECT -197.450 -176.250 -197.290 -175.460 ;
        RECT -196.950 -175.570 -196.630 -175.460 ;
        RECT -194.270 -175.320 -193.950 -175.290 ;
        RECT -194.270 -175.460 -193.450 -175.320 ;
        RECT -194.270 -175.570 -193.950 -175.460 ;
        RECT -199.230 -176.400 -197.290 -176.250 ;
        RECT -193.610 -176.250 -193.450 -175.460 ;
        RECT -192.490 -175.760 -192.330 -174.970 ;
        RECT -188.650 -174.970 -186.710 -174.820 ;
        RECT -191.990 -175.760 -191.670 -175.650 ;
        RECT -192.490 -175.900 -191.670 -175.760 ;
        RECT -191.990 -175.930 -191.670 -175.900 ;
        RECT -189.310 -175.760 -188.990 -175.650 ;
        RECT -188.650 -175.760 -188.490 -174.970 ;
        RECT -187.050 -175.120 -186.710 -174.970 ;
        RECT -184.350 -174.970 -182.410 -174.820 ;
        RECT -184.350 -175.120 -184.010 -174.970 ;
        RECT -187.030 -175.320 -186.710 -175.290 ;
        RECT -189.310 -175.900 -188.490 -175.760 ;
        RECT -187.530 -175.460 -186.710 -175.320 ;
        RECT -189.310 -175.930 -188.990 -175.900 ;
        RECT -192.010 -176.250 -191.670 -176.100 ;
        RECT -193.610 -176.400 -191.670 -176.250 ;
        RECT -189.310 -176.250 -188.970 -176.100 ;
        RECT -187.530 -176.250 -187.370 -175.460 ;
        RECT -187.030 -175.570 -186.710 -175.460 ;
        RECT -184.350 -175.320 -184.030 -175.290 ;
        RECT -184.350 -175.460 -183.530 -175.320 ;
        RECT -184.350 -175.570 -184.030 -175.460 ;
        RECT -189.310 -176.400 -187.370 -176.250 ;
        RECT -183.690 -176.250 -183.530 -175.460 ;
        RECT -182.570 -175.760 -182.410 -174.970 ;
        RECT -178.730 -174.970 -176.790 -174.820 ;
        RECT -182.070 -175.760 -181.750 -175.650 ;
        RECT -182.570 -175.900 -181.750 -175.760 ;
        RECT -182.070 -175.930 -181.750 -175.900 ;
        RECT -179.390 -175.760 -179.070 -175.650 ;
        RECT -178.730 -175.760 -178.570 -174.970 ;
        RECT -177.130 -175.120 -176.790 -174.970 ;
        RECT -174.430 -174.970 -172.490 -174.820 ;
        RECT -174.430 -175.120 -174.090 -174.970 ;
        RECT -177.110 -175.320 -176.790 -175.290 ;
        RECT -179.390 -175.900 -178.570 -175.760 ;
        RECT -177.610 -175.460 -176.790 -175.320 ;
        RECT -179.390 -175.930 -179.070 -175.900 ;
        RECT -182.090 -176.250 -181.750 -176.100 ;
        RECT -183.690 -176.400 -181.750 -176.250 ;
        RECT -179.390 -176.250 -179.050 -176.100 ;
        RECT -177.610 -176.250 -177.450 -175.460 ;
        RECT -177.110 -175.570 -176.790 -175.460 ;
        RECT -174.430 -175.320 -174.110 -175.290 ;
        RECT -174.430 -175.460 -173.610 -175.320 ;
        RECT -174.430 -175.570 -174.110 -175.460 ;
        RECT -179.390 -176.400 -177.450 -176.250 ;
        RECT -173.770 -176.250 -173.610 -175.460 ;
        RECT -172.650 -175.760 -172.490 -174.970 ;
        RECT -168.810 -174.970 -166.870 -174.820 ;
        RECT -172.150 -175.760 -171.830 -175.650 ;
        RECT -172.650 -175.900 -171.830 -175.760 ;
        RECT -172.150 -175.930 -171.830 -175.900 ;
        RECT -169.470 -175.760 -169.150 -175.650 ;
        RECT -168.810 -175.760 -168.650 -174.970 ;
        RECT -167.210 -175.120 -166.870 -174.970 ;
        RECT -164.510 -174.970 -162.570 -174.820 ;
        RECT -164.510 -175.120 -164.170 -174.970 ;
        RECT -167.190 -175.320 -166.870 -175.290 ;
        RECT -169.470 -175.900 -168.650 -175.760 ;
        RECT -167.690 -175.460 -166.870 -175.320 ;
        RECT -169.470 -175.930 -169.150 -175.900 ;
        RECT -172.170 -176.250 -171.830 -176.100 ;
        RECT -173.770 -176.400 -171.830 -176.250 ;
        RECT -169.470 -176.250 -169.130 -176.100 ;
        RECT -167.690 -176.250 -167.530 -175.460 ;
        RECT -167.190 -175.570 -166.870 -175.460 ;
        RECT -164.510 -175.320 -164.190 -175.290 ;
        RECT -164.510 -175.460 -163.690 -175.320 ;
        RECT -164.510 -175.570 -164.190 -175.460 ;
        RECT -169.470 -176.400 -167.530 -176.250 ;
        RECT -163.850 -176.250 -163.690 -175.460 ;
        RECT -162.730 -175.760 -162.570 -174.970 ;
        RECT -158.890 -174.970 -156.950 -174.820 ;
        RECT -162.230 -175.760 -161.910 -175.650 ;
        RECT -162.730 -175.900 -161.910 -175.760 ;
        RECT -162.230 -175.930 -161.910 -175.900 ;
        RECT -159.550 -175.760 -159.230 -175.650 ;
        RECT -158.890 -175.760 -158.730 -174.970 ;
        RECT -157.290 -175.120 -156.950 -174.970 ;
        RECT -154.590 -174.970 -152.650 -174.820 ;
        RECT -154.590 -175.120 -154.250 -174.970 ;
        RECT -157.270 -175.320 -156.950 -175.290 ;
        RECT -159.550 -175.900 -158.730 -175.760 ;
        RECT -157.770 -175.460 -156.950 -175.320 ;
        RECT -159.550 -175.930 -159.230 -175.900 ;
        RECT -162.250 -176.250 -161.910 -176.100 ;
        RECT -163.850 -176.400 -161.910 -176.250 ;
        RECT -159.550 -176.250 -159.210 -176.100 ;
        RECT -157.770 -176.250 -157.610 -175.460 ;
        RECT -157.270 -175.570 -156.950 -175.460 ;
        RECT -154.590 -175.320 -154.270 -175.290 ;
        RECT -154.590 -175.460 -153.770 -175.320 ;
        RECT -154.590 -175.570 -154.270 -175.460 ;
        RECT -159.550 -176.400 -157.610 -176.250 ;
        RECT -153.930 -176.250 -153.770 -175.460 ;
        RECT -152.810 -175.760 -152.650 -174.970 ;
        RECT -148.970 -174.970 -147.030 -174.820 ;
        RECT -152.310 -175.760 -151.990 -175.650 ;
        RECT -152.810 -175.900 -151.990 -175.760 ;
        RECT -152.310 -175.930 -151.990 -175.900 ;
        RECT -149.630 -175.760 -149.310 -175.650 ;
        RECT -148.970 -175.760 -148.810 -174.970 ;
        RECT -147.370 -175.120 -147.030 -174.970 ;
        RECT -144.670 -174.970 -142.730 -174.820 ;
        RECT -144.670 -175.120 -144.330 -174.970 ;
        RECT -147.350 -175.320 -147.030 -175.290 ;
        RECT -149.630 -175.900 -148.810 -175.760 ;
        RECT -147.850 -175.460 -147.030 -175.320 ;
        RECT -149.630 -175.930 -149.310 -175.900 ;
        RECT -152.330 -176.250 -151.990 -176.100 ;
        RECT -153.930 -176.400 -151.990 -176.250 ;
        RECT -149.630 -176.250 -149.290 -176.100 ;
        RECT -147.850 -176.250 -147.690 -175.460 ;
        RECT -147.350 -175.570 -147.030 -175.460 ;
        RECT -144.670 -175.320 -144.350 -175.290 ;
        RECT -144.670 -175.460 -143.850 -175.320 ;
        RECT -144.670 -175.570 -144.350 -175.460 ;
        RECT -149.630 -176.400 -147.690 -176.250 ;
        RECT -144.010 -176.250 -143.850 -175.460 ;
        RECT -142.890 -175.760 -142.730 -174.970 ;
        RECT -139.050 -174.970 -137.110 -174.820 ;
        RECT -142.390 -175.760 -142.070 -175.650 ;
        RECT -142.890 -175.900 -142.070 -175.760 ;
        RECT -142.390 -175.930 -142.070 -175.900 ;
        RECT -139.710 -175.760 -139.390 -175.650 ;
        RECT -139.050 -175.760 -138.890 -174.970 ;
        RECT -137.450 -175.120 -137.110 -174.970 ;
        RECT -134.750 -174.970 -132.810 -174.820 ;
        RECT -134.750 -175.120 -134.410 -174.970 ;
        RECT -137.430 -175.320 -137.110 -175.290 ;
        RECT -139.710 -175.900 -138.890 -175.760 ;
        RECT -137.930 -175.460 -137.110 -175.320 ;
        RECT -139.710 -175.930 -139.390 -175.900 ;
        RECT -142.410 -176.250 -142.070 -176.100 ;
        RECT -144.010 -176.400 -142.070 -176.250 ;
        RECT -139.710 -176.250 -139.370 -176.100 ;
        RECT -137.930 -176.250 -137.770 -175.460 ;
        RECT -137.430 -175.570 -137.110 -175.460 ;
        RECT -134.750 -175.320 -134.430 -175.290 ;
        RECT -134.750 -175.460 -133.930 -175.320 ;
        RECT -134.750 -175.570 -134.430 -175.460 ;
        RECT -139.710 -176.400 -137.770 -176.250 ;
        RECT -134.090 -176.250 -133.930 -175.460 ;
        RECT -132.970 -175.760 -132.810 -174.970 ;
        RECT -129.130 -174.970 -127.190 -174.820 ;
        RECT -132.470 -175.760 -132.150 -175.650 ;
        RECT -132.970 -175.900 -132.150 -175.760 ;
        RECT -132.470 -175.930 -132.150 -175.900 ;
        RECT -129.790 -175.760 -129.470 -175.650 ;
        RECT -129.130 -175.760 -128.970 -174.970 ;
        RECT -127.530 -175.120 -127.190 -174.970 ;
        RECT -124.830 -174.970 -122.890 -174.820 ;
        RECT -124.830 -175.120 -124.490 -174.970 ;
        RECT -127.510 -175.320 -127.190 -175.290 ;
        RECT -129.790 -175.900 -128.970 -175.760 ;
        RECT -128.010 -175.460 -127.190 -175.320 ;
        RECT -129.790 -175.930 -129.470 -175.900 ;
        RECT -132.490 -176.250 -132.150 -176.100 ;
        RECT -134.090 -176.400 -132.150 -176.250 ;
        RECT -129.790 -176.250 -129.450 -176.100 ;
        RECT -128.010 -176.250 -127.850 -175.460 ;
        RECT -127.510 -175.570 -127.190 -175.460 ;
        RECT -124.830 -175.320 -124.510 -175.290 ;
        RECT -124.830 -175.460 -124.010 -175.320 ;
        RECT -124.830 -175.570 -124.510 -175.460 ;
        RECT -129.790 -176.400 -127.850 -176.250 ;
        RECT -124.170 -176.250 -124.010 -175.460 ;
        RECT -123.050 -175.760 -122.890 -174.970 ;
        RECT -119.210 -174.970 -117.270 -174.820 ;
        RECT -122.550 -175.760 -122.230 -175.650 ;
        RECT -123.050 -175.900 -122.230 -175.760 ;
        RECT -122.550 -175.930 -122.230 -175.900 ;
        RECT -119.870 -175.760 -119.550 -175.650 ;
        RECT -119.210 -175.760 -119.050 -174.970 ;
        RECT -117.610 -175.120 -117.270 -174.970 ;
        RECT -114.910 -174.970 -112.970 -174.820 ;
        RECT -114.910 -175.120 -114.570 -174.970 ;
        RECT -117.590 -175.320 -117.270 -175.290 ;
        RECT -119.870 -175.900 -119.050 -175.760 ;
        RECT -118.090 -175.460 -117.270 -175.320 ;
        RECT -119.870 -175.930 -119.550 -175.900 ;
        RECT -122.570 -176.250 -122.230 -176.100 ;
        RECT -124.170 -176.400 -122.230 -176.250 ;
        RECT -119.870 -176.250 -119.530 -176.100 ;
        RECT -118.090 -176.250 -117.930 -175.460 ;
        RECT -117.590 -175.570 -117.270 -175.460 ;
        RECT -114.910 -175.320 -114.590 -175.290 ;
        RECT -114.910 -175.460 -114.090 -175.320 ;
        RECT -114.910 -175.570 -114.590 -175.460 ;
        RECT -119.870 -176.400 -117.930 -176.250 ;
        RECT -114.250 -176.250 -114.090 -175.460 ;
        RECT -113.130 -175.760 -112.970 -174.970 ;
        RECT -109.290 -174.970 -107.350 -174.820 ;
        RECT -112.630 -175.760 -112.310 -175.650 ;
        RECT -113.130 -175.900 -112.310 -175.760 ;
        RECT -112.630 -175.930 -112.310 -175.900 ;
        RECT -109.950 -175.760 -109.630 -175.650 ;
        RECT -109.290 -175.760 -109.130 -174.970 ;
        RECT -107.690 -175.120 -107.350 -174.970 ;
        RECT -104.990 -174.970 -103.050 -174.820 ;
        RECT -104.990 -175.120 -104.650 -174.970 ;
        RECT -107.670 -175.320 -107.350 -175.290 ;
        RECT -109.950 -175.900 -109.130 -175.760 ;
        RECT -108.170 -175.460 -107.350 -175.320 ;
        RECT -109.950 -175.930 -109.630 -175.900 ;
        RECT -112.650 -176.250 -112.310 -176.100 ;
        RECT -114.250 -176.400 -112.310 -176.250 ;
        RECT -109.950 -176.250 -109.610 -176.100 ;
        RECT -108.170 -176.250 -108.010 -175.460 ;
        RECT -107.670 -175.570 -107.350 -175.460 ;
        RECT -104.990 -175.320 -104.670 -175.290 ;
        RECT -104.990 -175.460 -104.170 -175.320 ;
        RECT -104.990 -175.570 -104.670 -175.460 ;
        RECT -109.950 -176.400 -108.010 -176.250 ;
        RECT -104.330 -176.250 -104.170 -175.460 ;
        RECT -103.210 -175.760 -103.050 -174.970 ;
        RECT -99.370 -174.970 -97.430 -174.820 ;
        RECT -102.710 -175.760 -102.390 -175.650 ;
        RECT -103.210 -175.900 -102.390 -175.760 ;
        RECT -102.710 -175.930 -102.390 -175.900 ;
        RECT -100.030 -175.760 -99.710 -175.650 ;
        RECT -99.370 -175.760 -99.210 -174.970 ;
        RECT -97.770 -175.120 -97.430 -174.970 ;
        RECT -95.070 -174.970 -93.130 -174.820 ;
        RECT -95.070 -175.120 -94.730 -174.970 ;
        RECT -97.750 -175.320 -97.430 -175.290 ;
        RECT -100.030 -175.900 -99.210 -175.760 ;
        RECT -98.250 -175.460 -97.430 -175.320 ;
        RECT -100.030 -175.930 -99.710 -175.900 ;
        RECT -102.730 -176.250 -102.390 -176.100 ;
        RECT -104.330 -176.400 -102.390 -176.250 ;
        RECT -100.030 -176.250 -99.690 -176.100 ;
        RECT -98.250 -176.250 -98.090 -175.460 ;
        RECT -97.750 -175.570 -97.430 -175.460 ;
        RECT -95.070 -175.320 -94.750 -175.290 ;
        RECT -95.070 -175.460 -94.250 -175.320 ;
        RECT -95.070 -175.570 -94.750 -175.460 ;
        RECT -100.030 -176.400 -98.090 -176.250 ;
        RECT -94.410 -176.250 -94.250 -175.460 ;
        RECT -93.290 -175.760 -93.130 -174.970 ;
        RECT -89.450 -174.970 -87.510 -174.820 ;
        RECT -92.790 -175.760 -92.470 -175.650 ;
        RECT -93.290 -175.900 -92.470 -175.760 ;
        RECT -92.790 -175.930 -92.470 -175.900 ;
        RECT -90.110 -175.760 -89.790 -175.650 ;
        RECT -89.450 -175.760 -89.290 -174.970 ;
        RECT -87.850 -175.120 -87.510 -174.970 ;
        RECT -85.150 -174.970 -83.210 -174.820 ;
        RECT -85.150 -175.120 -84.810 -174.970 ;
        RECT -87.830 -175.320 -87.510 -175.290 ;
        RECT -90.110 -175.900 -89.290 -175.760 ;
        RECT -88.330 -175.460 -87.510 -175.320 ;
        RECT -90.110 -175.930 -89.790 -175.900 ;
        RECT -92.810 -176.250 -92.470 -176.100 ;
        RECT -94.410 -176.400 -92.470 -176.250 ;
        RECT -90.110 -176.250 -89.770 -176.100 ;
        RECT -88.330 -176.250 -88.170 -175.460 ;
        RECT -87.830 -175.570 -87.510 -175.460 ;
        RECT -85.150 -175.320 -84.830 -175.290 ;
        RECT -85.150 -175.460 -84.330 -175.320 ;
        RECT -85.150 -175.570 -84.830 -175.460 ;
        RECT -90.110 -176.400 -88.170 -176.250 ;
        RECT -84.490 -176.250 -84.330 -175.460 ;
        RECT -83.370 -175.760 -83.210 -174.970 ;
        RECT -79.530 -174.970 -77.590 -174.820 ;
        RECT -82.870 -175.760 -82.550 -175.650 ;
        RECT -83.370 -175.900 -82.550 -175.760 ;
        RECT -82.870 -175.930 -82.550 -175.900 ;
        RECT -80.190 -175.760 -79.870 -175.650 ;
        RECT -79.530 -175.760 -79.370 -174.970 ;
        RECT -77.930 -175.120 -77.590 -174.970 ;
        RECT -75.230 -174.970 -73.290 -174.820 ;
        RECT -75.230 -175.120 -74.890 -174.970 ;
        RECT -77.910 -175.320 -77.590 -175.290 ;
        RECT -80.190 -175.900 -79.370 -175.760 ;
        RECT -78.410 -175.460 -77.590 -175.320 ;
        RECT -80.190 -175.930 -79.870 -175.900 ;
        RECT -82.890 -176.250 -82.550 -176.100 ;
        RECT -84.490 -176.400 -82.550 -176.250 ;
        RECT -80.190 -176.250 -79.850 -176.100 ;
        RECT -78.410 -176.250 -78.250 -175.460 ;
        RECT -77.910 -175.570 -77.590 -175.460 ;
        RECT -75.230 -175.320 -74.910 -175.290 ;
        RECT -75.230 -175.460 -74.410 -175.320 ;
        RECT -75.230 -175.570 -74.910 -175.460 ;
        RECT -80.190 -176.400 -78.250 -176.250 ;
        RECT -74.570 -176.250 -74.410 -175.460 ;
        RECT -73.450 -175.760 -73.290 -174.970 ;
        RECT -69.610 -174.970 -67.670 -174.820 ;
        RECT -72.950 -175.760 -72.630 -175.650 ;
        RECT -73.450 -175.900 -72.630 -175.760 ;
        RECT -72.950 -175.930 -72.630 -175.900 ;
        RECT -70.270 -175.760 -69.950 -175.650 ;
        RECT -69.610 -175.760 -69.450 -174.970 ;
        RECT -68.010 -175.120 -67.670 -174.970 ;
        RECT -65.310 -174.970 -63.370 -174.820 ;
        RECT -65.310 -175.120 -64.970 -174.970 ;
        RECT -67.990 -175.320 -67.670 -175.290 ;
        RECT -70.270 -175.900 -69.450 -175.760 ;
        RECT -68.490 -175.460 -67.670 -175.320 ;
        RECT -70.270 -175.930 -69.950 -175.900 ;
        RECT -72.970 -176.250 -72.630 -176.100 ;
        RECT -74.570 -176.400 -72.630 -176.250 ;
        RECT -70.270 -176.250 -69.930 -176.100 ;
        RECT -68.490 -176.250 -68.330 -175.460 ;
        RECT -67.990 -175.570 -67.670 -175.460 ;
        RECT -65.310 -175.320 -64.990 -175.290 ;
        RECT -65.310 -175.460 -64.490 -175.320 ;
        RECT -65.310 -175.570 -64.990 -175.460 ;
        RECT -70.270 -176.400 -68.330 -176.250 ;
        RECT -64.650 -176.250 -64.490 -175.460 ;
        RECT -63.530 -175.760 -63.370 -174.970 ;
        RECT -59.690 -174.970 -57.750 -174.820 ;
        RECT -63.030 -175.760 -62.710 -175.650 ;
        RECT -63.530 -175.900 -62.710 -175.760 ;
        RECT -63.030 -175.930 -62.710 -175.900 ;
        RECT -60.350 -175.760 -60.030 -175.650 ;
        RECT -59.690 -175.760 -59.530 -174.970 ;
        RECT -58.090 -175.120 -57.750 -174.970 ;
        RECT -55.390 -174.970 -53.450 -174.820 ;
        RECT -55.390 -175.120 -55.050 -174.970 ;
        RECT -58.070 -175.320 -57.750 -175.290 ;
        RECT -60.350 -175.900 -59.530 -175.760 ;
        RECT -58.570 -175.460 -57.750 -175.320 ;
        RECT -60.350 -175.930 -60.030 -175.900 ;
        RECT -63.050 -176.250 -62.710 -176.100 ;
        RECT -64.650 -176.400 -62.710 -176.250 ;
        RECT -60.350 -176.250 -60.010 -176.100 ;
        RECT -58.570 -176.250 -58.410 -175.460 ;
        RECT -58.070 -175.570 -57.750 -175.460 ;
        RECT -55.390 -175.320 -55.070 -175.290 ;
        RECT -55.390 -175.460 -54.570 -175.320 ;
        RECT -55.390 -175.570 -55.070 -175.460 ;
        RECT -60.350 -176.400 -58.410 -176.250 ;
        RECT -54.730 -176.250 -54.570 -175.460 ;
        RECT -53.610 -175.760 -53.450 -174.970 ;
        RECT -49.770 -174.970 -47.830 -174.820 ;
        RECT -53.110 -175.760 -52.790 -175.650 ;
        RECT -53.610 -175.900 -52.790 -175.760 ;
        RECT -53.110 -175.930 -52.790 -175.900 ;
        RECT -50.430 -175.760 -50.110 -175.650 ;
        RECT -49.770 -175.760 -49.610 -174.970 ;
        RECT -48.170 -175.120 -47.830 -174.970 ;
        RECT -45.470 -174.970 -43.530 -174.820 ;
        RECT -45.470 -175.120 -45.130 -174.970 ;
        RECT -48.150 -175.320 -47.830 -175.290 ;
        RECT -50.430 -175.900 -49.610 -175.760 ;
        RECT -48.650 -175.460 -47.830 -175.320 ;
        RECT -50.430 -175.930 -50.110 -175.900 ;
        RECT -53.130 -176.250 -52.790 -176.100 ;
        RECT -54.730 -176.400 -52.790 -176.250 ;
        RECT -50.430 -176.250 -50.090 -176.100 ;
        RECT -48.650 -176.250 -48.490 -175.460 ;
        RECT -48.150 -175.570 -47.830 -175.460 ;
        RECT -45.470 -175.320 -45.150 -175.290 ;
        RECT -45.470 -175.460 -44.650 -175.320 ;
        RECT -45.470 -175.570 -45.150 -175.460 ;
        RECT -50.430 -176.400 -48.490 -176.250 ;
        RECT -44.810 -176.250 -44.650 -175.460 ;
        RECT -43.690 -175.760 -43.530 -174.970 ;
        RECT -39.850 -174.970 -37.910 -174.820 ;
        RECT -43.190 -175.760 -42.870 -175.650 ;
        RECT -43.690 -175.900 -42.870 -175.760 ;
        RECT -43.190 -175.930 -42.870 -175.900 ;
        RECT -40.510 -175.760 -40.190 -175.650 ;
        RECT -39.850 -175.760 -39.690 -174.970 ;
        RECT -38.250 -175.120 -37.910 -174.970 ;
        RECT -35.550 -174.970 -33.610 -174.820 ;
        RECT -35.550 -175.120 -35.210 -174.970 ;
        RECT -38.230 -175.320 -37.910 -175.290 ;
        RECT -40.510 -175.900 -39.690 -175.760 ;
        RECT -38.730 -175.460 -37.910 -175.320 ;
        RECT -40.510 -175.930 -40.190 -175.900 ;
        RECT -43.210 -176.250 -42.870 -176.100 ;
        RECT -44.810 -176.400 -42.870 -176.250 ;
        RECT -40.510 -176.250 -40.170 -176.100 ;
        RECT -38.730 -176.250 -38.570 -175.460 ;
        RECT -38.230 -175.570 -37.910 -175.460 ;
        RECT -35.550 -175.320 -35.230 -175.290 ;
        RECT -35.550 -175.460 -34.730 -175.320 ;
        RECT -35.550 -175.570 -35.230 -175.460 ;
        RECT -40.510 -176.400 -38.570 -176.250 ;
        RECT -34.890 -176.250 -34.730 -175.460 ;
        RECT -33.770 -175.760 -33.610 -174.970 ;
        RECT -29.930 -174.970 -27.990 -174.820 ;
        RECT -33.270 -175.760 -32.950 -175.650 ;
        RECT -33.770 -175.900 -32.950 -175.760 ;
        RECT -33.270 -175.930 -32.950 -175.900 ;
        RECT -30.590 -175.760 -30.270 -175.650 ;
        RECT -29.930 -175.760 -29.770 -174.970 ;
        RECT -28.330 -175.120 -27.990 -174.970 ;
        RECT -25.630 -174.970 -23.690 -174.820 ;
        RECT -25.630 -175.120 -25.290 -174.970 ;
        RECT -28.310 -175.320 -27.990 -175.290 ;
        RECT -30.590 -175.900 -29.770 -175.760 ;
        RECT -28.810 -175.460 -27.990 -175.320 ;
        RECT -30.590 -175.930 -30.270 -175.900 ;
        RECT -33.290 -176.250 -32.950 -176.100 ;
        RECT -34.890 -176.400 -32.950 -176.250 ;
        RECT -30.590 -176.250 -30.250 -176.100 ;
        RECT -28.810 -176.250 -28.650 -175.460 ;
        RECT -28.310 -175.570 -27.990 -175.460 ;
        RECT -25.630 -175.320 -25.310 -175.290 ;
        RECT -25.630 -175.460 -24.810 -175.320 ;
        RECT -25.630 -175.570 -25.310 -175.460 ;
        RECT -30.590 -176.400 -28.650 -176.250 ;
        RECT -24.970 -176.250 -24.810 -175.460 ;
        RECT -23.850 -175.760 -23.690 -174.970 ;
        RECT -20.010 -174.970 -18.070 -174.820 ;
        RECT -23.350 -175.760 -23.030 -175.650 ;
        RECT -23.850 -175.900 -23.030 -175.760 ;
        RECT -23.350 -175.930 -23.030 -175.900 ;
        RECT -20.670 -175.760 -20.350 -175.650 ;
        RECT -20.010 -175.760 -19.850 -174.970 ;
        RECT -18.410 -175.120 -18.070 -174.970 ;
        RECT -15.710 -174.970 -13.770 -174.820 ;
        RECT -15.710 -175.120 -15.370 -174.970 ;
        RECT -18.390 -175.320 -18.070 -175.290 ;
        RECT -20.670 -175.900 -19.850 -175.760 ;
        RECT -18.890 -175.460 -18.070 -175.320 ;
        RECT -20.670 -175.930 -20.350 -175.900 ;
        RECT -23.370 -176.250 -23.030 -176.100 ;
        RECT -24.970 -176.400 -23.030 -176.250 ;
        RECT -20.670 -176.250 -20.330 -176.100 ;
        RECT -18.890 -176.250 -18.730 -175.460 ;
        RECT -18.390 -175.570 -18.070 -175.460 ;
        RECT -15.710 -175.320 -15.390 -175.290 ;
        RECT -15.710 -175.460 -14.890 -175.320 ;
        RECT -15.710 -175.570 -15.390 -175.460 ;
        RECT -20.670 -176.400 -18.730 -176.250 ;
        RECT -15.050 -176.250 -14.890 -175.460 ;
        RECT -13.930 -175.760 -13.770 -174.970 ;
        RECT -10.090 -174.970 -8.150 -174.820 ;
        RECT -13.430 -175.760 -13.110 -175.650 ;
        RECT -13.930 -175.900 -13.110 -175.760 ;
        RECT -13.430 -175.930 -13.110 -175.900 ;
        RECT -10.750 -175.760 -10.430 -175.650 ;
        RECT -10.090 -175.760 -9.930 -174.970 ;
        RECT -8.490 -175.120 -8.150 -174.970 ;
        RECT -5.790 -174.970 -3.850 -174.820 ;
        RECT -5.790 -175.120 -5.450 -174.970 ;
        RECT -8.470 -175.320 -8.150 -175.290 ;
        RECT -10.750 -175.900 -9.930 -175.760 ;
        RECT -8.970 -175.460 -8.150 -175.320 ;
        RECT -10.750 -175.930 -10.430 -175.900 ;
        RECT -13.450 -176.250 -13.110 -176.100 ;
        RECT -15.050 -176.400 -13.110 -176.250 ;
        RECT -10.750 -176.250 -10.410 -176.100 ;
        RECT -8.970 -176.250 -8.810 -175.460 ;
        RECT -8.470 -175.570 -8.150 -175.460 ;
        RECT -5.790 -175.320 -5.470 -175.290 ;
        RECT -5.790 -175.460 -4.970 -175.320 ;
        RECT -5.790 -175.570 -5.470 -175.460 ;
        RECT -10.750 -176.400 -8.810 -176.250 ;
        RECT -5.130 -176.250 -4.970 -175.460 ;
        RECT -4.010 -175.760 -3.850 -174.970 ;
        RECT -0.170 -174.970 1.770 -174.820 ;
        RECT -3.510 -175.760 -3.190 -175.650 ;
        RECT -4.010 -175.900 -3.190 -175.760 ;
        RECT -3.510 -175.930 -3.190 -175.900 ;
        RECT -0.830 -175.760 -0.510 -175.650 ;
        RECT -0.170 -175.760 -0.010 -174.970 ;
        RECT 1.430 -175.120 1.770 -174.970 ;
        RECT 4.130 -174.970 6.070 -174.820 ;
        RECT 4.130 -175.120 4.470 -174.970 ;
        RECT 1.450 -175.320 1.770 -175.290 ;
        RECT -0.830 -175.900 -0.010 -175.760 ;
        RECT 0.950 -175.460 1.770 -175.320 ;
        RECT -0.830 -175.930 -0.510 -175.900 ;
        RECT -3.530 -176.250 -3.190 -176.100 ;
        RECT -5.130 -176.400 -3.190 -176.250 ;
        RECT -0.830 -176.250 -0.490 -176.100 ;
        RECT 0.950 -176.250 1.110 -175.460 ;
        RECT 1.450 -175.570 1.770 -175.460 ;
        RECT 4.130 -175.320 4.450 -175.290 ;
        RECT 4.130 -175.460 4.950 -175.320 ;
        RECT 4.130 -175.570 4.450 -175.460 ;
        RECT -0.830 -176.400 1.110 -176.250 ;
        RECT 4.790 -176.250 4.950 -175.460 ;
        RECT 5.910 -175.760 6.070 -174.970 ;
        RECT 9.750 -174.970 11.690 -174.820 ;
        RECT 6.410 -175.760 6.730 -175.650 ;
        RECT 5.910 -175.900 6.730 -175.760 ;
        RECT 6.410 -175.930 6.730 -175.900 ;
        RECT 9.090 -175.760 9.410 -175.650 ;
        RECT 9.750 -175.760 9.910 -174.970 ;
        RECT 11.350 -175.120 11.690 -174.970 ;
        RECT 14.050 -174.970 15.990 -174.820 ;
        RECT 14.050 -175.120 14.390 -174.970 ;
        RECT 11.370 -175.320 11.690 -175.290 ;
        RECT 9.090 -175.900 9.910 -175.760 ;
        RECT 10.870 -175.460 11.690 -175.320 ;
        RECT 9.090 -175.930 9.410 -175.900 ;
        RECT 6.390 -176.250 6.730 -176.100 ;
        RECT 4.790 -176.400 6.730 -176.250 ;
        RECT 9.090 -176.250 9.430 -176.100 ;
        RECT 10.870 -176.250 11.030 -175.460 ;
        RECT 11.370 -175.570 11.690 -175.460 ;
        RECT 14.050 -175.320 14.370 -175.290 ;
        RECT 14.050 -175.460 14.870 -175.320 ;
        RECT 14.050 -175.570 14.370 -175.460 ;
        RECT 9.090 -176.400 11.030 -176.250 ;
        RECT 14.710 -176.250 14.870 -175.460 ;
        RECT 15.830 -175.760 15.990 -174.970 ;
        RECT 19.670 -174.970 21.610 -174.820 ;
        RECT 16.330 -175.760 16.650 -175.650 ;
        RECT 15.830 -175.900 16.650 -175.760 ;
        RECT 16.330 -175.930 16.650 -175.900 ;
        RECT 19.010 -175.760 19.330 -175.650 ;
        RECT 19.670 -175.760 19.830 -174.970 ;
        RECT 21.270 -175.120 21.610 -174.970 ;
        RECT 21.290 -175.320 21.610 -175.290 ;
        RECT 19.010 -175.900 19.830 -175.760 ;
        RECT 20.790 -175.460 21.610 -175.320 ;
        RECT 19.010 -175.930 19.330 -175.900 ;
        RECT 16.310 -176.250 16.650 -176.100 ;
        RECT 14.710 -176.400 16.650 -176.250 ;
        RECT 19.010 -176.250 19.350 -176.100 ;
        RECT 20.790 -176.250 20.950 -175.460 ;
        RECT 21.290 -175.570 21.610 -175.460 ;
        RECT 19.010 -176.400 20.950 -176.250 ;
        RECT -294.880 -177.210 -293.040 -176.730 ;
        RECT -293.120 -178.300 -292.640 -177.400 ;
        RECT -291.820 -177.530 -291.630 -176.400 ;
        RECT -287.750 -177.530 -287.560 -176.400 ;
        RECT -281.900 -177.530 -281.710 -176.400 ;
        RECT -277.830 -177.530 -277.640 -176.400 ;
        RECT -271.980 -177.530 -271.790 -176.400 ;
        RECT -267.910 -177.530 -267.720 -176.400 ;
        RECT -262.060 -177.530 -261.870 -176.400 ;
        RECT -257.990 -177.530 -257.800 -176.400 ;
        RECT -252.140 -177.530 -251.950 -176.400 ;
        RECT -248.070 -177.530 -247.880 -176.400 ;
        RECT -242.220 -177.530 -242.030 -176.400 ;
        RECT -238.150 -177.530 -237.960 -176.400 ;
        RECT -232.300 -177.530 -232.110 -176.400 ;
        RECT -228.230 -177.530 -228.040 -176.400 ;
        RECT -222.380 -177.530 -222.190 -176.400 ;
        RECT -218.310 -177.530 -218.120 -176.400 ;
        RECT -212.460 -177.530 -212.270 -176.400 ;
        RECT -208.390 -177.530 -208.200 -176.400 ;
        RECT -202.540 -177.530 -202.350 -176.400 ;
        RECT -198.470 -177.530 -198.280 -176.400 ;
        RECT -192.620 -177.530 -192.430 -176.400 ;
        RECT -188.550 -177.530 -188.360 -176.400 ;
        RECT -182.700 -177.530 -182.510 -176.400 ;
        RECT -178.630 -177.530 -178.440 -176.400 ;
        RECT -172.780 -177.530 -172.590 -176.400 ;
        RECT -168.710 -177.530 -168.520 -176.400 ;
        RECT -162.860 -177.530 -162.670 -176.400 ;
        RECT -158.790 -177.530 -158.600 -176.400 ;
        RECT -152.940 -177.530 -152.750 -176.400 ;
        RECT -148.870 -177.530 -148.680 -176.400 ;
        RECT -143.020 -177.530 -142.830 -176.400 ;
        RECT -138.950 -177.530 -138.760 -176.400 ;
        RECT -133.100 -177.530 -132.910 -176.400 ;
        RECT -129.030 -177.530 -128.840 -176.400 ;
        RECT -123.180 -177.530 -122.990 -176.400 ;
        RECT -119.110 -177.530 -118.920 -176.400 ;
        RECT -113.260 -177.530 -113.070 -176.400 ;
        RECT -109.190 -177.530 -109.000 -176.400 ;
        RECT -103.340 -177.530 -103.150 -176.400 ;
        RECT -99.270 -177.530 -99.080 -176.400 ;
        RECT -93.420 -177.530 -93.230 -176.400 ;
        RECT -89.350 -177.530 -89.160 -176.400 ;
        RECT -83.500 -177.530 -83.310 -176.400 ;
        RECT -79.430 -177.530 -79.240 -176.400 ;
        RECT -73.580 -177.530 -73.390 -176.400 ;
        RECT -69.510 -177.530 -69.320 -176.400 ;
        RECT -63.660 -177.530 -63.470 -176.400 ;
        RECT -59.590 -177.530 -59.400 -176.400 ;
        RECT -53.740 -177.530 -53.550 -176.400 ;
        RECT -49.670 -177.530 -49.480 -176.400 ;
        RECT -43.820 -177.530 -43.630 -176.400 ;
        RECT -39.750 -177.530 -39.560 -176.400 ;
        RECT -33.900 -177.530 -33.710 -176.400 ;
        RECT -29.830 -177.530 -29.640 -176.400 ;
        RECT -23.980 -177.530 -23.790 -176.400 ;
        RECT -19.910 -177.530 -19.720 -176.400 ;
        RECT -14.060 -177.530 -13.870 -176.400 ;
        RECT -9.990 -177.530 -9.800 -176.400 ;
        RECT -4.140 -177.530 -3.950 -176.400 ;
        RECT -0.070 -177.530 0.120 -176.400 ;
        RECT 5.780 -177.530 5.970 -176.400 ;
        RECT 9.850 -177.530 10.040 -176.400 ;
        RECT 15.700 -177.530 15.890 -176.400 ;
        RECT 19.770 -177.530 19.960 -176.400 ;
        RECT -291.870 -177.820 -291.550 -177.530 ;
        RECT -287.830 -177.820 -287.510 -177.530 ;
        RECT -281.950 -177.820 -281.630 -177.530 ;
        RECT -277.910 -177.820 -277.590 -177.530 ;
        RECT -272.030 -177.820 -271.710 -177.530 ;
        RECT -267.990 -177.820 -267.670 -177.530 ;
        RECT -262.110 -177.820 -261.790 -177.530 ;
        RECT -258.070 -177.820 -257.750 -177.530 ;
        RECT -252.190 -177.820 -251.870 -177.530 ;
        RECT -248.150 -177.820 -247.830 -177.530 ;
        RECT -242.270 -177.820 -241.950 -177.530 ;
        RECT -238.230 -177.820 -237.910 -177.530 ;
        RECT -232.350 -177.820 -232.030 -177.530 ;
        RECT -228.310 -177.820 -227.990 -177.530 ;
        RECT -222.430 -177.820 -222.110 -177.530 ;
        RECT -218.390 -177.820 -218.070 -177.530 ;
        RECT -212.510 -177.820 -212.190 -177.530 ;
        RECT -208.470 -177.820 -208.150 -177.530 ;
        RECT -202.590 -177.820 -202.270 -177.530 ;
        RECT -198.550 -177.820 -198.230 -177.530 ;
        RECT -192.670 -177.820 -192.350 -177.530 ;
        RECT -188.630 -177.820 -188.310 -177.530 ;
        RECT -182.750 -177.820 -182.430 -177.530 ;
        RECT -178.710 -177.820 -178.390 -177.530 ;
        RECT -172.830 -177.820 -172.510 -177.530 ;
        RECT -168.790 -177.820 -168.470 -177.530 ;
        RECT -162.910 -177.820 -162.590 -177.530 ;
        RECT -158.870 -177.820 -158.550 -177.530 ;
        RECT -152.990 -177.820 -152.670 -177.530 ;
        RECT -148.950 -177.820 -148.630 -177.530 ;
        RECT -143.070 -177.820 -142.750 -177.530 ;
        RECT -139.030 -177.820 -138.710 -177.530 ;
        RECT -133.150 -177.820 -132.830 -177.530 ;
        RECT -129.110 -177.820 -128.790 -177.530 ;
        RECT -123.230 -177.820 -122.910 -177.530 ;
        RECT -119.190 -177.820 -118.870 -177.530 ;
        RECT -113.310 -177.820 -112.990 -177.530 ;
        RECT -109.270 -177.820 -108.950 -177.530 ;
        RECT -103.390 -177.820 -103.070 -177.530 ;
        RECT -99.350 -177.820 -99.030 -177.530 ;
        RECT -93.470 -177.820 -93.150 -177.530 ;
        RECT -89.430 -177.820 -89.110 -177.530 ;
        RECT -83.550 -177.820 -83.230 -177.530 ;
        RECT -79.510 -177.820 -79.190 -177.530 ;
        RECT -73.630 -177.820 -73.310 -177.530 ;
        RECT -69.590 -177.820 -69.270 -177.530 ;
        RECT -63.710 -177.820 -63.390 -177.530 ;
        RECT -59.670 -177.820 -59.350 -177.530 ;
        RECT -53.790 -177.820 -53.470 -177.530 ;
        RECT -49.750 -177.820 -49.430 -177.530 ;
        RECT -43.870 -177.820 -43.550 -177.530 ;
        RECT -39.830 -177.820 -39.510 -177.530 ;
        RECT -33.950 -177.820 -33.630 -177.530 ;
        RECT -29.910 -177.820 -29.590 -177.530 ;
        RECT -24.030 -177.820 -23.710 -177.530 ;
        RECT -19.990 -177.820 -19.670 -177.530 ;
        RECT -14.110 -177.820 -13.790 -177.530 ;
        RECT -10.070 -177.820 -9.750 -177.530 ;
        RECT -4.190 -177.820 -3.870 -177.530 ;
        RECT -0.150 -177.820 0.170 -177.530 ;
        RECT 5.730 -177.820 6.050 -177.530 ;
        RECT 9.770 -177.820 10.090 -177.530 ;
        RECT 15.650 -177.820 15.970 -177.530 ;
        RECT 19.690 -177.820 20.010 -177.530 ;
        RECT -293.580 -178.780 -292.640 -178.300 ;
        RECT 20.780 -178.300 21.260 -177.400 ;
        RECT -288.570 -178.700 -286.880 -178.400 ;
        RECT -278.650 -178.700 -276.960 -178.400 ;
        RECT -268.730 -178.700 -267.040 -178.400 ;
        RECT -258.810 -178.700 -257.120 -178.400 ;
        RECT -248.890 -178.700 -247.200 -178.400 ;
        RECT -238.970 -178.700 -237.280 -178.400 ;
        RECT -229.050 -178.700 -227.360 -178.400 ;
        RECT -219.130 -178.700 -217.440 -178.400 ;
        RECT -209.210 -178.700 -207.520 -178.400 ;
        RECT -199.290 -178.700 -197.600 -178.400 ;
        RECT -189.370 -178.700 -187.680 -178.400 ;
        RECT -179.450 -178.700 -177.760 -178.400 ;
        RECT -169.530 -178.700 -167.840 -178.400 ;
        RECT -159.610 -178.700 -157.920 -178.400 ;
        RECT -149.690 -178.700 -148.000 -178.400 ;
        RECT -139.770 -178.700 -138.080 -178.400 ;
        RECT -129.850 -178.700 -128.160 -178.400 ;
        RECT -119.930 -178.700 -118.240 -178.400 ;
        RECT -110.010 -178.700 -108.320 -178.400 ;
        RECT -100.090 -178.700 -98.400 -178.400 ;
        RECT -90.170 -178.700 -88.480 -178.400 ;
        RECT -80.250 -178.700 -78.560 -178.400 ;
        RECT -70.330 -178.700 -68.640 -178.400 ;
        RECT -60.410 -178.700 -58.720 -178.400 ;
        RECT -50.490 -178.700 -48.800 -178.400 ;
        RECT -40.570 -178.700 -38.880 -178.400 ;
        RECT -30.650 -178.700 -28.960 -178.400 ;
        RECT -20.730 -178.700 -19.040 -178.400 ;
        RECT -10.810 -178.700 -9.120 -178.400 ;
        RECT -0.890 -178.700 0.800 -178.400 ;
        RECT 9.030 -178.700 10.720 -178.400 ;
        RECT 18.950 -178.700 20.640 -178.400 ;
        RECT -288.060 -179.400 -287.060 -178.700 ;
        RECT -278.140 -179.400 -277.140 -178.700 ;
        RECT -268.220 -179.400 -267.220 -178.700 ;
        RECT -258.300 -179.400 -257.300 -178.700 ;
        RECT -248.380 -179.400 -247.380 -178.700 ;
        RECT -238.460 -179.400 -237.460 -178.700 ;
        RECT -228.540 -179.400 -227.540 -178.700 ;
        RECT -218.620 -179.400 -217.620 -178.700 ;
        RECT -208.700 -179.400 -207.700 -178.700 ;
        RECT -198.780 -179.400 -197.780 -178.700 ;
        RECT -188.860 -179.400 -187.860 -178.700 ;
        RECT -178.940 -179.400 -177.940 -178.700 ;
        RECT -169.020 -179.400 -168.020 -178.700 ;
        RECT -159.100 -179.400 -158.100 -178.700 ;
        RECT -149.180 -179.400 -148.180 -178.700 ;
        RECT -139.260 -179.400 -138.260 -178.700 ;
        RECT -129.340 -179.400 -128.340 -178.700 ;
        RECT -119.420 -179.400 -118.420 -178.700 ;
        RECT -109.500 -179.400 -108.500 -178.700 ;
        RECT -99.580 -179.400 -98.580 -178.700 ;
        RECT -89.660 -179.400 -88.660 -178.700 ;
        RECT -79.740 -179.400 -78.740 -178.700 ;
        RECT -69.820 -179.400 -68.820 -178.700 ;
        RECT -59.900 -179.400 -58.900 -178.700 ;
        RECT -49.980 -179.400 -48.980 -178.700 ;
        RECT -40.060 -179.400 -39.060 -178.700 ;
        RECT -30.140 -179.400 -29.140 -178.700 ;
        RECT -20.220 -179.400 -19.220 -178.700 ;
        RECT -10.300 -179.400 -9.300 -178.700 ;
        RECT -0.380 -179.400 0.620 -178.700 ;
        RECT 9.540 -179.400 10.540 -178.700 ;
        RECT 19.460 -179.400 20.460 -178.700 ;
        RECT 20.780 -178.780 21.720 -178.300 ;
  END
END meta_srlatch_stack
END LIBRARY

